magic
tech sky130A
magscale 1 2
timestamp 1685641953
<< viali >>
rect 5917 9673 5951 9707
rect 6929 9673 6963 9707
rect 26525 9673 26559 9707
rect 27353 9673 27387 9707
rect 29101 9673 29135 9707
rect 30389 9673 30423 9707
rect 32505 9673 32539 9707
rect 39313 9673 39347 9707
rect 55689 9673 55723 9707
rect 56517 9673 56551 9707
rect 57345 9673 57379 9707
rect 58265 9673 58299 9707
rect 61761 9673 61795 9707
rect 62497 9673 62531 9707
rect 63417 9673 63451 9707
rect 84025 9673 84059 9707
rect 87015 9673 87049 9707
rect 92765 9673 92799 9707
rect 93501 9673 93535 9707
rect 96077 9673 96111 9707
rect 96905 9673 96939 9707
rect 99481 9673 99515 9707
rect 100493 9673 100527 9707
rect 104725 9673 104759 9707
rect 105461 9673 105495 9707
rect 106197 9673 106231 9707
rect 107577 9673 107611 9707
rect 121745 9673 121779 9707
rect 125241 9673 125275 9707
rect 126345 9673 126379 9707
rect 129565 9673 129599 9707
rect 130761 9673 130795 9707
rect 131497 9673 131531 9707
rect 133429 9673 133463 9707
rect 134165 9673 134199 9707
rect 169033 9673 169067 9707
rect 215861 9673 215895 9707
rect 259193 9673 259227 9707
rect 260021 9673 260055 9707
rect 266277 9673 266311 9707
rect 1685 9605 1719 9639
rect 2421 9605 2455 9639
rect 3249 9605 3283 9639
rect 4353 9605 4387 9639
rect 5089 9605 5123 9639
rect 5825 9605 5859 9639
rect 6837 9605 6871 9639
rect 7573 9605 7607 9639
rect 8401 9605 8435 9639
rect 9505 9605 9539 9639
rect 10241 9605 10275 9639
rect 10977 9605 11011 9639
rect 11989 9605 12023 9639
rect 12725 9605 12759 9639
rect 13553 9605 13587 9639
rect 14657 9605 14691 9639
rect 15393 9605 15427 9639
rect 16129 9605 16163 9639
rect 17141 9605 17175 9639
rect 17877 9605 17911 9639
rect 18061 9605 18095 9639
rect 18613 9605 18647 9639
rect 60749 9605 60783 9639
rect 79241 9605 79275 9639
rect 79425 9605 79459 9639
rect 83105 9605 83139 9639
rect 83933 9605 83967 9639
rect 84669 9605 84703 9639
rect 85405 9605 85439 9639
rect 175381 9605 175415 9639
rect 175565 9605 175599 9639
rect 265633 9605 265667 9639
rect 268117 9605 268151 9639
rect 8585 9537 8619 9571
rect 22477 9537 22511 9571
rect 22569 9537 22603 9571
rect 23489 9537 23523 9571
rect 24685 9537 24719 9571
rect 25697 9537 25731 9571
rect 25881 9537 25915 9571
rect 26341 9537 26375 9571
rect 27169 9537 27203 9571
rect 28917 9537 28951 9571
rect 30205 9537 30239 9571
rect 32321 9537 32355 9571
rect 35633 9537 35667 9571
rect 36277 9537 36311 9571
rect 36921 9537 36955 9571
rect 38117 9537 38151 9571
rect 38853 9537 38887 9571
rect 39497 9537 39531 9571
rect 40785 9537 40819 9571
rect 41429 9537 41463 9571
rect 42073 9537 42107 9571
rect 43269 9537 43303 9571
rect 44005 9537 44039 9571
rect 44649 9537 44683 9571
rect 45937 9537 45971 9571
rect 46581 9537 46615 9571
rect 47225 9537 47259 9571
rect 48421 9537 48455 9571
rect 49157 9537 49191 9571
rect 49801 9537 49835 9571
rect 50629 9537 50663 9571
rect 51365 9537 51399 9571
rect 52101 9537 52135 9571
rect 53113 9537 53147 9571
rect 54493 9537 54527 9571
rect 55505 9537 55539 9571
rect 56333 9537 56367 9571
rect 57161 9537 57195 9571
rect 58081 9537 58115 9571
rect 61577 9537 61611 9571
rect 62313 9537 62347 9571
rect 63233 9537 63267 9571
rect 69121 9537 69155 9571
rect 69581 9537 69615 9571
rect 71513 9537 71547 9571
rect 72157 9537 72191 9571
rect 74733 9537 74767 9571
rect 77309 9537 77343 9571
rect 79885 9537 79919 9571
rect 81633 9537 81667 9571
rect 86785 9537 86819 9571
rect 89361 9537 89395 9571
rect 90189 9537 90223 9571
rect 91569 9537 91603 9571
rect 92581 9537 92615 9571
rect 93317 9537 93351 9571
rect 94789 9537 94823 9571
rect 94973 9537 95007 9571
rect 95893 9537 95927 9571
rect 96721 9537 96755 9571
rect 99297 9537 99331 9571
rect 100309 9537 100343 9571
rect 103253 9537 103287 9571
rect 103897 9537 103931 9571
rect 104909 9537 104943 9571
rect 105645 9537 105679 9571
rect 106381 9537 106415 9571
rect 107761 9537 107795 9571
rect 108405 9537 108439 9571
rect 109049 9537 109083 9571
rect 110061 9537 110095 9571
rect 110797 9537 110831 9571
rect 111533 9537 111567 9571
rect 112913 9537 112947 9571
rect 113557 9537 113591 9571
rect 114201 9537 114235 9571
rect 115213 9537 115247 9571
rect 115949 9537 115983 9571
rect 116685 9537 116719 9571
rect 118065 9537 118099 9571
rect 118709 9537 118743 9571
rect 119353 9537 119387 9571
rect 120365 9537 120399 9571
rect 121101 9537 121135 9571
rect 121561 9537 121595 9571
rect 125057 9537 125091 9571
rect 126161 9537 126195 9571
rect 128461 9537 128495 9571
rect 129381 9537 129415 9571
rect 130577 9537 130611 9571
rect 131313 9537 131347 9571
rect 133245 9537 133279 9571
rect 133981 9537 134015 9571
rect 138121 9537 138155 9571
rect 138765 9537 138799 9571
rect 139409 9537 139443 9571
rect 140697 9537 140731 9571
rect 141341 9537 141375 9571
rect 141985 9537 142019 9571
rect 143273 9537 143307 9571
rect 143917 9537 143951 9571
rect 144561 9537 144595 9571
rect 145849 9537 145883 9571
rect 146493 9537 146527 9571
rect 147137 9537 147171 9571
rect 148425 9537 148459 9571
rect 149069 9537 149103 9571
rect 149713 9537 149747 9571
rect 151001 9537 151035 9571
rect 151645 9537 151679 9571
rect 152289 9537 152323 9571
rect 153577 9537 153611 9571
rect 154221 9537 154255 9571
rect 154865 9537 154899 9571
rect 156521 9537 156555 9571
rect 157441 9537 157475 9571
rect 159005 9537 159039 9571
rect 159741 9537 159775 9571
rect 161305 9537 161339 9571
rect 162133 9537 162167 9571
rect 162777 9537 162811 9571
rect 162961 9537 162995 9571
rect 163881 9537 163915 9571
rect 164709 9537 164743 9571
rect 165537 9537 165571 9571
rect 166641 9537 166675 9571
rect 167285 9537 167319 9571
rect 167469 9537 167503 9571
rect 167653 9537 167687 9571
rect 168849 9537 168883 9571
rect 169585 9537 169619 9571
rect 171701 9537 171735 9571
rect 172253 9537 172287 9571
rect 174001 9537 174035 9571
rect 176669 9537 176703 9571
rect 177773 9537 177807 9571
rect 178049 9537 178083 9571
rect 179153 9537 179187 9571
rect 180533 9537 180567 9571
rect 180717 9537 180751 9571
rect 181821 9537 181855 9571
rect 182557 9537 182591 9571
rect 184305 9537 184339 9571
rect 186881 9537 186915 9571
rect 188629 9537 188663 9571
rect 190837 9537 190871 9571
rect 192033 9537 192067 9571
rect 192769 9537 192803 9571
rect 194609 9537 194643 9571
rect 195345 9537 195379 9571
rect 196357 9537 196391 9571
rect 197645 9537 197679 9571
rect 197829 9537 197863 9571
rect 198289 9537 198323 9571
rect 202337 9537 202371 9571
rect 203073 9537 203107 9571
rect 205833 9537 205867 9571
rect 206569 9537 206603 9571
rect 207673 9537 207707 9571
rect 208317 9537 208351 9571
rect 208961 9537 208995 9571
rect 210249 9537 210283 9571
rect 210893 9537 210927 9571
rect 211537 9537 211571 9571
rect 212825 9537 212859 9571
rect 213469 9537 213503 9571
rect 214113 9537 214147 9571
rect 215401 9537 215435 9571
rect 216045 9537 216079 9571
rect 216689 9537 216723 9571
rect 217977 9537 218011 9571
rect 218621 9537 218655 9571
rect 219265 9537 219299 9571
rect 220553 9537 220587 9571
rect 221197 9537 221231 9571
rect 221841 9537 221875 9571
rect 223129 9537 223163 9571
rect 223865 9537 223899 9571
rect 224785 9541 224819 9575
rect 228097 9537 228131 9571
rect 228833 9537 228867 9571
rect 229661 9537 229695 9571
rect 230673 9537 230707 9571
rect 230857 9537 230891 9571
rect 231777 9537 231811 9571
rect 233249 9537 233283 9571
rect 234813 9537 234847 9571
rect 234997 9537 235031 9571
rect 235825 9537 235859 9571
rect 239965 9537 239999 9571
rect 240977 9537 241011 9571
rect 242357 9537 242391 9571
rect 243645 9537 243679 9571
rect 244381 9537 244415 9571
rect 245117 9537 245151 9571
rect 246405 9537 246439 9571
rect 247969 9537 248003 9571
rect 249349 9537 249383 9571
rect 251557 9537 251591 9571
rect 253857 9537 253891 9571
rect 256433 9537 256467 9571
rect 257997 9537 258031 9571
rect 258089 9537 258123 9571
rect 259009 9537 259043 9571
rect 260205 9537 260239 9571
rect 260849 9537 260883 9571
rect 261769 9537 261803 9571
rect 262597 9537 262631 9571
rect 263425 9537 263459 9571
rect 264253 9537 264287 9571
rect 264897 9537 264931 9571
rect 265265 9537 265299 9571
rect 266093 9537 266127 9571
rect 267105 9537 267139 9571
rect 267933 9537 267967 9571
rect 268761 9537 268795 9571
rect 269129 9537 269163 9571
rect 269589 9537 269623 9571
rect 270141 9537 270175 9571
rect 12173 9469 12207 9503
rect 23305 9469 23339 9503
rect 24501 9469 24535 9503
rect 25513 9469 25547 9503
rect 54309 9469 54343 9503
rect 69857 9469 69891 9503
rect 72433 9469 72467 9503
rect 75009 9469 75043 9503
rect 77585 9469 77619 9503
rect 80161 9469 80195 9503
rect 81909 9469 81943 9503
rect 89177 9469 89211 9503
rect 127909 9469 127943 9503
rect 128277 9469 128311 9503
rect 157257 9469 157291 9503
rect 158821 9469 158855 9503
rect 160017 9469 160051 9503
rect 161121 9469 161155 9503
rect 161949 9469 161983 9503
rect 163697 9469 163731 9503
rect 164525 9469 164559 9503
rect 165353 9469 165387 9503
rect 166457 9469 166491 9503
rect 172529 9469 172563 9503
rect 179429 9469 179463 9503
rect 182005 9469 182039 9503
rect 182833 9469 182867 9503
rect 184581 9469 184615 9503
rect 187157 9469 187191 9503
rect 189457 9469 189491 9503
rect 189733 9469 189767 9503
rect 197461 9469 197495 9503
rect 234629 9469 234663 9503
rect 241253 9469 241287 9503
rect 242541 9469 242575 9503
rect 246681 9469 246715 9503
rect 249625 9469 249659 9503
rect 251833 9469 251867 9503
rect 254133 9469 254167 9503
rect 256709 9469 256743 9503
rect 260665 9469 260699 9503
rect 261585 9469 261619 9503
rect 262413 9469 262447 9503
rect 263241 9469 263275 9503
rect 265081 9469 265115 9503
rect 265449 9469 265483 9503
rect 266921 9469 266955 9503
rect 267749 9469 267783 9503
rect 268577 9469 268611 9503
rect 270417 9469 270451 9503
rect 2605 9401 2639 9435
rect 9689 9401 9723 9435
rect 12909 9401 12943 9435
rect 13737 9401 13771 9435
rect 15577 9401 15611 9435
rect 16313 9401 16347 9435
rect 49617 9401 49651 9435
rect 51181 9401 51215 9435
rect 61301 9401 61335 9435
rect 83289 9401 83323 9435
rect 84853 9401 84887 9435
rect 85589 9401 85623 9435
rect 89545 9401 89579 9435
rect 90373 9401 90407 9435
rect 91753 9401 91787 9435
rect 108865 9401 108899 9435
rect 111349 9401 111383 9435
rect 114017 9401 114051 9435
rect 120181 9401 120215 9435
rect 143733 9401 143767 9435
rect 146309 9401 146343 9435
rect 151461 9401 151495 9435
rect 153393 9401 153427 9435
rect 154681 9401 154715 9435
rect 156705 9401 156739 9435
rect 169769 9401 169803 9435
rect 192217 9401 192251 9435
rect 192953 9401 192987 9435
rect 194793 9401 194827 9435
rect 195529 9401 195563 9435
rect 196541 9401 196575 9435
rect 198473 9401 198507 9435
rect 202521 9401 202555 9435
rect 208133 9401 208167 9435
rect 213929 9401 213963 9435
rect 228281 9401 228315 9435
rect 229017 9401 229051 9435
rect 229845 9401 229879 9435
rect 231961 9401 231995 9435
rect 233433 9401 233467 9435
rect 236009 9401 236043 9435
rect 243829 9401 243863 9435
rect 264437 9401 264471 9435
rect 265817 9401 265851 9435
rect 268945 9401 268979 9435
rect 1777 9333 1811 9367
rect 3341 9333 3375 9367
rect 4445 9333 4479 9367
rect 5181 9333 5215 9367
rect 7665 9333 7699 9367
rect 10333 9333 10367 9367
rect 11069 9333 11103 9367
rect 14749 9333 14783 9367
rect 17233 9333 17267 9367
rect 18705 9333 18739 9367
rect 22753 9333 22787 9367
rect 23673 9333 23707 9367
rect 24869 9333 24903 9367
rect 25145 9333 25179 9367
rect 35449 9333 35483 9367
rect 36093 9333 36127 9367
rect 36737 9333 36771 9367
rect 37933 9333 37967 9367
rect 38669 9333 38703 9367
rect 40601 9333 40635 9367
rect 41245 9333 41279 9367
rect 41889 9333 41923 9367
rect 43085 9333 43119 9367
rect 43821 9333 43855 9367
rect 44465 9333 44499 9367
rect 45753 9333 45787 9367
rect 46397 9333 46431 9367
rect 47041 9333 47075 9367
rect 48237 9333 48271 9367
rect 48973 9333 49007 9367
rect 50445 9333 50479 9367
rect 51917 9333 51951 9367
rect 52929 9333 52963 9367
rect 54677 9333 54711 9367
rect 60841 9333 60875 9367
rect 71329 9333 71363 9367
rect 103713 9333 103747 9367
rect 108221 9333 108255 9367
rect 109877 9333 109911 9367
rect 110613 9333 110647 9367
rect 112729 9333 112763 9367
rect 113373 9333 113407 9367
rect 115029 9333 115063 9367
rect 115765 9333 115799 9367
rect 116501 9333 116535 9367
rect 117881 9333 117915 9367
rect 118525 9333 118559 9367
rect 119169 9333 119203 9367
rect 120917 9333 120951 9367
rect 128645 9333 128679 9367
rect 138581 9333 138615 9367
rect 139225 9333 139259 9367
rect 140513 9333 140547 9367
rect 141157 9333 141191 9367
rect 141801 9333 141835 9367
rect 143089 9333 143123 9367
rect 144377 9333 144411 9367
rect 145665 9333 145699 9367
rect 146953 9333 146987 9367
rect 148241 9333 148275 9367
rect 148885 9333 148919 9367
rect 149529 9333 149563 9367
rect 150817 9333 150851 9367
rect 152105 9333 152139 9367
rect 154037 9333 154071 9367
rect 157625 9333 157659 9367
rect 159189 9333 159223 9367
rect 161489 9333 161523 9367
rect 162317 9333 162351 9367
rect 163145 9333 163179 9367
rect 164065 9333 164099 9367
rect 164893 9333 164927 9367
rect 165721 9333 165755 9367
rect 166825 9333 166859 9367
rect 174231 9333 174265 9367
rect 176761 9333 176795 9367
rect 188445 9333 188479 9367
rect 190929 9333 190963 9367
rect 203257 9333 203291 9367
rect 206385 9333 206419 9367
rect 207489 9333 207523 9367
rect 208777 9333 208811 9367
rect 210065 9333 210099 9367
rect 210709 9333 210743 9367
rect 211353 9333 211387 9367
rect 212641 9333 212675 9367
rect 213285 9333 213319 9367
rect 215217 9333 215251 9367
rect 216505 9333 216539 9367
rect 217793 9333 217827 9367
rect 218437 9333 218471 9367
rect 219081 9333 219115 9367
rect 220369 9333 220403 9367
rect 221013 9333 221047 9367
rect 221657 9333 221691 9367
rect 222945 9333 222979 9367
rect 224049 9333 224083 9367
rect 224601 9333 224635 9367
rect 231041 9333 231075 9367
rect 244473 9333 244507 9367
rect 245209 9333 245243 9367
rect 248061 9333 248095 9367
rect 258273 9333 258307 9367
rect 261033 9333 261067 9367
rect 261953 9333 261987 9367
rect 262781 9333 262815 9367
rect 263609 9333 263643 9367
rect 267289 9333 267323 9367
rect 269221 9333 269255 9367
rect 269681 9333 269715 9367
rect 1777 9129 1811 9163
rect 23949 9129 23983 9163
rect 30389 9129 30423 9163
rect 32137 9129 32171 9163
rect 33057 9129 33091 9163
rect 35173 9129 35207 9163
rect 53297 9129 53331 9163
rect 53849 9129 53883 9163
rect 54953 9129 54987 9163
rect 55689 9129 55723 9163
rect 56609 9129 56643 9163
rect 57253 9129 57287 9163
rect 58541 9129 58575 9163
rect 62221 9129 62255 9163
rect 62773 9129 62807 9163
rect 88441 9129 88475 9163
rect 90189 9129 90223 9163
rect 91753 9129 91787 9163
rect 93685 9129 93719 9163
rect 98929 9129 98963 9163
rect 100585 9129 100619 9163
rect 101229 9129 101263 9163
rect 107025 9129 107059 9163
rect 124413 9129 124447 9163
rect 124689 9129 124723 9163
rect 126253 9129 126287 9163
rect 130577 9129 130611 9163
rect 131405 9129 131439 9163
rect 133061 9129 133095 9163
rect 134073 9129 134107 9163
rect 134717 9129 134751 9163
rect 176853 9129 176887 9163
rect 177589 9129 177623 9163
rect 192769 9129 192803 9163
rect 195805 9129 195839 9163
rect 199117 9129 199151 9163
rect 203441 9129 203475 9163
rect 204085 9129 204119 9163
rect 228373 9129 228407 9163
rect 233985 9129 234019 9163
rect 236837 9129 236871 9163
rect 252523 9129 252557 9163
rect 259377 9129 259411 9163
rect 261769 9129 261803 9163
rect 262689 9129 262723 9163
rect 270601 9129 270635 9163
rect 121101 9061 121135 9095
rect 170229 9061 170263 9095
rect 174277 9061 174311 9095
rect 182097 9061 182131 9095
rect 223773 9061 223807 9095
rect 268853 9061 268887 9095
rect 23213 8993 23247 9027
rect 25513 8993 25547 9027
rect 31493 8993 31527 9027
rect 31769 8993 31803 9027
rect 60657 8993 60691 9027
rect 66821 8993 66855 9027
rect 72065 8993 72099 9027
rect 73445 8993 73479 9027
rect 81265 8993 81299 9027
rect 81541 8993 81575 9027
rect 82829 8993 82863 9027
rect 86417 8993 86451 9027
rect 94973 8993 95007 9027
rect 95985 8993 96019 9027
rect 99205 8993 99239 9027
rect 123401 8993 123435 9027
rect 128553 8993 128587 9027
rect 128829 8993 128863 9027
rect 156153 8993 156187 9027
rect 157349 8993 157383 9027
rect 184305 8993 184339 9027
rect 185593 8993 185627 9027
rect 186881 8993 186915 9027
rect 189457 8993 189491 9027
rect 197645 8993 197679 9027
rect 197921 8993 197955 9027
rect 230673 8993 230707 9027
rect 232789 8993 232823 9027
rect 255053 8993 255087 9027
rect 256433 8993 256467 9027
rect 257721 8993 257755 9027
rect 265817 8993 265851 9027
rect 3157 8925 3191 8959
rect 8309 8925 8343 8959
rect 13461 8925 13495 8959
rect 20269 8925 20303 8959
rect 20913 8925 20947 8959
rect 21097 8925 21131 8959
rect 21189 8925 21223 8959
rect 21649 8925 21683 8959
rect 22109 8925 22143 8959
rect 22201 8925 22235 8959
rect 22937 8925 22971 8959
rect 23765 8925 23799 8959
rect 24685 8925 24719 8959
rect 25789 8925 25823 8959
rect 26709 8925 26743 8959
rect 27077 8925 27111 8959
rect 27169 8925 27203 8959
rect 27813 8925 27847 8959
rect 27997 8925 28031 8959
rect 28641 8925 28675 8959
rect 28825 8925 28859 8959
rect 30113 8925 30147 8959
rect 30205 8925 30239 8959
rect 30757 8925 30791 8959
rect 30941 8925 30975 8959
rect 31953 8925 31987 8959
rect 32873 8925 32907 8959
rect 40325 8925 40359 8959
rect 45477 8925 45511 8959
rect 53113 8925 53147 8959
rect 53665 8925 53699 8959
rect 54585 8925 54619 8959
rect 54769 8925 54803 8959
rect 55505 8925 55539 8959
rect 56333 8925 56367 8959
rect 56425 8925 56459 8959
rect 56885 8925 56919 8959
rect 57069 8925 57103 8959
rect 57621 8925 57655 8959
rect 57897 8925 57931 8959
rect 58081 8925 58115 8959
rect 58909 8925 58943 8959
rect 59093 8925 59127 8959
rect 59737 8925 59771 8959
rect 59921 8925 59955 8959
rect 60841 8925 60875 8959
rect 61853 8925 61887 8959
rect 62037 8925 62071 8959
rect 62405 8925 62439 8959
rect 62589 8925 62623 8959
rect 63233 8925 63267 8959
rect 63417 8925 63451 8959
rect 64061 8925 64095 8959
rect 64245 8925 64279 8959
rect 64981 8925 65015 8959
rect 65073 8925 65107 8959
rect 66085 8925 66119 8959
rect 66255 8935 66289 8969
rect 67005 8925 67039 8959
rect 70041 8925 70075 8959
rect 72341 8925 72375 8959
rect 73721 8925 73755 8959
rect 74733 8925 74767 8959
rect 75009 8925 75043 8959
rect 77217 8925 77251 8959
rect 77493 8925 77527 8959
rect 78689 8925 78723 8959
rect 78965 8925 78999 8959
rect 82645 8925 82679 8959
rect 86693 8925 86727 8959
rect 88257 8925 88291 8959
rect 89085 8925 89119 8959
rect 89177 8925 89211 8959
rect 89913 8925 89947 8959
rect 90005 8925 90039 8959
rect 90741 8925 90775 8959
rect 90833 8925 90867 8959
rect 91569 8925 91603 8959
rect 92397 8925 92431 8959
rect 92489 8925 92523 8959
rect 93041 8925 93075 8959
rect 93409 8925 93443 8959
rect 93501 8925 93535 8959
rect 94145 8925 94179 8959
rect 94329 8925 94363 8959
rect 95157 8925 95191 8959
rect 96997 8925 97031 8959
rect 97089 8925 97123 8959
rect 97733 8925 97767 8959
rect 97917 8925 97951 8959
rect 98101 8925 98135 8959
rect 98561 8925 98595 8959
rect 98745 8925 98779 8959
rect 99389 8925 99423 8959
rect 99941 8925 99975 8959
rect 100309 8925 100343 8959
rect 100401 8925 100435 8959
rect 101045 8925 101079 8959
rect 107209 8925 107243 8959
rect 112361 8925 112395 8959
rect 117513 8925 117547 8959
rect 120917 8925 120951 8959
rect 121653 8925 121687 8959
rect 121745 8925 121779 8959
rect 122665 8925 122699 8959
rect 122757 8925 122791 8959
rect 123585 8925 123619 8959
rect 124137 8925 124171 8959
rect 124229 8925 124263 8959
rect 125057 8925 125091 8959
rect 125241 8925 125275 8959
rect 125885 8925 125919 8959
rect 126069 8925 126103 8959
rect 126713 8925 126747 8959
rect 126897 8925 126931 8959
rect 127633 8925 127667 8959
rect 127817 8925 127851 8959
rect 130209 8925 130243 8959
rect 130393 8925 130427 8959
rect 131037 8925 131071 8959
rect 131221 8925 131255 8959
rect 131865 8925 131899 8959
rect 132049 8925 132083 8959
rect 132785 8925 132819 8959
rect 132877 8925 132911 8959
rect 133797 8925 133831 8959
rect 133889 8925 133923 8959
rect 134533 8925 134567 8959
rect 139777 8925 139811 8959
rect 144929 8925 144963 8959
rect 150081 8925 150115 8959
rect 155233 8925 155267 8959
rect 156337 8925 156371 8959
rect 157073 8925 157107 8959
rect 157165 8925 157199 8959
rect 158637 8925 158671 8959
rect 159649 8925 159683 8959
rect 160385 8925 160419 8959
rect 161581 8925 161615 8959
rect 161949 8925 161983 8959
rect 163145 8925 163179 8959
rect 163789 8925 163823 8959
rect 164985 8925 165019 8959
rect 166181 8925 166215 8959
rect 166549 8925 166583 8959
rect 167377 8925 167411 8959
rect 168941 8925 168975 8959
rect 170045 8925 170079 8959
rect 174093 8925 174127 8959
rect 175289 8925 175323 8959
rect 176761 8925 176795 8959
rect 177497 8925 177531 8959
rect 180441 8925 180475 8959
rect 181913 8925 181947 8959
rect 184581 8925 184615 8959
rect 185869 8925 185903 8959
rect 187157 8925 187191 8959
rect 189733 8925 189767 8959
rect 190745 8925 190779 8959
rect 190929 8925 190963 8959
rect 191573 8925 191607 8959
rect 191757 8925 191791 8959
rect 192401 8925 192435 8959
rect 192585 8925 192619 8959
rect 193321 8925 193355 8959
rect 193413 8925 193447 8959
rect 194701 8925 194735 8959
rect 194793 8925 194827 8959
rect 195529 8925 195563 8959
rect 195621 8925 195655 8959
rect 196357 8925 196391 8959
rect 196449 8925 196483 8959
rect 198933 8925 198967 8959
rect 199761 8925 199795 8959
rect 199945 8925 199979 8959
rect 200681 8925 200715 8959
rect 200773 8925 200807 8959
rect 201417 8925 201451 8959
rect 201601 8925 201635 8959
rect 202337 8925 202371 8959
rect 202429 8925 202463 8959
rect 203073 8925 203107 8959
rect 203257 8925 203291 8959
rect 203901 8925 203935 8959
rect 211721 8925 211755 8959
rect 216873 8925 216907 8959
rect 222025 8925 222059 8959
rect 223405 8925 223439 8959
rect 223589 8925 223623 8959
rect 224325 8925 224359 8959
rect 224417 8925 224451 8959
rect 225613 8925 225647 8959
rect 225705 8925 225739 8959
rect 226441 8925 226475 8959
rect 226533 8925 226567 8959
rect 227177 8925 227211 8959
rect 227361 8925 227395 8959
rect 228097 8925 228131 8959
rect 228189 8925 228223 8959
rect 228833 8925 228867 8959
rect 229017 8925 229051 8959
rect 229661 8925 229695 8959
rect 229845 8925 229879 8959
rect 230029 8925 230063 8959
rect 230949 8925 230983 8959
rect 231961 8925 231995 8959
rect 232145 8925 232179 8959
rect 232329 8925 232363 8959
rect 232973 8925 233007 8959
rect 233617 8925 233651 8959
rect 233801 8925 233835 8959
rect 234537 8925 234571 8959
rect 234629 8925 234663 8959
rect 235825 8925 235859 8959
rect 236009 8925 236043 8959
rect 236193 8925 236227 8959
rect 236653 8925 236687 8959
rect 241253 8925 241287 8959
rect 241529 8925 241563 8959
rect 245025 8925 245059 8959
rect 246221 8925 246255 8959
rect 247141 8925 247175 8959
rect 247417 8925 247451 8959
rect 248705 8925 248739 8959
rect 250177 8925 250211 8959
rect 251373 8925 251407 8959
rect 252293 8925 252327 8959
rect 253765 8925 253799 8959
rect 254041 8925 254075 8959
rect 255329 8925 255363 8959
rect 256709 8925 256743 8959
rect 257997 8925 258031 8959
rect 259101 8925 259135 8959
rect 259193 8925 259227 8959
rect 259837 8925 259871 8959
rect 260021 8925 260055 8959
rect 260665 8925 260699 8959
rect 260849 8925 260883 8959
rect 261677 8925 261711 8959
rect 262321 8925 262355 8959
rect 263425 8925 263459 8959
rect 263609 8925 263643 8959
rect 264253 8925 264287 8959
rect 264529 8925 264563 8959
rect 267749 8925 267783 8959
rect 268669 8925 268703 8959
rect 269313 8925 269347 8959
rect 3341 8857 3375 8891
rect 8493 8857 8527 8891
rect 13645 8857 13679 8891
rect 89361 8857 89395 8891
rect 92673 8857 92707 8891
rect 95617 8857 95651 8891
rect 123217 8857 123251 8891
rect 159189 8857 159223 8891
rect 161029 8857 161063 8891
rect 162317 8857 162351 8891
rect 164157 8857 164191 8891
rect 165353 8857 165387 8891
rect 167745 8857 167779 8891
rect 169309 8857 169343 8891
rect 180625 8857 180659 8891
rect 262597 8857 262631 8891
rect 266829 8857 266863 8891
rect 270141 8857 270175 8891
rect 270509 8857 270543 8891
rect 20453 8789 20487 8823
rect 21373 8789 21407 8823
rect 22385 8789 22419 8823
rect 24777 8789 24811 8823
rect 27353 8789 27387 8823
rect 28181 8789 28215 8823
rect 29009 8789 29043 8823
rect 31125 8789 31159 8823
rect 40141 8789 40175 8823
rect 45293 8789 45327 8823
rect 54217 8789 54251 8823
rect 58265 8789 58299 8823
rect 59277 8789 59311 8823
rect 60105 8789 60139 8823
rect 61025 8789 61059 8823
rect 61485 8789 61519 8823
rect 63601 8789 63635 8823
rect 64429 8789 64463 8823
rect 65257 8789 65291 8823
rect 66453 8789 66487 8823
rect 67189 8789 67223 8823
rect 69857 8789 69891 8823
rect 91017 8789 91051 8823
rect 94513 8789 94547 8823
rect 95341 8789 95375 8823
rect 97273 8789 97307 8823
rect 99573 8789 99607 8823
rect 112177 8789 112211 8823
rect 117329 8789 117363 8823
rect 121929 8789 121963 8823
rect 122941 8789 122975 8823
rect 123769 8789 123803 8823
rect 125425 8789 125459 8823
rect 127081 8789 127115 8823
rect 128001 8789 128035 8823
rect 132233 8789 132267 8823
rect 133429 8789 133463 8823
rect 139593 8789 139627 8823
rect 144745 8789 144779 8823
rect 149897 8789 149931 8823
rect 155049 8789 155083 8823
rect 156521 8789 156555 8823
rect 165997 8789 166031 8823
rect 175381 8789 175415 8823
rect 191113 8789 191147 8823
rect 191941 8789 191975 8823
rect 193597 8789 193631 8823
rect 194977 8789 195011 8823
rect 195345 8789 195379 8823
rect 196633 8789 196667 8823
rect 200129 8789 200163 8823
rect 200957 8789 200991 8823
rect 201785 8789 201819 8823
rect 202613 8789 202647 8823
rect 211537 8789 211571 8823
rect 216689 8789 216723 8823
rect 221841 8789 221875 8823
rect 224601 8789 224635 8823
rect 225889 8789 225923 8823
rect 226717 8789 226751 8823
rect 227545 8789 227579 8823
rect 229201 8789 229235 8823
rect 233157 8789 233191 8823
rect 234813 8789 234847 8823
rect 245117 8789 245151 8823
rect 246313 8789 246347 8823
rect 248797 8789 248831 8823
rect 250269 8789 250303 8823
rect 251465 8789 251499 8823
rect 260205 8789 260239 8823
rect 261033 8789 261067 8823
rect 263793 8789 263827 8823
rect 266185 8789 266219 8823
rect 266921 8789 266955 8823
rect 267841 8789 267875 8823
rect 21373 8585 21407 8619
rect 24041 8585 24075 8619
rect 26525 8585 26559 8619
rect 27445 8585 27479 8619
rect 28181 8585 28215 8619
rect 28917 8585 28951 8619
rect 29837 8585 29871 8619
rect 31033 8585 31067 8619
rect 33149 8585 33183 8619
rect 54861 8585 54895 8619
rect 55873 8585 55907 8619
rect 56609 8585 56643 8619
rect 57345 8585 57379 8619
rect 58817 8585 58851 8619
rect 59553 8585 59587 8619
rect 60289 8585 60323 8619
rect 61669 8585 61703 8619
rect 62589 8585 62623 8619
rect 63969 8585 64003 8619
rect 64705 8585 64739 8619
rect 88993 8585 89027 8619
rect 90833 8585 90867 8619
rect 91937 8585 91971 8619
rect 93409 8585 93443 8619
rect 94605 8585 94639 8619
rect 95065 8585 95099 8619
rect 95433 8585 95467 8619
rect 96169 8585 96203 8619
rect 96905 8585 96939 8619
rect 97549 8585 97583 8619
rect 98285 8585 98319 8619
rect 99849 8585 99883 8619
rect 121653 8585 121687 8619
rect 122389 8585 122423 8619
rect 123217 8585 123251 8619
rect 124045 8585 124079 8619
rect 125609 8585 125643 8619
rect 126989 8585 127023 8619
rect 127725 8585 127759 8619
rect 128277 8585 128311 8619
rect 130577 8585 130611 8619
rect 132141 8585 132175 8619
rect 134533 8585 134567 8619
rect 156153 8585 156187 8619
rect 224693 8585 224727 8619
rect 225521 8585 225555 8619
rect 226257 8585 226291 8619
rect 226993 8585 227027 8619
rect 228465 8585 228499 8619
rect 229201 8585 229235 8619
rect 230949 8585 230983 8619
rect 231685 8585 231719 8619
rect 232605 8585 232639 8619
rect 234445 8585 234479 8619
rect 236285 8585 236319 8619
rect 258273 8585 258307 8619
rect 259193 8585 259227 8619
rect 259929 8585 259963 8619
rect 260481 8585 260515 8619
rect 262321 8585 262355 8619
rect 265817 8585 265851 8619
rect 270509 8585 270543 8619
rect 22385 8517 22419 8551
rect 23397 8517 23431 8551
rect 89361 8517 89395 8551
rect 223865 8517 223899 8551
rect 264253 8517 264287 8551
rect 264897 8517 264931 8551
rect 266921 8517 266955 8551
rect 21189 8449 21223 8483
rect 22201 8449 22235 8483
rect 22845 8449 22879 8483
rect 23765 8449 23799 8483
rect 23857 8449 23891 8483
rect 24869 8449 24903 8483
rect 25881 8449 25915 8483
rect 26157 8449 26191 8483
rect 26341 8449 26375 8483
rect 27261 8449 27295 8483
rect 27997 8449 28031 8483
rect 28733 8449 28767 8483
rect 29561 8449 29595 8483
rect 29653 8449 29687 8483
rect 30849 8449 30883 8483
rect 32873 8449 32907 8483
rect 32965 8449 32999 8483
rect 33701 8449 33735 8483
rect 54677 8449 54711 8483
rect 55597 8449 55631 8483
rect 55689 8449 55723 8483
rect 57161 8449 57195 8483
rect 58633 8449 58667 8483
rect 59369 8449 59403 8483
rect 60105 8449 60139 8483
rect 60841 8449 60875 8483
rect 62221 8449 62255 8483
rect 62405 8449 62439 8483
rect 63785 8449 63819 8483
rect 64521 8449 64555 8483
rect 65349 8449 65383 8483
rect 66085 8449 66119 8483
rect 67281 8449 67315 8483
rect 74273 8449 74307 8483
rect 74549 8449 74583 8483
rect 76481 8449 76515 8483
rect 88809 8449 88843 8483
rect 89729 8449 89763 8483
rect 89913 8449 89947 8483
rect 90649 8449 90683 8483
rect 91293 8449 91327 8483
rect 91569 8449 91603 8483
rect 91753 8449 91787 8483
rect 93225 8449 93259 8483
rect 94421 8449 94455 8483
rect 94881 8449 94915 8483
rect 95801 8449 95835 8483
rect 95985 8449 96019 8483
rect 96721 8449 96755 8483
rect 97365 8449 97399 8483
rect 98101 8449 98135 8483
rect 99665 8449 99699 8483
rect 121469 8449 121503 8483
rect 122205 8449 122239 8483
rect 123033 8449 123067 8483
rect 123861 8449 123895 8483
rect 125425 8449 125459 8483
rect 126805 8449 126839 8483
rect 127541 8449 127575 8483
rect 128093 8449 128127 8483
rect 129197 8449 129231 8483
rect 130393 8449 130427 8483
rect 131957 8449 131991 8483
rect 132877 8449 132911 8483
rect 134257 8449 134291 8483
rect 134349 8449 134383 8483
rect 155969 8449 156003 8483
rect 156889 8449 156923 8483
rect 157993 8449 158027 8483
rect 158545 8449 158579 8483
rect 158913 8449 158947 8483
rect 160201 8449 160235 8483
rect 161213 8449 161247 8483
rect 161765 8449 161799 8483
rect 162133 8449 162167 8483
rect 163329 8449 163363 8483
rect 163697 8449 163731 8483
rect 164709 8449 164743 8483
rect 165077 8449 165111 8483
rect 166365 8449 166399 8483
rect 166457 8449 166491 8483
rect 167009 8449 167043 8483
rect 167377 8449 167411 8483
rect 186973 8449 187007 8483
rect 190377 8449 190411 8483
rect 191113 8449 191147 8483
rect 192401 8449 192435 8483
rect 192493 8449 192527 8483
rect 192677 8449 192711 8483
rect 193137 8449 193171 8483
rect 193873 8449 193907 8483
rect 195437 8449 195471 8483
rect 195621 8449 195655 8483
rect 196081 8449 196115 8483
rect 197369 8449 197403 8483
rect 197553 8449 197587 8483
rect 198381 8449 198415 8483
rect 198565 8449 198599 8483
rect 199025 8449 199059 8483
rect 199761 8449 199795 8483
rect 200589 8449 200623 8483
rect 201325 8449 201359 8483
rect 202521 8449 202555 8483
rect 202705 8449 202739 8483
rect 203349 8449 203383 8483
rect 203533 8449 203567 8483
rect 223681 8449 223715 8483
rect 224509 8449 224543 8483
rect 225337 8449 225371 8483
rect 226073 8449 226107 8483
rect 226809 8449 226843 8483
rect 228097 8449 228131 8483
rect 228281 8449 228315 8483
rect 229017 8449 229051 8483
rect 230029 8449 230063 8483
rect 230121 8449 230155 8483
rect 230305 8449 230339 8483
rect 230765 8449 230799 8483
rect 231501 8449 231535 8483
rect 232421 8449 232455 8483
rect 233617 8449 233651 8483
rect 233801 8449 233835 8483
rect 234261 8449 234295 8483
rect 235273 8449 235307 8483
rect 235457 8449 235491 8483
rect 236101 8449 236135 8483
rect 256709 8449 256743 8483
rect 258089 8449 258123 8483
rect 259101 8449 259135 8483
rect 259745 8449 259779 8483
rect 260297 8449 260331 8483
rect 261309 8449 261343 8483
rect 262137 8449 262171 8483
rect 262965 8449 262999 8483
rect 265357 8449 265391 8483
rect 265725 8449 265759 8483
rect 266737 8449 266771 8483
rect 267657 8449 267691 8483
rect 268393 8449 268427 8483
rect 269589 8449 269623 8483
rect 270417 8449 270451 8483
rect 270693 8449 270727 8483
rect 22017 8381 22051 8415
rect 22661 8381 22695 8415
rect 24409 8381 24443 8415
rect 24685 8381 24719 8415
rect 33885 8381 33919 8415
rect 54493 8381 54527 8415
rect 56977 8381 57011 8415
rect 67005 8381 67039 8415
rect 76757 8381 76791 8415
rect 93041 8381 93075 8415
rect 96537 8381 96571 8415
rect 100677 8381 100711 8415
rect 100953 8381 100987 8415
rect 101965 8381 101999 8415
rect 121285 8381 121319 8415
rect 128645 8381 128679 8415
rect 129013 8381 129047 8415
rect 130209 8381 130243 8415
rect 130853 8381 130887 8415
rect 132693 8381 132727 8415
rect 156705 8381 156739 8415
rect 157809 8381 157843 8415
rect 159465 8381 159499 8415
rect 160017 8381 160051 8415
rect 161029 8381 161063 8415
rect 162685 8381 162719 8415
rect 163973 8381 164007 8415
rect 165353 8381 165387 8415
rect 167653 8381 167687 8415
rect 168665 8381 168699 8415
rect 168941 8381 168975 8415
rect 169953 8381 169987 8415
rect 187249 8381 187283 8415
rect 195253 8381 195287 8415
rect 197185 8381 197219 8415
rect 198197 8381 198231 8415
rect 202337 8381 202371 8415
rect 203165 8381 203199 8415
rect 233433 8381 233467 8415
rect 235089 8381 235123 8415
rect 256985 8381 257019 8415
rect 260941 8381 260975 8415
rect 261585 8381 261619 8415
rect 266553 8381 266587 8415
rect 267473 8381 267507 8415
rect 267841 8381 267875 8415
rect 269497 8381 269531 8415
rect 23029 8313 23063 8347
rect 65533 8313 65567 8347
rect 66269 8313 66303 8347
rect 158177 8313 158211 8347
rect 161397 8313 161431 8347
rect 190561 8313 190595 8347
rect 191297 8313 191331 8347
rect 193321 8313 193355 8347
rect 194057 8313 194091 8347
rect 196265 8313 196299 8347
rect 199209 8313 199243 8347
rect 199945 8313 199979 8347
rect 200773 8313 200807 8347
rect 201509 8313 201543 8347
rect 264437 8313 264471 8347
rect 25053 8245 25087 8279
rect 61025 8245 61059 8279
rect 90097 8245 90131 8279
rect 129381 8245 129415 8279
rect 133061 8245 133095 8279
rect 157073 8245 157107 8279
rect 160385 8245 160419 8279
rect 166641 8245 166675 8279
rect 263057 8245 263091 8279
rect 268485 8245 268519 8279
rect 269957 8245 269991 8279
rect 67281 8041 67315 8075
rect 100861 8041 100895 8075
rect 129289 8041 129323 8075
rect 132969 8041 133003 8075
rect 157257 8041 157291 8075
rect 158729 8041 158763 8075
rect 160201 8041 160235 8075
rect 160937 8041 160971 8075
rect 161673 8041 161707 8075
rect 162409 8041 162443 8075
rect 163881 8041 163915 8075
rect 164617 8041 164651 8075
rect 166089 8041 166123 8075
rect 259561 8041 259595 8075
rect 260849 8041 260883 8075
rect 261769 8041 261803 8075
rect 262505 8041 262539 8075
rect 263333 8041 263367 8075
rect 264989 8041 265023 8075
rect 267473 8041 267507 8075
rect 268853 8041 268887 8075
rect 21925 7973 21959 8007
rect 22937 7973 22971 8007
rect 23673 7973 23707 8007
rect 25237 7973 25271 8007
rect 109877 7973 109911 8007
rect 168205 7973 168239 8007
rect 169217 7973 169251 8007
rect 270233 7973 270267 8007
rect 32873 7905 32907 7939
rect 66913 7905 66947 7939
rect 67741 7905 67775 7939
rect 100493 7905 100527 7939
rect 134257 7905 134291 7939
rect 168849 7905 168883 7939
rect 267105 7905 267139 7939
rect 21741 7837 21775 7871
rect 22753 7837 22787 7871
rect 23489 7837 23523 7871
rect 25053 7837 25087 7871
rect 67097 7837 67131 7871
rect 89545 7837 89579 7871
rect 100677 7837 100711 7871
rect 109325 7837 109359 7871
rect 110061 7837 110095 7871
rect 114937 7837 114971 7871
rect 116133 7837 116167 7871
rect 129105 7837 129139 7871
rect 132785 7837 132819 7871
rect 157073 7837 157107 7871
rect 158545 7837 158579 7871
rect 159281 7837 159315 7871
rect 160017 7837 160051 7871
rect 160753 7837 160787 7871
rect 161489 7837 161523 7871
rect 162225 7837 162259 7871
rect 163697 7837 163731 7871
rect 164433 7837 164467 7871
rect 165169 7837 165203 7871
rect 165905 7837 165939 7871
rect 166629 7837 166663 7871
rect 167837 7837 167871 7871
rect 168021 7837 168055 7871
rect 169033 7837 169067 7871
rect 202981 7837 203015 7871
rect 225521 7837 225555 7871
rect 234721 7837 234755 7871
rect 260389 7837 260423 7871
rect 261033 7837 261067 7871
rect 261585 7837 261619 7871
rect 262321 7837 262355 7871
rect 263149 7837 263183 7871
rect 263977 7837 264011 7871
rect 264161 7837 264195 7871
rect 264345 7837 264379 7871
rect 264805 7837 264839 7871
rect 265633 7837 265667 7871
rect 265725 7837 265759 7871
rect 267289 7837 267323 7871
rect 268025 7837 268059 7871
rect 268117 7837 268151 7871
rect 268761 7837 268795 7871
rect 269681 7837 269715 7871
rect 269865 7837 269899 7871
rect 270101 7837 270135 7871
rect 270785 7837 270819 7871
rect 115305 7769 115339 7803
rect 116225 7769 116259 7803
rect 224417 7769 224451 7803
rect 259929 7769 259963 7803
rect 269957 7769 269991 7803
rect 89729 7701 89763 7735
rect 97825 7701 97859 7735
rect 109141 7701 109175 7735
rect 115121 7701 115155 7735
rect 115213 7701 115247 7735
rect 115489 7701 115523 7735
rect 159465 7701 159499 7735
rect 165353 7701 165387 7735
rect 166825 7701 166859 7735
rect 224509 7701 224543 7735
rect 225705 7701 225739 7735
rect 234905 7701 234939 7735
rect 235825 7701 235859 7735
rect 260205 7701 260239 7735
rect 265909 7701 265943 7735
rect 268301 7701 268335 7735
rect 269221 7701 269255 7735
rect 270877 7701 270911 7735
rect 76389 7497 76423 7531
rect 101321 7497 101355 7531
rect 110613 7497 110647 7531
rect 111533 7497 111567 7531
rect 115305 7497 115339 7531
rect 115397 7497 115431 7531
rect 117513 7497 117547 7531
rect 119905 7497 119939 7531
rect 163145 7497 163179 7531
rect 166917 7497 166951 7531
rect 168573 7497 168607 7531
rect 221473 7497 221507 7531
rect 261493 7497 261527 7531
rect 262137 7497 262171 7531
rect 262781 7497 262815 7531
rect 263425 7497 263459 7531
rect 264345 7497 264379 7531
rect 265449 7497 265483 7531
rect 266185 7497 266219 7531
rect 270877 7497 270911 7531
rect 162317 7429 162351 7463
rect 226349 7429 226383 7463
rect 252109 7429 252143 7463
rect 253121 7429 253155 7463
rect 269865 7429 269899 7463
rect 76573 7361 76607 7395
rect 78781 7361 78815 7395
rect 94973 7361 95007 7395
rect 95847 7361 95881 7395
rect 97365 7361 97399 7395
rect 97549 7361 97583 7395
rect 98653 7361 98687 7395
rect 99481 7361 99515 7395
rect 100125 7361 100159 7395
rect 101505 7361 101539 7395
rect 107117 7361 107151 7395
rect 108405 7361 108439 7395
rect 109049 7361 109083 7395
rect 109785 7361 109819 7395
rect 110797 7361 110831 7395
rect 111257 7361 111291 7395
rect 111901 7361 111935 7395
rect 112085 7361 112119 7395
rect 112821 7361 112855 7395
rect 113097 7361 113131 7395
rect 115029 7361 115063 7395
rect 116317 7361 116351 7395
rect 117421 7361 117455 7395
rect 118065 7361 118099 7395
rect 120089 7361 120123 7395
rect 151829 7361 151863 7395
rect 152749 7361 152783 7395
rect 162501 7361 162535 7395
rect 162961 7361 162995 7395
rect 166733 7361 166767 7395
rect 168757 7361 168791 7395
rect 213469 7361 213503 7395
rect 218529 7361 218563 7395
rect 221657 7361 221691 7395
rect 223957 7361 223991 7395
rect 224601 7361 224635 7395
rect 225981 7361 226015 7395
rect 250177 7361 250211 7395
rect 251005 7361 251039 7395
rect 251925 7361 251959 7395
rect 252845 7361 252879 7395
rect 252937 7361 252971 7395
rect 260389 7361 260423 7395
rect 260849 7361 260883 7395
rect 261677 7361 261711 7395
rect 262321 7361 262355 7395
rect 262965 7361 262999 7395
rect 263609 7361 263643 7395
rect 264161 7361 264195 7395
rect 265265 7361 265299 7395
rect 266007 7361 266041 7395
rect 267289 7361 267323 7395
rect 268117 7361 268151 7395
rect 269577 7361 269611 7395
rect 269682 7361 269716 7395
rect 269957 7361 269991 7395
rect 270095 7361 270129 7395
rect 270785 7361 270819 7395
rect 94789 7293 94823 7327
rect 95709 7293 95743 7327
rect 95985 7293 96019 7327
rect 112959 7293 112993 7327
rect 115489 7293 115523 7327
rect 152013 7293 152047 7327
rect 213653 7293 213687 7327
rect 225061 7293 225095 7327
rect 249993 7293 250027 7327
rect 250821 7293 250855 7327
rect 251189 7293 251223 7327
rect 251741 7293 251775 7327
rect 261217 7293 261251 7327
rect 267105 7293 267139 7327
rect 267933 7293 267967 7327
rect 78965 7225 78999 7259
rect 95433 7225 95467 7259
rect 106933 7225 106967 7259
rect 108865 7225 108899 7259
rect 112545 7225 112579 7259
rect 115673 7225 115707 7259
rect 218713 7225 218747 7259
rect 223773 7225 223807 7259
rect 260665 7225 260699 7259
rect 96629 7157 96663 7191
rect 97457 7157 97491 7191
rect 97733 7157 97767 7191
rect 98469 7157 98503 7191
rect 99297 7157 99331 7191
rect 99941 7157 99975 7191
rect 108221 7157 108255 7191
rect 109601 7157 109635 7191
rect 111073 7157 111107 7191
rect 113741 7157 113775 7191
rect 116593 7157 116627 7191
rect 118157 7157 118191 7191
rect 152933 7157 152967 7191
rect 250361 7157 250395 7191
rect 260205 7157 260239 7191
rect 267473 7157 267507 7191
rect 268301 7157 268335 7191
rect 270233 7157 270267 7191
rect 97641 6953 97675 6987
rect 98285 6953 98319 6987
rect 100493 6953 100527 6987
rect 108773 6953 108807 6987
rect 108957 6953 108991 6987
rect 110337 6953 110371 6987
rect 151093 6953 151127 6987
rect 151829 6953 151863 6987
rect 153393 6953 153427 6987
rect 269221 6953 269255 6987
rect 106197 6885 106231 6919
rect 110613 6885 110647 6919
rect 112177 6885 112211 6919
rect 116685 6885 116719 6919
rect 190193 6885 190227 6919
rect 223497 6885 223531 6919
rect 261769 6885 261803 6919
rect 97549 6817 97583 6851
rect 109693 6817 109727 6851
rect 113741 6817 113775 6851
rect 114569 6817 114603 6851
rect 116317 6817 116351 6851
rect 216873 6817 216907 6851
rect 226993 6817 227027 6851
rect 263609 6817 263643 6851
rect 268577 6817 268611 6851
rect 270509 6817 270543 6851
rect 96169 6749 96203 6783
rect 96905 6749 96939 6783
rect 97457 6749 97491 6783
rect 98285 6749 98319 6783
rect 98469 6749 98503 6783
rect 99849 6749 99883 6783
rect 100403 6749 100437 6783
rect 101321 6749 101355 6783
rect 102057 6749 102091 6783
rect 102701 6749 102735 6783
rect 106381 6749 106415 6783
rect 107485 6749 107519 6783
rect 108129 6749 108163 6783
rect 108589 6749 108623 6783
rect 108681 6749 108715 6783
rect 110245 6749 110279 6783
rect 110429 6749 110463 6783
rect 111257 6749 111291 6783
rect 112361 6749 112395 6783
rect 113005 6749 113039 6783
rect 116041 6749 116075 6783
rect 151001 6749 151035 6783
rect 151369 6749 151403 6783
rect 152197 6749 152231 6783
rect 153577 6749 153611 6783
rect 190377 6749 190411 6783
rect 213193 6749 213227 6783
rect 216597 6749 216631 6783
rect 217333 6749 217367 6783
rect 223313 6749 223347 6783
rect 225613 6749 225647 6783
rect 226717 6749 226751 6783
rect 238401 6749 238435 6783
rect 248705 6749 248739 6783
rect 249349 6749 249383 6783
rect 251373 6749 251407 6783
rect 251465 6749 251499 6783
rect 253029 6749 253063 6783
rect 253305 6749 253339 6783
rect 256617 6749 256651 6783
rect 261033 6749 261067 6783
rect 261953 6749 261987 6783
rect 262413 6749 262447 6783
rect 262781 6749 262815 6783
rect 263241 6749 263275 6783
rect 263701 6749 263735 6783
rect 264437 6749 264471 6783
rect 265909 6749 265943 6783
rect 266829 6749 266863 6783
rect 266921 6749 266955 6783
rect 268025 6749 268059 6783
rect 269221 6749 269255 6783
rect 269865 6749 269899 6783
rect 270049 6749 270083 6783
rect 270601 6749 270635 6783
rect 109509 6681 109543 6715
rect 113925 6681 113959 6715
rect 116526 6681 116560 6715
rect 117421 6681 117455 6715
rect 118341 6681 118375 6715
rect 152473 6681 152507 6715
rect 213837 6681 213871 6715
rect 216045 6681 216079 6715
rect 216321 6681 216355 6715
rect 224141 6681 224175 6715
rect 239045 6681 239079 6715
rect 255697 6681 255731 6715
rect 264897 6681 264931 6715
rect 95985 6613 96019 6647
rect 96721 6613 96755 6647
rect 97825 6613 97859 6647
rect 98653 6613 98687 6647
rect 99665 6613 99699 6647
rect 101137 6613 101171 6647
rect 101873 6613 101907 6647
rect 102517 6613 102551 6647
rect 107301 6613 107335 6647
rect 107945 6613 107979 6647
rect 111073 6613 111107 6647
rect 112821 6613 112855 6647
rect 116409 6613 116443 6647
rect 117513 6613 117547 6647
rect 118433 6613 118467 6647
rect 151553 6613 151587 6647
rect 216505 6613 216539 6647
rect 216689 6613 216723 6647
rect 217425 6613 217459 6647
rect 224233 6613 224267 6647
rect 225705 6613 225739 6647
rect 248521 6613 248555 6647
rect 249165 6613 249199 6647
rect 251649 6613 251683 6647
rect 255789 6613 255823 6647
rect 256433 6613 256467 6647
rect 262229 6613 262263 6647
rect 263057 6613 263091 6647
rect 263793 6613 263827 6647
rect 266093 6613 266127 6647
rect 267105 6613 267139 6647
rect 98745 6409 98779 6443
rect 100033 6409 100067 6443
rect 102333 6409 102367 6443
rect 108129 6409 108163 6443
rect 112821 6409 112855 6443
rect 118157 6409 118191 6443
rect 118985 6409 119019 6443
rect 119169 6409 119203 6443
rect 151369 6409 151403 6443
rect 188813 6409 188847 6443
rect 189365 6409 189399 6443
rect 189457 6409 189491 6443
rect 189733 6409 189767 6443
rect 216413 6409 216447 6443
rect 224969 6409 225003 6443
rect 249349 6409 249383 6443
rect 253121 6409 253155 6443
rect 254685 6409 254719 6443
rect 255789 6409 255823 6443
rect 256709 6409 256743 6443
rect 95525 6341 95559 6375
rect 102885 6341 102919 6375
rect 107117 6341 107151 6375
rect 109785 6341 109819 6375
rect 111441 6341 111475 6375
rect 141525 6341 141559 6375
rect 168757 6341 168791 6375
rect 169953 6341 169987 6375
rect 189181 6341 189215 6375
rect 190009 6341 190043 6375
rect 256249 6341 256283 6375
rect 262045 6341 262079 6375
rect 52929 6273 52963 6307
rect 91937 6273 91971 6307
rect 92949 6273 92983 6307
rect 94881 6273 94915 6307
rect 97917 6273 97951 6307
rect 98377 6273 98411 6307
rect 99481 6273 99515 6307
rect 99849 6273 99883 6307
rect 100677 6273 100711 6307
rect 101137 6273 101171 6307
rect 101321 6273 101355 6307
rect 101965 6273 101999 6307
rect 102057 6273 102091 6307
rect 103069 6273 103103 6307
rect 104633 6273 104667 6307
rect 105645 6273 105679 6307
rect 106289 6273 106323 6307
rect 107761 6273 107795 6307
rect 108589 6273 108623 6307
rect 109601 6273 109635 6307
rect 112085 6273 112119 6307
rect 113005 6273 113039 6307
rect 113465 6273 113499 6307
rect 113741 6273 113775 6307
rect 115029 6273 115063 6307
rect 115949 6273 115983 6307
rect 117605 6273 117639 6307
rect 118801 6273 118835 6307
rect 118893 6273 118927 6307
rect 135361 6273 135395 6307
rect 137017 6273 137051 6307
rect 140513 6273 140547 6307
rect 142261 6273 142295 6307
rect 150265 6273 150299 6307
rect 150817 6273 150851 6307
rect 151829 6273 151863 6307
rect 152841 6273 152875 6307
rect 153853 6273 153887 6307
rect 154865 6273 154899 6307
rect 156153 6273 156187 6307
rect 168113 6273 168147 6307
rect 168389 6273 168423 6307
rect 169585 6273 169619 6307
rect 189549 6273 189583 6307
rect 208225 6273 208259 6307
rect 209145 6273 209179 6307
rect 209283 6273 209317 6307
rect 213101 6273 213135 6307
rect 216137 6273 216171 6307
rect 217149 6273 217183 6307
rect 217885 6273 217919 6307
rect 217977 6273 218011 6307
rect 218069 6273 218103 6307
rect 218805 6273 218839 6307
rect 221657 6273 221691 6307
rect 221749 6273 221783 6307
rect 221841 6273 221875 6307
rect 224601 6273 224635 6307
rect 226165 6273 226199 6307
rect 226441 6273 226475 6307
rect 248153 6273 248187 6307
rect 248889 6273 248923 6307
rect 249165 6273 249199 6307
rect 249993 6273 250027 6307
rect 250637 6273 250671 6307
rect 252845 6273 252879 6307
rect 252937 6273 252971 6307
rect 254869 6273 254903 6307
rect 255329 6273 255363 6307
rect 255605 6273 255639 6307
rect 256525 6273 256559 6307
rect 257353 6273 257387 6307
rect 260113 6273 260147 6307
rect 260941 6273 260975 6307
rect 261677 6273 261711 6307
rect 262965 6273 262999 6307
rect 264253 6273 264287 6307
rect 265449 6273 265483 6307
rect 266645 6273 266679 6307
rect 267197 6273 267231 6307
rect 267841 6273 267875 6307
rect 269405 6273 269439 6307
rect 270693 6273 270727 6307
rect 53113 6205 53147 6239
rect 91753 6205 91787 6239
rect 92673 6205 92707 6239
rect 92811 6205 92845 6239
rect 93593 6205 93627 6239
rect 95341 6205 95375 6239
rect 96905 6205 96939 6239
rect 98469 6205 98503 6239
rect 107853 6205 107887 6239
rect 108681 6205 108715 6239
rect 115213 6205 115247 6239
rect 115673 6205 115707 6239
rect 116087 6205 116121 6239
rect 116235 6205 116269 6239
rect 117881 6205 117915 6239
rect 118617 6205 118651 6239
rect 135545 6205 135579 6239
rect 137201 6205 137235 6239
rect 140789 6205 140823 6239
rect 151093 6205 151127 6239
rect 152105 6205 152139 6239
rect 153025 6205 153059 6239
rect 168665 6205 168699 6239
rect 168874 6205 168908 6239
rect 208409 6205 208443 6239
rect 209421 6205 209455 6239
rect 213285 6205 213319 6239
rect 216505 6205 216539 6239
rect 216622 6205 216656 6239
rect 218989 6205 219023 6239
rect 219725 6205 219759 6239
rect 219863 6205 219897 6239
rect 220001 6205 220035 6239
rect 222761 6205 222795 6239
rect 222945 6205 222979 6239
rect 225245 6205 225279 6239
rect 225429 6205 225463 6239
rect 226282 6205 226316 6239
rect 248981 6205 249015 6239
rect 255513 6205 255547 6239
rect 256433 6205 256467 6239
rect 259929 6205 259963 6239
rect 260757 6205 260791 6239
rect 263241 6205 263275 6239
rect 264529 6205 264563 6239
rect 265725 6205 265759 6239
rect 268393 6205 268427 6239
rect 269681 6205 269715 6239
rect 270509 6205 270543 6239
rect 53757 6137 53791 6171
rect 92397 6137 92431 6171
rect 101505 6137 101539 6171
rect 104449 6137 104483 6171
rect 107301 6137 107335 6171
rect 114017 6137 114051 6171
rect 152381 6137 152415 6171
rect 155969 6137 156003 6171
rect 167745 6137 167779 6171
rect 169033 6137 169067 6171
rect 208869 6137 208903 6171
rect 216781 6137 216815 6171
rect 219449 6137 219483 6171
rect 225889 6137 225923 6171
rect 94697 6069 94731 6103
rect 97733 6069 97767 6103
rect 98377 6069 98411 6103
rect 99573 6069 99607 6103
rect 100493 6069 100527 6103
rect 101137 6069 101171 6103
rect 101965 6069 101999 6103
rect 103713 6069 103747 6103
rect 105461 6069 105495 6103
rect 106105 6069 106139 6103
rect 107945 6069 107979 6103
rect 108773 6069 108807 6103
rect 108957 6069 108991 6103
rect 111901 6069 111935 6103
rect 113557 6069 113591 6103
rect 116869 6069 116903 6103
rect 117973 6069 118007 6103
rect 141617 6069 141651 6103
rect 142353 6069 142387 6103
rect 150081 6069 150115 6103
rect 150909 6069 150943 6103
rect 151921 6069 151955 6103
rect 153945 6069 153979 6103
rect 154681 6069 154715 6103
rect 210065 6069 210099 6103
rect 215861 6069 215895 6103
rect 218253 6069 218287 6103
rect 220645 6069 220679 6103
rect 222025 6069 222059 6103
rect 227085 6069 227119 6103
rect 247969 6069 248003 6103
rect 248889 6069 248923 6103
rect 249809 6069 249843 6103
rect 250453 6069 250487 6103
rect 255605 6069 255639 6103
rect 256433 6069 256467 6103
rect 257169 6069 257203 6103
rect 260297 6069 260331 6103
rect 261125 6069 261159 6103
rect 270877 6069 270911 6103
rect 46673 5865 46707 5899
rect 95985 5865 96019 5899
rect 96169 5865 96203 5899
rect 96721 5865 96755 5899
rect 97089 5865 97123 5899
rect 100125 5865 100159 5899
rect 100953 5865 100987 5899
rect 101873 5865 101907 5899
rect 104357 5865 104391 5899
rect 107209 5865 107243 5899
rect 113465 5865 113499 5899
rect 114293 5865 114327 5899
rect 116593 5865 116627 5899
rect 116777 5865 116811 5899
rect 148333 5865 148367 5899
rect 150081 5865 150115 5899
rect 155969 5865 156003 5899
rect 157717 5865 157751 5899
rect 169217 5865 169251 5899
rect 217425 5865 217459 5899
rect 224969 5865 225003 5899
rect 225705 5865 225739 5899
rect 248061 5865 248095 5899
rect 248245 5865 248279 5899
rect 248889 5865 248923 5899
rect 249717 5865 249751 5899
rect 259377 5865 259411 5899
rect 263149 5865 263183 5899
rect 265265 5865 265299 5899
rect 95157 5797 95191 5831
rect 100401 5797 100435 5831
rect 101321 5797 101355 5831
rect 102241 5797 102275 5831
rect 102977 5797 103011 5831
rect 107669 5797 107703 5831
rect 108405 5797 108439 5831
rect 112453 5797 112487 5831
rect 114661 5797 114695 5831
rect 138949 5797 138983 5831
rect 148793 5797 148827 5831
rect 150541 5797 150575 5831
rect 188813 5797 188847 5831
rect 190101 5797 190135 5831
rect 249165 5797 249199 5831
rect 250545 5797 250579 5831
rect 254593 5797 254627 5831
rect 270509 5797 270543 5831
rect 47593 5729 47627 5763
rect 97549 5729 97583 5763
rect 97733 5729 97767 5763
rect 98469 5729 98503 5763
rect 101045 5729 101079 5763
rect 101965 5729 101999 5763
rect 109049 5729 109083 5763
rect 109233 5729 109267 5763
rect 114385 5729 114419 5763
rect 115397 5729 115431 5763
rect 115581 5729 115615 5763
rect 116501 5729 116535 5763
rect 117329 5729 117363 5763
rect 120114 5729 120148 5763
rect 140053 5729 140087 5763
rect 140789 5729 140823 5763
rect 148517 5729 148551 5763
rect 151645 5729 151679 5763
rect 153761 5729 153795 5763
rect 154405 5729 154439 5763
rect 154681 5729 154715 5763
rect 154819 5729 154853 5763
rect 189825 5729 189859 5763
rect 190377 5729 190411 5763
rect 216413 5729 216447 5763
rect 216781 5729 216815 5763
rect 217057 5729 217091 5763
rect 220553 5729 220587 5763
rect 220829 5729 220863 5763
rect 223129 5729 223163 5763
rect 223773 5729 223807 5763
rect 224049 5729 224083 5763
rect 224187 5729 224221 5763
rect 247877 5729 247911 5763
rect 248889 5729 248923 5763
rect 249809 5729 249843 5763
rect 255053 5729 255087 5763
rect 259377 5729 259411 5763
rect 269865 5729 269899 5763
rect 45661 5661 45695 5695
rect 46121 5661 46155 5695
rect 48145 5661 48179 5695
rect 51549 5661 51583 5695
rect 52285 5661 52319 5695
rect 52377 5661 52411 5695
rect 94697 5661 94731 5695
rect 95341 5661 95375 5695
rect 95801 5661 95835 5695
rect 95985 5661 96019 5695
rect 96721 5661 96755 5695
rect 96905 5661 96939 5695
rect 99849 5661 99883 5695
rect 100217 5661 100251 5695
rect 100953 5661 100987 5695
rect 101873 5661 101907 5695
rect 103621 5661 103655 5695
rect 104541 5661 104575 5695
rect 105185 5661 105219 5695
rect 105829 5661 105863 5695
rect 106473 5661 106507 5695
rect 107117 5661 107151 5695
rect 107393 5661 107427 5695
rect 112269 5661 112303 5695
rect 113465 5661 113499 5695
rect 113649 5661 113683 5695
rect 114293 5661 114327 5695
rect 115121 5661 115155 5695
rect 115489 5661 115523 5695
rect 116409 5661 116443 5695
rect 119169 5661 119203 5695
rect 119629 5661 119663 5695
rect 121009 5661 121043 5695
rect 121561 5661 121595 5695
rect 121929 5661 121963 5695
rect 127725 5661 127759 5695
rect 128093 5661 128127 5695
rect 136097 5661 136131 5695
rect 139133 5661 139167 5695
rect 139777 5661 139811 5695
rect 140605 5661 140639 5695
rect 142445 5661 142479 5695
rect 143273 5661 143307 5695
rect 144837 5661 144871 5695
rect 145481 5661 145515 5695
rect 146493 5661 146527 5695
rect 146769 5661 146803 5695
rect 148241 5661 148275 5695
rect 149529 5661 149563 5695
rect 149989 5661 150023 5695
rect 150265 5661 150299 5695
rect 151001 5661 151035 5695
rect 151185 5661 151219 5695
rect 151921 5661 151955 5695
rect 152059 5661 152093 5695
rect 152197 5661 152231 5695
rect 153945 5661 153979 5695
rect 154957 5661 154991 5695
rect 156705 5661 156739 5695
rect 168021 5661 168055 5695
rect 168849 5661 168883 5695
rect 169217 5661 169251 5695
rect 169861 5661 169895 5695
rect 189457 5661 189491 5695
rect 207305 5661 207339 5695
rect 212825 5661 212859 5695
rect 213285 5661 213319 5695
rect 213377 5661 213411 5695
rect 213653 5661 213687 5695
rect 215401 5661 215435 5695
rect 218253 5661 218287 5695
rect 218345 5661 218379 5695
rect 218529 5661 218563 5695
rect 220369 5661 220403 5695
rect 223313 5661 223347 5695
rect 224325 5661 224359 5695
rect 225521 5661 225555 5695
rect 247325 5661 247359 5695
rect 248061 5661 248095 5695
rect 248981 5661 249015 5695
rect 249901 5661 249935 5695
rect 250729 5661 250763 5695
rect 253857 5661 253891 5695
rect 255329 5661 255363 5695
rect 256433 5661 256467 5695
rect 256709 5661 256743 5695
rect 257905 5661 257939 5695
rect 259285 5661 259319 5695
rect 259561 5661 259595 5695
rect 260389 5661 260423 5695
rect 261677 5661 261711 5695
rect 262873 5661 262907 5695
rect 262965 5661 262999 5695
rect 263793 5661 263827 5695
rect 264345 5661 264379 5695
rect 264897 5661 264931 5695
rect 265081 5661 265115 5695
rect 265909 5661 265943 5695
rect 266921 5661 266955 5695
rect 268393 5661 268427 5695
rect 269589 5661 269623 5695
rect 269681 5661 269715 5695
rect 270325 5661 270359 5695
rect 156797 5627 156831 5661
rect 45753 5593 45787 5627
rect 47317 5593 47351 5627
rect 52745 5593 52779 5627
rect 102793 5593 102827 5627
rect 108221 5593 108255 5627
rect 110889 5593 110923 5627
rect 111441 5593 111475 5627
rect 117513 5593 117547 5627
rect 119905 5593 119939 5627
rect 119997 5593 120031 5627
rect 132877 5593 132911 5627
rect 133245 5593 133279 5627
rect 144101 5593 144135 5627
rect 145757 5593 145791 5627
rect 155601 5593 155635 5627
rect 156383 5593 156417 5627
rect 157165 5593 157199 5627
rect 157533 5593 157567 5627
rect 169953 5593 169987 5627
rect 189942 5593 189976 5627
rect 207489 5593 207523 5627
rect 209145 5593 209179 5627
rect 216137 5593 216171 5627
rect 217266 5593 217300 5627
rect 218897 5593 218931 5627
rect 247785 5593 247819 5627
rect 248705 5593 248739 5627
rect 249625 5593 249659 5627
rect 254409 5593 254443 5627
rect 260757 5593 260791 5627
rect 262045 5593 262079 5627
rect 267289 5593 267323 5627
rect 268761 5593 268795 5627
rect 45385 5525 45419 5559
rect 46489 5525 46523 5559
rect 48329 5525 48363 5559
rect 51181 5525 51215 5559
rect 52009 5525 52043 5559
rect 53113 5525 53147 5559
rect 53297 5525 53331 5559
rect 94513 5525 94547 5559
rect 103437 5525 103471 5559
rect 105001 5525 105035 5559
rect 105645 5525 105679 5559
rect 106289 5525 106323 5559
rect 111533 5525 111567 5559
rect 113833 5525 113867 5559
rect 115765 5525 115799 5559
rect 120273 5525 120307 5559
rect 120825 5525 120859 5559
rect 136281 5525 136315 5559
rect 143089 5525 143123 5559
rect 149345 5525 149379 5559
rect 152841 5525 152875 5559
rect 168205 5525 168239 5559
rect 169401 5525 169435 5559
rect 189733 5525 189767 5559
rect 215217 5525 215251 5559
rect 217149 5525 217183 5559
rect 247141 5525 247175 5559
rect 250085 5525 250119 5559
rect 253673 5525 253707 5559
rect 257721 5525 257755 5559
rect 259745 5525 259779 5559
rect 265725 5525 265759 5559
rect 35541 5321 35575 5355
rect 99849 5321 99883 5355
rect 100861 5321 100895 5355
rect 101873 5321 101907 5355
rect 102701 5321 102735 5355
rect 108957 5321 108991 5355
rect 113189 5321 113223 5355
rect 116041 5321 116075 5355
rect 143733 5321 143767 5355
rect 206937 5321 206971 5355
rect 247233 5321 247267 5355
rect 248153 5321 248187 5355
rect 262505 5321 262539 5355
rect 263425 5321 263459 5355
rect 265081 5321 265115 5355
rect 266829 5321 266863 5355
rect 267749 5321 267783 5355
rect 268577 5321 268611 5355
rect 269681 5321 269715 5355
rect 35817 5253 35851 5287
rect 36277 5253 36311 5287
rect 36645 5253 36679 5287
rect 45845 5253 45879 5287
rect 46121 5253 46155 5287
rect 46949 5253 46983 5287
rect 50997 5253 51031 5287
rect 52101 5253 52135 5287
rect 110981 5253 111015 5287
rect 112637 5253 112671 5287
rect 153301 5253 153335 5287
rect 156153 5253 156187 5287
rect 216505 5253 216539 5287
rect 220369 5253 220403 5287
rect 223129 5253 223163 5287
rect 225429 5253 225463 5287
rect 246773 5253 246807 5287
rect 247693 5253 247727 5287
rect 248889 5253 248923 5287
rect 251097 5253 251131 5287
rect 254225 5253 254259 5287
rect 255329 5253 255363 5287
rect 256985 5253 257019 5287
rect 265817 5253 265851 5287
rect 270509 5253 270543 5287
rect 35909 5185 35943 5219
rect 46213 5185 46247 5219
rect 46581 5185 46615 5219
rect 50445 5185 50479 5219
rect 51273 5185 51307 5219
rect 51365 5185 51399 5219
rect 51733 5185 51767 5219
rect 52929 5185 52963 5219
rect 53573 5185 53607 5219
rect 93593 5185 93627 5219
rect 94329 5185 94363 5219
rect 98469 5185 98503 5219
rect 99297 5185 99331 5219
rect 100309 5185 100343 5219
rect 101321 5185 101355 5219
rect 101689 5185 101723 5219
rect 102333 5185 102367 5219
rect 103345 5185 103379 5219
rect 105001 5185 105035 5219
rect 105737 5185 105771 5219
rect 107025 5185 107059 5219
rect 108589 5185 108623 5219
rect 108681 5185 108715 5219
rect 109785 5185 109819 5219
rect 110153 5185 110187 5219
rect 110797 5185 110831 5219
rect 113373 5185 113407 5219
rect 113833 5185 113867 5219
rect 114753 5185 114787 5219
rect 114845 5185 114879 5219
rect 115857 5185 115891 5219
rect 116225 5185 116259 5219
rect 116501 5185 116535 5219
rect 116961 5185 116995 5219
rect 118801 5185 118835 5219
rect 119905 5185 119939 5219
rect 120641 5185 120675 5219
rect 121009 5185 121043 5219
rect 121837 5185 121871 5219
rect 122481 5185 122515 5219
rect 137477 5185 137511 5219
rect 138765 5185 138799 5219
rect 139409 5185 139443 5219
rect 140513 5185 140547 5219
rect 142169 5185 142203 5219
rect 143181 5185 143215 5219
rect 144377 5185 144411 5219
rect 145021 5185 145055 5219
rect 145665 5185 145699 5219
rect 148241 5185 148275 5219
rect 148517 5185 148551 5219
rect 149718 5185 149752 5219
rect 150817 5185 150851 5219
rect 151737 5185 151771 5219
rect 155969 5185 156003 5219
rect 169953 5185 169987 5219
rect 206569 5185 206603 5219
rect 206661 5185 206695 5219
rect 206753 5185 206787 5219
rect 207489 5185 207523 5219
rect 209881 5185 209915 5219
rect 213193 5185 213227 5219
rect 213469 5185 213503 5219
rect 214389 5185 214423 5219
rect 214506 5185 214540 5219
rect 215861 5185 215895 5219
rect 215953 5185 215987 5219
rect 216321 5185 216355 5219
rect 217149 5185 217183 5219
rect 217885 5185 217919 5219
rect 218069 5185 218103 5219
rect 218805 5185 218839 5219
rect 219081 5185 219115 5219
rect 220185 5185 220219 5219
rect 246129 5185 246163 5219
rect 247049 5185 247083 5219
rect 247877 5185 247911 5219
rect 247969 5185 248003 5219
rect 248705 5185 248739 5219
rect 251925 5185 251959 5219
rect 253305 5185 253339 5219
rect 254501 5185 254535 5219
rect 255145 5185 255179 5219
rect 257445 5185 257479 5219
rect 257721 5185 257755 5219
rect 259837 5185 259871 5219
rect 261033 5185 261067 5219
rect 262321 5185 262355 5219
rect 263609 5185 263643 5219
rect 264621 5185 264655 5219
rect 265265 5185 265299 5219
rect 266553 5185 266587 5219
rect 266645 5185 266679 5219
rect 267473 5185 267507 5219
rect 267565 5185 267599 5219
rect 268393 5185 268427 5219
rect 269313 5185 269347 5219
rect 269497 5185 269531 5219
rect 270325 5185 270359 5219
rect 94513 5117 94547 5151
rect 96169 5117 96203 5151
rect 96629 5117 96663 5151
rect 96813 5117 96847 5151
rect 99573 5117 99607 5151
rect 100585 5117 100619 5151
rect 102425 5117 102459 5151
rect 105277 5117 105311 5151
rect 107301 5117 107335 5151
rect 113925 5117 113959 5151
rect 117145 5117 117179 5151
rect 137753 5117 137787 5151
rect 139685 5117 139719 5151
rect 140789 5117 140823 5151
rect 142445 5117 142479 5151
rect 143457 5117 143491 5151
rect 145849 5117 145883 5151
rect 146401 5117 146435 5151
rect 149989 5117 150023 5151
rect 151001 5117 151035 5151
rect 151875 5117 151909 5151
rect 152013 5117 152047 5151
rect 153117 5117 153151 5151
rect 154773 5117 154807 5151
rect 157809 5117 157843 5151
rect 168113 5117 168147 5151
rect 168297 5117 168331 5151
rect 207673 5117 207707 5151
rect 208409 5117 208443 5151
rect 208547 5117 208581 5151
rect 208685 5117 208719 5151
rect 213653 5117 213687 5151
rect 214113 5117 214147 5151
rect 214665 5117 214699 5151
rect 218529 5117 218563 5151
rect 218943 5117 218977 5151
rect 220829 5117 220863 5151
rect 222945 5117 222979 5151
rect 223773 5117 223807 5151
rect 225245 5117 225279 5151
rect 227085 5117 227119 5151
rect 246865 5117 246899 5151
rect 250545 5117 250579 5151
rect 254409 5117 254443 5151
rect 257537 5117 257571 5151
rect 260113 5117 260147 5151
rect 261401 5117 261435 5151
rect 262137 5117 262171 5151
rect 268209 5117 268243 5151
rect 270141 5117 270175 5151
rect 47133 5049 47167 5083
rect 52285 5049 52319 5083
rect 53113 5049 53147 5083
rect 115121 5049 115155 5083
rect 121193 5049 121227 5083
rect 138029 5049 138063 5083
rect 138949 5049 138983 5083
rect 139961 5049 139995 5083
rect 144193 5049 144227 5083
rect 148793 5049 148827 5083
rect 150265 5049 150299 5083
rect 151461 5049 151495 5083
rect 208133 5049 208167 5083
rect 257905 5049 257939 5083
rect 264437 5049 264471 5083
rect 36829 4981 36863 5015
rect 93409 4981 93443 5015
rect 99665 4981 99699 5015
rect 100401 4981 100435 5015
rect 101413 4981 101447 5015
rect 102333 4981 102367 5015
rect 103161 4981 103195 5015
rect 104817 4981 104851 5015
rect 105829 4981 105863 5015
rect 108773 4981 108807 5015
rect 109877 4981 109911 5015
rect 110337 4981 110371 5015
rect 113833 4981 113867 5015
rect 114201 4981 114235 5015
rect 114753 4981 114787 5015
rect 116317 4981 116351 5015
rect 120089 4981 120123 5015
rect 120917 4981 120951 5015
rect 121653 4981 121687 5015
rect 122297 4981 122331 5015
rect 137569 4981 137603 5015
rect 139501 4981 139535 5015
rect 142261 4981 142295 5015
rect 142721 4981 142755 5015
rect 143457 4981 143491 5015
rect 144837 4981 144871 5015
rect 148333 4981 148367 5015
rect 149805 4981 149839 5015
rect 152657 4981 152691 5015
rect 209329 4981 209363 5015
rect 209973 4981 210007 5015
rect 215309 4981 215343 5015
rect 216965 4981 216999 5015
rect 219725 4981 219759 5015
rect 220093 4981 220127 5015
rect 245945 4981 245979 5015
rect 246957 4981 246991 5015
rect 247969 4981 248003 5015
rect 251189 4981 251223 5015
rect 251741 4981 251775 5015
rect 253121 4981 253155 5015
rect 254501 4981 254535 5015
rect 254685 4981 254719 5015
rect 257721 4981 257755 5015
rect 265909 4981 265943 5015
rect 37013 4777 37047 4811
rect 40969 4777 41003 4811
rect 42809 4777 42843 4811
rect 48053 4777 48087 4811
rect 100125 4777 100159 4811
rect 100861 4777 100895 4811
rect 101321 4777 101355 4811
rect 106013 4777 106047 4811
rect 107117 4777 107151 4811
rect 108129 4777 108163 4811
rect 112177 4777 112211 4811
rect 114109 4777 114143 4811
rect 114477 4777 114511 4811
rect 117697 4777 117731 4811
rect 120641 4777 120675 4811
rect 121653 4777 121687 4811
rect 121837 4777 121871 4811
rect 122757 4777 122791 4811
rect 143181 4777 143215 4811
rect 143641 4777 143675 4811
rect 151369 4777 151403 4811
rect 152381 4777 152415 4811
rect 165629 4777 165663 4811
rect 168113 4777 168147 4811
rect 222945 4777 222979 4811
rect 223865 4777 223899 4811
rect 224509 4777 224543 4811
rect 246957 4777 246991 4811
rect 251557 4777 251591 4811
rect 252569 4777 252603 4811
rect 258733 4777 258767 4811
rect 259193 4777 259227 4811
rect 264713 4777 264747 4811
rect 265357 4777 265391 4811
rect 266001 4777 266035 4811
rect 270693 4777 270727 4811
rect 92213 4709 92247 4743
rect 106473 4709 106507 4743
rect 108589 4709 108623 4743
rect 112821 4709 112855 4743
rect 113465 4709 113499 4743
rect 117789 4709 117823 4743
rect 117973 4709 118007 4743
rect 118709 4709 118743 4743
rect 119629 4709 119663 4743
rect 120825 4709 120859 4743
rect 141157 4709 141191 4743
rect 169125 4709 169159 4743
rect 212181 4709 212215 4743
rect 212549 4709 212583 4743
rect 244749 4709 244783 4743
rect 91569 4641 91603 4675
rect 92489 4641 92523 4675
rect 92627 4641 92661 4675
rect 94513 4641 94547 4675
rect 97457 4641 97491 4675
rect 97641 4641 97675 4675
rect 98653 4641 98687 4675
rect 102333 4641 102367 4675
rect 102517 4641 102551 4675
rect 106197 4641 106231 4675
rect 107301 4641 107335 4675
rect 109325 4641 109359 4675
rect 117881 4641 117915 4675
rect 121561 4641 121595 4675
rect 122757 4641 122791 4675
rect 138213 4641 138247 4675
rect 138857 4641 138891 4675
rect 139250 4641 139284 4675
rect 139409 4641 139443 4675
rect 140513 4641 140547 4675
rect 140697 4641 140731 4675
rect 141433 4641 141467 4675
rect 141709 4641 141743 4675
rect 143365 4641 143399 4675
rect 144469 4641 144503 4675
rect 144653 4641 144687 4675
rect 145113 4641 145147 4675
rect 145389 4641 145423 4675
rect 145665 4641 145699 4675
rect 148977 4641 149011 4675
rect 149161 4641 149195 4675
rect 149621 4641 149655 4675
rect 149897 4641 149931 4675
rect 150173 4641 150207 4675
rect 152565 4641 152599 4675
rect 153393 4641 153427 4675
rect 153577 4641 153611 4675
rect 154589 4641 154623 4675
rect 155877 4641 155911 4675
rect 156153 4641 156187 4675
rect 158545 4641 158579 4675
rect 159189 4641 159223 4675
rect 166457 4641 166491 4675
rect 166917 4641 166951 4675
rect 167331 4641 167365 4675
rect 206477 4641 206511 4675
rect 212825 4641 212859 4675
rect 213469 4641 213503 4675
rect 213862 4641 213896 4675
rect 215401 4641 215435 4675
rect 217977 4641 218011 4675
rect 218161 4641 218195 4675
rect 219449 4641 219483 4675
rect 221105 4641 221139 4675
rect 221749 4641 221783 4675
rect 247601 4641 247635 4675
rect 249073 4641 249107 4675
rect 250729 4641 250763 4675
rect 251465 4641 251499 4675
rect 252753 4641 252787 4675
rect 256617 4641 256651 4675
rect 258825 4641 258859 4675
rect 270049 4641 270083 4675
rect 36001 4573 36035 4607
rect 41797 4573 41831 4607
rect 42257 4573 42291 4607
rect 47041 4573 47075 4607
rect 47501 4573 47535 4607
rect 91753 4573 91787 4607
rect 92765 4573 92799 4607
rect 94329 4573 94363 4607
rect 96721 4573 96755 4607
rect 99757 4573 99791 4607
rect 100125 4573 100159 4607
rect 100769 4573 100803 4607
rect 101045 4573 101079 4607
rect 104817 4573 104851 4607
rect 105461 4573 105495 4607
rect 105921 4573 105955 4607
rect 107025 4573 107059 4607
rect 108037 4573 108071 4607
rect 108405 4573 108439 4607
rect 109141 4573 109175 4607
rect 111625 4573 111659 4607
rect 112361 4573 112395 4607
rect 113005 4573 113039 4607
rect 113649 4573 113683 4607
rect 114109 4573 114143 4607
rect 114293 4573 114327 4607
rect 114937 4573 114971 4607
rect 117329 4573 117363 4607
rect 118893 4573 118927 4607
rect 119445 4573 119479 4607
rect 120273 4573 120307 4607
rect 120641 4573 120675 4607
rect 121285 4573 121319 4607
rect 122481 4573 122515 4607
rect 138397 4573 138431 4607
rect 139133 4573 139167 4607
rect 141571 4573 141605 4607
rect 143089 4573 143123 4607
rect 145527 4573 145561 4607
rect 147137 4573 147171 4607
rect 148425 4573 148459 4607
rect 150035 4573 150069 4607
rect 151277 4573 151311 4607
rect 151553 4573 151587 4607
rect 152289 4573 152323 4607
rect 155693 4573 155727 4607
rect 158729 4573 158763 4607
rect 159465 4573 159499 4607
rect 159603 4573 159637 4607
rect 159741 4573 159775 4607
rect 166273 4573 166307 4607
rect 167193 4573 167227 4607
rect 167469 4573 167503 4607
rect 168941 4573 168975 4607
rect 205649 4573 205683 4607
rect 205741 4573 205775 4607
rect 205833 4573 205867 4607
rect 208869 4573 208903 4607
rect 208961 4573 208995 4607
rect 209053 4573 209087 4607
rect 211537 4573 211571 4607
rect 211629 4573 211663 4607
rect 211813 4573 211847 4607
rect 213009 4573 213043 4607
rect 213745 4573 213779 4607
rect 214021 4573 214055 4607
rect 214665 4573 214699 4607
rect 215217 4573 215251 4607
rect 220553 4573 220587 4607
rect 221289 4573 221323 4607
rect 222025 4573 222059 4607
rect 222142 4573 222176 4607
rect 222301 4573 222335 4607
rect 223681 4573 223715 4607
rect 223865 4573 223899 4607
rect 224693 4573 224727 4607
rect 225521 4573 225555 4607
rect 227361 4573 227395 4607
rect 244933 4573 244967 4607
rect 245577 4573 245611 4607
rect 246865 4573 246899 4607
rect 246957 4573 246991 4607
rect 247877 4573 247911 4607
rect 248889 4573 248923 4607
rect 251557 4573 251591 4607
rect 252845 4573 252879 4607
rect 253397 4573 253431 4607
rect 255881 4573 255915 4607
rect 256433 4573 256467 4607
rect 259009 4573 259043 4607
rect 259837 4573 259871 4607
rect 261769 4573 261803 4607
rect 264253 4573 264287 4607
rect 264897 4573 264931 4607
rect 265541 4573 265575 4607
rect 266185 4573 266219 4607
rect 266921 4573 266955 4607
rect 268577 4573 268611 4607
rect 269681 4573 269715 4607
rect 269865 4573 269899 4607
rect 270509 4573 270543 4607
rect 36093 4505 36127 4539
rect 36461 4505 36495 4539
rect 41889 4505 41923 4539
rect 47133 4505 47167 4539
rect 96169 4505 96203 4539
rect 104173 4505 104207 4539
rect 110981 4505 111015 4539
rect 115121 4505 115155 4539
rect 116777 4505 116811 4539
rect 147321 4505 147355 4539
rect 206017 4505 206051 4539
rect 206661 4505 206695 4539
rect 208317 4505 208351 4539
rect 210157 4505 210191 4539
rect 217057 4505 217091 4539
rect 223405 4505 223439 4539
rect 225705 4505 225739 4539
rect 246681 4505 246715 4539
rect 251281 4505 251315 4539
rect 252569 4505 252603 4539
rect 252937 4505 252971 4539
rect 253581 4505 253615 4539
rect 255237 4505 255271 4539
rect 258273 4505 258307 4539
rect 258733 4505 258767 4539
rect 267289 4505 267323 4539
rect 268945 4505 268979 4539
rect 35173 4437 35207 4471
rect 35725 4437 35759 4471
rect 36829 4437 36863 4471
rect 41521 4437 41555 4471
rect 42625 4437 42659 4471
rect 46765 4437 46799 4471
rect 47869 4437 47903 4471
rect 93409 4437 93443 4471
rect 96905 4437 96939 4471
rect 100309 4437 100343 4471
rect 104633 4437 104667 4471
rect 105277 4437 105311 4471
rect 107577 4437 107611 4471
rect 111441 4437 111475 4471
rect 123033 4437 123067 4471
rect 140053 4437 140087 4471
rect 142353 4437 142387 4471
rect 146309 4437 146343 4471
rect 148241 4437 148275 4471
rect 150817 4437 150851 4471
rect 151829 4437 151863 4471
rect 152841 4437 152875 4471
rect 160385 4437 160419 4471
rect 165997 4437 166031 4471
rect 209237 4437 209271 4471
rect 210249 4437 210283 4471
rect 220369 4437 220403 4471
rect 224049 4437 224083 4471
rect 245393 4437 245427 4471
rect 247141 4437 247175 4471
rect 251741 4437 251775 4471
rect 255697 4437 255731 4471
rect 259653 4437 259687 4471
rect 261585 4437 261619 4471
rect 264069 4437 264103 4471
rect 41797 4233 41831 4267
rect 49617 4233 49651 4267
rect 49801 4233 49835 4267
rect 50537 4233 50571 4267
rect 110797 4233 110831 4267
rect 148517 4233 148551 4267
rect 155049 4233 155083 4267
rect 244381 4233 244415 4267
rect 267289 4233 267323 4267
rect 268577 4233 268611 4267
rect 270785 4233 270819 4267
rect 37657 4165 37691 4199
rect 38761 4165 38795 4199
rect 39313 4165 39347 4199
rect 41705 4165 41739 4199
rect 44465 4165 44499 4199
rect 44833 4165 44867 4199
rect 45569 4165 45603 4199
rect 48513 4165 48547 4199
rect 49249 4165 49283 4199
rect 50813 4165 50847 4199
rect 51273 4165 51307 4199
rect 51641 4165 51675 4199
rect 98745 4165 98779 4199
rect 205833 4165 205867 4199
rect 215769 4165 215803 4199
rect 216689 4165 216723 4199
rect 217057 4165 217091 4199
rect 252845 4165 252879 4199
rect 259837 4165 259871 4199
rect 36829 4097 36863 4131
rect 37933 4097 37967 4131
rect 38025 4097 38059 4131
rect 38393 4097 38427 4131
rect 39681 4097 39715 4131
rect 42625 4097 42659 4131
rect 44741 4097 44775 4131
rect 45201 4097 45235 4131
rect 48789 4097 48823 4131
rect 48881 4097 48915 4131
rect 50905 4097 50939 4131
rect 66913 4097 66947 4131
rect 92949 4097 92983 4131
rect 93593 4097 93627 4131
rect 94605 4097 94639 4131
rect 102057 4097 102091 4131
rect 104725 4097 104759 4131
rect 108497 4097 108531 4131
rect 108773 4097 108807 4131
rect 109785 4097 109819 4131
rect 110245 4097 110279 4131
rect 114201 4097 114235 4131
rect 117053 4097 117087 4131
rect 118249 4097 118283 4131
rect 120457 4097 120491 4131
rect 120825 4097 120859 4131
rect 138397 4097 138431 4131
rect 139409 4097 139443 4131
rect 142813 4097 142847 4131
rect 143825 4097 143859 4131
rect 145021 4097 145055 4131
rect 146861 4097 146895 4131
rect 147505 4097 147539 4131
rect 147965 4097 147999 4131
rect 148977 4097 149011 4131
rect 150265 4097 150299 4131
rect 150817 4097 150851 4131
rect 153209 4097 153243 4131
rect 167653 4097 167687 4131
rect 168113 4097 168147 4131
rect 190469 4097 190503 4131
rect 206017 4097 206051 4131
rect 206569 4097 206603 4131
rect 206661 4097 206695 4131
rect 206753 4097 206787 4131
rect 213193 4097 213227 4131
rect 217977 4097 218011 4131
rect 220277 4097 220311 4131
rect 222945 4097 222979 4131
rect 223865 4097 223899 4131
rect 224003 4097 224037 4131
rect 224141 4097 224175 4131
rect 224785 4097 224819 4131
rect 236561 4097 236595 4131
rect 244565 4097 244599 4131
rect 245030 4097 245064 4131
rect 247325 4097 247359 4131
rect 247601 4097 247635 4131
rect 251005 4097 251039 4131
rect 253121 4097 253155 4131
rect 254133 4097 254167 4131
rect 254409 4097 254443 4131
rect 256893 4097 256927 4131
rect 257353 4097 257387 4131
rect 257537 4097 257571 4131
rect 257629 4097 257663 4131
rect 258457 4097 258491 4131
rect 259009 4097 259043 4131
rect 265173 4097 265207 4131
rect 265817 4097 265851 4131
rect 266461 4097 266495 4131
rect 267013 4097 267047 4131
rect 267105 4097 267139 4131
rect 267933 4097 267967 4131
rect 269313 4097 269347 4131
rect 270049 4097 270083 4131
rect 270969 4097 271003 4131
rect 42809 4029 42843 4063
rect 66453 4029 66487 4063
rect 94789 4029 94823 4063
rect 96169 4029 96203 4063
rect 96905 4029 96939 4063
rect 97089 4029 97123 4063
rect 99297 4029 99331 4063
rect 99481 4029 99515 4063
rect 101137 4029 101171 4063
rect 102241 4029 102275 4063
rect 103897 4029 103931 4063
rect 105001 4029 105035 4063
rect 105737 4029 105771 4063
rect 105921 4029 105955 4063
rect 107577 4029 107611 4063
rect 110521 4029 110555 4063
rect 111625 4029 111659 4063
rect 111809 4029 111843 4063
rect 112085 4029 112119 4063
rect 114753 4029 114787 4063
rect 114937 4029 114971 4063
rect 116593 4029 116627 4063
rect 117237 4029 117271 4063
rect 117697 4029 117731 4063
rect 117973 4029 118007 4063
rect 118090 4029 118124 4063
rect 121469 4029 121503 4063
rect 121653 4029 121687 4063
rect 123309 4029 123343 4063
rect 138673 4029 138707 4063
rect 139685 4029 139719 4063
rect 140513 4029 140547 4063
rect 140697 4029 140731 4063
rect 140973 4029 141007 4063
rect 143089 4029 143123 4063
rect 144101 4029 144135 4063
rect 145665 4029 145699 4063
rect 145849 4029 145883 4063
rect 146309 4029 146343 4063
rect 146585 4029 146619 4063
rect 146723 4029 146757 4063
rect 148241 4029 148275 4063
rect 149253 4029 149287 4063
rect 151001 4029 151035 4063
rect 152013 4029 152047 4063
rect 153393 4029 153427 4063
rect 153853 4029 153887 4063
rect 154129 4029 154163 4063
rect 154246 4029 154280 4063
rect 154405 4029 154439 4063
rect 155969 4029 156003 4063
rect 156153 4029 156187 4063
rect 157073 4029 157107 4063
rect 158269 4029 158303 4063
rect 158453 4029 158487 4063
rect 160017 4029 160051 4063
rect 168021 4029 168055 4063
rect 207489 4029 207523 4063
rect 207673 4029 207707 4063
rect 209329 4029 209363 4063
rect 209789 4029 209823 4063
rect 209973 4029 210007 4063
rect 210249 4029 210283 4063
rect 213377 4029 213411 4063
rect 213929 4029 213963 4063
rect 217793 4029 217827 4063
rect 218437 4029 218471 4063
rect 218713 4029 218747 4063
rect 218830 4029 218864 4063
rect 218989 4029 219023 4063
rect 220093 4029 220127 4063
rect 221013 4029 221047 4063
rect 221151 4029 221185 4063
rect 221289 4029 221323 4063
rect 223129 4029 223163 4063
rect 223589 4029 223623 4063
rect 225245 4029 225279 4063
rect 225429 4029 225463 4063
rect 226717 4029 226751 4063
rect 236837 4029 236871 4063
rect 245209 4029 245243 4063
rect 246865 4029 246899 4063
rect 248705 4029 248739 4063
rect 248889 4029 248923 4063
rect 250545 4029 250579 4063
rect 251281 4029 251315 4063
rect 253029 4029 253063 4063
rect 254317 4029 254351 4063
rect 255053 4029 255087 4063
rect 255237 4029 255271 4063
rect 259653 4029 259687 4063
rect 260757 4029 260791 4063
rect 267749 4029 267783 4063
rect 38945 3961 38979 3995
rect 51825 3961 51859 3995
rect 93409 3961 93443 3995
rect 105277 3961 105311 3995
rect 109601 3961 109635 3995
rect 114017 3961 114051 3995
rect 121009 3961 121043 3995
rect 144377 3961 144411 3995
rect 150081 3961 150115 3995
rect 206937 3961 206971 3995
rect 220737 3961 220771 3995
rect 257813 3961 257847 3995
rect 266277 3961 266311 3995
rect 269497 3961 269531 3995
rect 270233 3961 270267 3995
rect 45753 3893 45787 3927
rect 47961 3893 47995 3927
rect 66729 3893 66763 3927
rect 92765 3893 92799 3927
rect 104817 3893 104851 3927
rect 108865 3893 108899 3927
rect 109049 3893 109083 3927
rect 110613 3893 110647 3927
rect 118893 3893 118927 3927
rect 120825 3893 120859 3927
rect 138765 3893 138799 3927
rect 138949 3893 138983 3927
rect 139593 3893 139627 3927
rect 139961 3893 139995 3927
rect 142905 3893 142939 3927
rect 143365 3893 143399 3927
rect 143917 3893 143951 3927
rect 144837 3893 144871 3927
rect 148057 3893 148091 3927
rect 149069 3893 149103 3927
rect 149529 3893 149563 3927
rect 167745 3893 167779 3927
rect 168297 3893 168331 3927
rect 190285 3893 190319 3927
rect 216045 3893 216079 3927
rect 219633 3893 219667 3927
rect 221933 3893 221967 3927
rect 225153 3893 225187 3927
rect 252845 3893 252879 3927
rect 253305 3893 253339 3927
rect 254133 3893 254167 3927
rect 254593 3893 254627 3927
rect 257353 3893 257387 3927
rect 258273 3893 258307 3927
rect 258825 3893 258859 3927
rect 259285 3893 259319 3927
rect 264989 3893 265023 3927
rect 268117 3893 268151 3927
rect 92581 3689 92615 3723
rect 95801 3689 95835 3723
rect 96997 3689 97031 3723
rect 101873 3689 101907 3723
rect 102241 3689 102275 3723
rect 105369 3689 105403 3723
rect 106197 3689 106231 3723
rect 106473 3689 106507 3723
rect 111625 3689 111659 3723
rect 119629 3689 119663 3723
rect 122481 3689 122515 3723
rect 138949 3689 138983 3723
rect 141985 3689 142019 3723
rect 148241 3689 148275 3723
rect 149253 3689 149287 3723
rect 155233 3689 155267 3723
rect 208869 3689 208903 3723
rect 214389 3689 214423 3723
rect 244473 3689 244507 3723
rect 245393 3689 245427 3723
rect 246497 3689 246531 3723
rect 246681 3689 246715 3723
rect 252569 3689 252603 3723
rect 258733 3689 258767 3723
rect 260573 3689 260607 3723
rect 267933 3689 267967 3723
rect 269221 3689 269255 3723
rect 270049 3689 270083 3723
rect 68845 3621 68879 3655
rect 92029 3621 92063 3655
rect 94605 3621 94639 3655
rect 102793 3621 102827 3655
rect 104173 3621 104207 3655
rect 118433 3621 118467 3655
rect 152565 3621 152599 3655
rect 154037 3621 154071 3655
rect 156337 3621 156371 3655
rect 212089 3621 212123 3655
rect 220369 3621 220403 3655
rect 227361 3621 227395 3655
rect 253029 3621 253063 3655
rect 268577 3621 268611 3655
rect 94881 3553 94915 3587
rect 95019 3553 95053 3587
rect 95157 3553 95191 3587
rect 99113 3553 99147 3587
rect 99297 3553 99331 3587
rect 101965 3553 101999 3587
rect 103713 3553 103747 3587
rect 104449 3553 104483 3587
rect 104566 3553 104600 3587
rect 104725 3553 104759 3587
rect 107209 3553 107243 3587
rect 108865 3553 108899 3587
rect 109785 3553 109819 3587
rect 110429 3553 110463 3587
rect 110705 3553 110739 3587
rect 110981 3553 111015 3587
rect 112177 3553 112211 3587
rect 113741 3553 113775 3587
rect 115121 3553 115155 3587
rect 118709 3553 118743 3587
rect 120089 3553 120123 3587
rect 120273 3553 120307 3587
rect 150265 3553 150299 3587
rect 153393 3553 153427 3587
rect 153577 3553 153611 3587
rect 154313 3553 154347 3587
rect 155877 3553 155911 3587
rect 156613 3553 156647 3587
rect 156751 3553 156785 3587
rect 207029 3553 207063 3587
rect 207213 3553 207247 3587
rect 207673 3553 207707 3587
rect 208087 3553 208121 3587
rect 217425 3553 217459 3587
rect 221105 3553 221139 3587
rect 222577 3553 222611 3587
rect 224141 3553 224175 3587
rect 226165 3553 226199 3587
rect 226441 3553 226475 3587
rect 226579 3553 226613 3587
rect 245301 3553 245335 3587
rect 246405 3553 246439 3587
rect 247325 3553 247359 3587
rect 248705 3553 248739 3587
rect 251557 3553 251591 3587
rect 252661 3553 252695 3587
rect 254041 3553 254075 3587
rect 255881 3553 255915 3587
rect 258273 3553 258307 3587
rect 258825 3553 258859 3587
rect 266001 3553 266035 3587
rect 23397 3485 23431 3519
rect 36645 3485 36679 3519
rect 37105 3485 37139 3519
rect 41061 3485 41095 3519
rect 41153 3485 41187 3519
rect 43545 3485 43579 3519
rect 44005 3485 44039 3519
rect 48973 3485 49007 3519
rect 50813 3485 50847 3519
rect 50905 3485 50939 3519
rect 68753 3485 68787 3519
rect 91937 3485 91971 3519
rect 92765 3485 92799 3519
rect 93225 3485 93259 3519
rect 93961 3485 93995 3519
rect 94145 3485 94179 3519
rect 96997 3485 97031 3519
rect 97181 3485 97215 3519
rect 97825 3485 97859 3519
rect 98101 3485 98135 3519
rect 101873 3485 101907 3519
rect 102609 3485 102643 3519
rect 103529 3485 103563 3519
rect 105921 3485 105955 3519
rect 106197 3485 106231 3519
rect 107025 3485 107059 3519
rect 109969 3485 110003 3519
rect 110843 3485 110877 3519
rect 114937 3485 114971 3519
rect 117789 3485 117823 3519
rect 117973 3485 118007 3519
rect 118847 3485 118881 3519
rect 118985 3485 119019 3519
rect 121929 3485 121963 3519
rect 122665 3485 122699 3519
rect 138489 3485 138523 3519
rect 139133 3485 139167 3519
rect 139593 3485 139627 3519
rect 141433 3485 141467 3519
rect 141893 3485 141927 3519
rect 142261 3485 142295 3519
rect 143089 3485 143123 3519
rect 145389 3485 145423 3519
rect 148425 3485 148459 3519
rect 149161 3485 149195 3519
rect 149437 3485 149471 3519
rect 152749 3485 152783 3519
rect 154451 3485 154485 3519
rect 154589 3485 154623 3519
rect 155693 3485 155727 3519
rect 156889 3485 156923 3519
rect 158729 3485 158763 3519
rect 159373 3485 159407 3519
rect 167653 3485 167687 3519
rect 207949 3485 207983 3519
rect 208225 3485 208259 3519
rect 210249 3485 210283 3519
rect 210341 3485 210375 3519
rect 210525 3485 210559 3519
rect 211445 3485 211479 3519
rect 211537 3485 211571 3519
rect 211721 3485 211755 3519
rect 212641 3485 212675 3519
rect 212733 3485 212767 3519
rect 213009 3485 213043 3519
rect 213929 3485 213963 3519
rect 214573 3485 214607 3519
rect 215585 3485 215619 3519
rect 215769 3485 215803 3519
rect 216505 3485 216539 3519
rect 216597 3485 216631 3519
rect 216689 3485 216723 3519
rect 220553 3485 220587 3519
rect 223497 3485 223531 3519
rect 223589 3485 223623 3519
rect 223773 3485 223807 3519
rect 224601 3485 224635 3519
rect 225521 3485 225555 3519
rect 225705 3485 225739 3519
rect 226717 3485 226751 3519
rect 244381 3485 244415 3519
rect 244473 3485 244507 3519
rect 245393 3485 245427 3519
rect 246497 3485 246531 3519
rect 247049 3485 247083 3519
rect 248521 3485 248555 3519
rect 251281 3485 251315 3519
rect 252845 3485 252879 3519
rect 256433 3485 256467 3519
rect 259009 3485 259043 3519
rect 260389 3485 260423 3519
rect 267473 3485 267507 3519
rect 268117 3485 268151 3519
rect 268761 3485 268795 3519
rect 269405 3485 269439 3519
rect 269865 3485 269899 3519
rect 270969 3485 271003 3519
rect 36737 3417 36771 3451
rect 40233 3417 40267 3451
rect 41521 3417 41555 3451
rect 41889 3417 41923 3451
rect 43637 3417 43671 3451
rect 48237 3417 48271 3451
rect 48513 3417 48547 3451
rect 48605 3417 48639 3451
rect 51273 3417 51307 3451
rect 100953 3417 100987 3451
rect 103161 3417 103195 3451
rect 112361 3417 112395 3451
rect 116777 3417 116811 3451
rect 139777 3417 139811 3451
rect 143273 3417 143307 3451
rect 144929 3417 144963 3451
rect 145573 3417 145607 3451
rect 147229 3417 147263 3451
rect 150449 3417 150483 3451
rect 152105 3417 152139 3451
rect 210893 3417 210927 3451
rect 213285 3417 213319 3451
rect 216873 3417 216907 3451
rect 217609 3417 217643 3451
rect 219265 3417 219299 3451
rect 221289 3417 221323 3451
rect 244197 3417 244231 3451
rect 245117 3417 245151 3451
rect 246221 3417 246255 3451
rect 248153 3417 248187 3451
rect 250361 3417 250395 3451
rect 252569 3417 252603 3451
rect 254225 3417 254259 3451
rect 256617 3417 256651 3451
rect 258733 3417 258767 3451
rect 259745 3417 259779 3451
rect 23581 3349 23615 3383
rect 36369 3349 36403 3383
rect 37473 3349 37507 3383
rect 37657 3349 37691 3383
rect 40785 3349 40819 3383
rect 42073 3349 42107 3383
rect 43269 3349 43303 3383
rect 44373 3349 44407 3383
rect 44557 3349 44591 3383
rect 49341 3349 49375 3383
rect 49525 3349 49559 3383
rect 50537 3349 50571 3383
rect 51641 3349 51675 3383
rect 51825 3349 51859 3383
rect 93409 3349 93443 3383
rect 97365 3349 97399 3383
rect 138305 3349 138339 3383
rect 142445 3349 142479 3383
rect 149713 3349 149747 3383
rect 157533 3349 157567 3383
rect 158545 3349 158579 3383
rect 159189 3349 159223 3383
rect 167745 3349 167779 3383
rect 213745 3349 213779 3383
rect 224693 3349 224727 3383
rect 227729 3349 227763 3383
rect 244657 3349 244691 3383
rect 245577 3349 245611 3383
rect 259193 3349 259227 3383
rect 259837 3349 259871 3383
rect 267289 3349 267323 3383
rect 270785 3349 270819 3383
rect 38761 3145 38795 3179
rect 38945 3145 38979 3179
rect 44097 3145 44131 3179
rect 44281 3145 44315 3179
rect 96445 3145 96479 3179
rect 106289 3145 106323 3179
rect 148057 3145 148091 3179
rect 153761 3145 153795 3179
rect 154405 3145 154439 3179
rect 210801 3145 210835 3179
rect 220921 3145 220955 3179
rect 225705 3145 225739 3179
rect 244473 3145 244507 3179
rect 257675 3145 257709 3179
rect 267289 3145 267323 3179
rect 268577 3145 268611 3179
rect 270785 3145 270819 3179
rect 37657 3077 37691 3111
rect 37933 3077 37967 3111
rect 38025 3077 38059 3111
rect 42993 3077 43027 3111
rect 43269 3077 43303 3111
rect 43361 3077 43395 3111
rect 43729 3077 43763 3111
rect 47961 3077 47995 3111
rect 49065 3077 49099 3111
rect 95249 3077 95283 3111
rect 97089 3077 97123 3111
rect 99757 3077 99791 3111
rect 102057 3077 102091 3111
rect 103713 3077 103747 3111
rect 107393 3077 107427 3111
rect 140697 3077 140731 3111
rect 143089 3077 143123 3111
rect 145849 3077 145883 3111
rect 212825 3077 212859 3111
rect 215125 3077 215159 3111
rect 225245 3077 225279 3111
rect 244013 3077 244047 3111
rect 245117 3077 245151 3111
rect 248889 3077 248923 3111
rect 252845 3077 252879 3111
rect 22661 3009 22695 3043
rect 22845 3009 22879 3043
rect 23673 3009 23707 3043
rect 24501 3009 24535 3043
rect 24593 3009 24627 3043
rect 25605 3009 25639 3043
rect 26341 3009 26375 3043
rect 38393 3009 38427 3043
rect 48230 3009 48264 3043
rect 48329 3009 48363 3043
rect 48697 3009 48731 3043
rect 49617 3009 49651 3043
rect 54309 3009 54343 3043
rect 89361 3009 89395 3043
rect 90649 3009 90683 3043
rect 91845 3009 91879 3043
rect 92581 3009 92615 3043
rect 93317 3009 93351 3043
rect 94145 3009 94179 3043
rect 94973 3009 95007 3043
rect 95065 3009 95099 3043
rect 96261 3009 96295 3043
rect 96905 3009 96939 3043
rect 99573 3009 99607 3043
rect 104449 3009 104483 3043
rect 104633 3009 104667 3043
rect 105369 3009 105403 3043
rect 105645 3009 105679 3043
rect 109785 3009 109819 3043
rect 110245 3009 110279 3043
rect 115029 3009 115063 3043
rect 119353 3009 119387 3043
rect 119997 3009 120031 3043
rect 138397 3009 138431 3043
rect 139041 3009 139075 3043
rect 139685 3009 139719 3043
rect 148425 3009 148459 3043
rect 149345 3009 149379 3043
rect 149621 3009 149655 3043
rect 153301 3009 153335 3043
rect 153945 3009 153979 3043
rect 154589 3009 154623 3043
rect 155233 3009 155267 3043
rect 156153 3009 156187 3043
rect 158453 3009 158487 3043
rect 159189 3009 159223 3043
rect 190929 3009 190963 3043
rect 207673 3009 207707 3043
rect 207765 3009 207799 3043
rect 207949 3009 207983 3043
rect 208961 3009 208995 3043
rect 209998 3009 210032 3043
rect 210157 3009 210191 3043
rect 211353 3009 211387 3043
rect 211445 3009 211479 3043
rect 211629 3009 211663 3043
rect 220553 3009 220587 3043
rect 220645 3009 220679 3043
rect 220749 3015 220783 3049
rect 221473 3009 221507 3043
rect 221657 3009 221691 3043
rect 221841 3009 221875 3043
rect 223405 3009 223439 3043
rect 224325 3009 224359 3043
rect 224601 3009 224635 3043
rect 225889 3009 225923 3043
rect 226533 3009 226567 3043
rect 244289 3009 244323 3043
rect 246773 3009 246807 3043
rect 248705 3009 248739 3043
rect 251005 3009 251039 3043
rect 254133 3009 254167 3043
rect 257445 3009 257479 3043
rect 259101 3009 259135 3043
rect 259745 3009 259779 3043
rect 260481 3009 260515 3043
rect 261125 3009 261159 3043
rect 261861 3009 261895 3043
rect 267473 3009 267507 3043
rect 268117 3009 268151 3043
rect 268761 3009 268795 3043
rect 269865 3009 269899 3043
rect 270969 3009 271003 3043
rect 32321 2941 32355 2975
rect 66361 2941 66395 2975
rect 96077 2941 96111 2975
rect 98745 2941 98779 2975
rect 101413 2941 101447 2975
rect 101873 2941 101907 2975
rect 105486 2941 105520 2975
rect 107209 2941 107243 2975
rect 108957 2941 108991 2975
rect 110521 2941 110555 2975
rect 111809 2941 111843 2975
rect 111993 2941 112027 2975
rect 113465 2941 113499 2975
rect 115213 2941 115247 2975
rect 116869 2941 116903 2975
rect 117513 2941 117547 2975
rect 117697 2941 117731 2975
rect 120181 2941 120215 2975
rect 120733 2941 120767 2975
rect 120917 2941 120951 2975
rect 121837 2941 121871 2975
rect 135361 2941 135395 2975
rect 140513 2941 140547 2975
rect 142077 2941 142111 2975
rect 142905 2941 142939 2975
rect 143549 2941 143583 2975
rect 145665 2941 145699 2975
rect 146493 2941 146527 2975
rect 148609 2941 148643 2975
rect 149483 2941 149517 2975
rect 150265 2941 150299 2975
rect 150817 2941 150851 2975
rect 151001 2941 151035 2975
rect 152657 2941 152691 2975
rect 156337 2941 156371 2975
rect 156613 2941 156647 2975
rect 167929 2941 167963 2975
rect 203165 2941 203199 2975
rect 209145 2941 209179 2975
rect 209881 2941 209915 2975
rect 212641 2941 212675 2975
rect 214297 2941 214331 2975
rect 214941 2941 214975 2975
rect 215401 2941 215435 2975
rect 218161 2941 218195 2975
rect 218345 2941 218379 2975
rect 219633 2941 219667 2975
rect 223589 2941 223623 2975
rect 224049 2941 224083 2975
rect 224463 2941 224497 2975
rect 235733 2941 235767 2975
rect 244197 2941 244231 2975
rect 244933 2941 244967 2975
rect 247233 2941 247267 2975
rect 247509 2941 247543 2975
rect 250545 2941 250579 2975
rect 251189 2941 251223 2975
rect 253857 2941 253891 2975
rect 255145 2941 255179 2975
rect 255329 2941 255363 2975
rect 256985 2941 257019 2975
rect 260297 2941 260331 2975
rect 260665 2941 260699 2975
rect 266645 2941 266679 2975
rect 44649 2873 44683 2907
rect 49249 2873 49283 2907
rect 93501 2873 93535 2907
rect 105093 2873 105127 2907
rect 110797 2873 110831 2907
rect 139501 2873 139535 2907
rect 149069 2873 149103 2907
rect 153117 2873 153151 2907
rect 208317 2873 208351 2907
rect 209605 2873 209639 2907
rect 211905 2873 211939 2907
rect 262045 2873 262079 2907
rect 23029 2805 23063 2839
rect 23857 2805 23891 2839
rect 24777 2805 24811 2839
rect 25789 2805 25823 2839
rect 26525 2805 26559 2839
rect 54493 2805 54527 2839
rect 89545 2805 89579 2839
rect 90833 2805 90867 2839
rect 92029 2805 92063 2839
rect 92765 2805 92799 2839
rect 94329 2805 94363 2839
rect 109601 2805 109635 2839
rect 110521 2805 110555 2839
rect 138213 2805 138247 2839
rect 138857 2805 138891 2839
rect 155049 2805 155083 2839
rect 158637 2805 158671 2839
rect 159373 2805 159407 2839
rect 191113 2805 191147 2839
rect 208685 2805 208719 2839
rect 221565 2805 221599 2839
rect 226349 2805 226383 2839
rect 244289 2805 244323 2839
rect 259193 2805 259227 2839
rect 261309 2805 261343 2839
rect 266185 2805 266219 2839
rect 267933 2805 267967 2839
rect 270049 2805 270083 2839
rect 1777 2601 1811 2635
rect 22017 2601 22051 2635
rect 23765 2601 23799 2635
rect 24593 2601 24627 2635
rect 27629 2601 27663 2635
rect 43545 2601 43579 2635
rect 55689 2601 55723 2635
rect 76711 2601 76745 2635
rect 124229 2601 124263 2635
rect 133981 2601 134015 2635
rect 138673 2601 138707 2635
rect 141157 2601 141191 2635
rect 141985 2601 142019 2635
rect 153393 2601 153427 2635
rect 154681 2601 154715 2635
rect 155785 2601 155819 2635
rect 190561 2601 190595 2635
rect 192033 2601 192067 2635
rect 198749 2601 198783 2635
rect 219357 2601 219391 2635
rect 226993 2601 227027 2635
rect 268301 2601 268335 2635
rect 270141 2601 270175 2635
rect 24961 2533 24995 2567
rect 94973 2533 95007 2567
rect 200405 2533 200439 2567
rect 201969 2533 202003 2567
rect 218161 2533 218195 2567
rect 230949 2533 230983 2567
rect 262597 2533 262631 2567
rect 4813 2465 4847 2499
rect 22569 2465 22603 2499
rect 23397 2465 23431 2499
rect 25329 2465 25363 2499
rect 26433 2465 26467 2499
rect 66821 2465 66855 2499
rect 81909 2465 81943 2499
rect 84117 2465 84151 2499
rect 94329 2465 94363 2499
rect 94513 2465 94547 2499
rect 95249 2465 95283 2499
rect 95387 2465 95421 2499
rect 97365 2465 97399 2499
rect 99665 2465 99699 2499
rect 101965 2465 101999 2499
rect 102149 2465 102183 2499
rect 104817 2465 104851 2499
rect 106197 2465 106231 2499
rect 107209 2465 107243 2499
rect 107669 2465 107703 2499
rect 109509 2465 109543 2499
rect 111165 2465 111199 2499
rect 112637 2465 112671 2499
rect 115029 2465 115063 2499
rect 119721 2465 119755 2499
rect 120273 2465 120307 2499
rect 124781 2465 124815 2499
rect 129749 2465 129783 2499
rect 134625 2465 134659 2499
rect 139317 2465 139351 2499
rect 139961 2465 139995 2499
rect 145573 2465 145607 2499
rect 146309 2465 146343 2499
rect 148609 2465 148643 2499
rect 148793 2465 148827 2499
rect 150265 2465 150299 2499
rect 151093 2465 151127 2499
rect 151369 2465 151403 2499
rect 182097 2465 182131 2499
rect 185041 2465 185075 2499
rect 187249 2465 187283 2499
rect 210065 2465 210099 2499
rect 212549 2465 212583 2499
rect 215401 2465 215435 2499
rect 216781 2465 216815 2499
rect 217517 2465 217551 2499
rect 223129 2465 223163 2499
rect 246129 2465 246163 2499
rect 248981 2465 249015 2499
rect 250637 2465 250671 2499
rect 251465 2465 251499 2499
rect 253857 2465 253891 2499
rect 256617 2465 256651 2499
rect 258273 2465 258307 2499
rect 261585 2465 261619 2499
rect 263977 2465 264011 2499
rect 264897 2465 264931 2499
rect 269773 2465 269807 2499
rect 4537 2397 4571 2431
rect 6745 2397 6779 2431
rect 7021 2397 7055 2431
rect 14841 2397 14875 2431
rect 15117 2397 15151 2431
rect 21833 2397 21867 2431
rect 22753 2397 22787 2431
rect 23581 2397 23615 2431
rect 24409 2397 24443 2431
rect 25513 2397 25547 2431
rect 26157 2397 26191 2431
rect 27445 2397 27479 2431
rect 29745 2397 29779 2431
rect 31953 2397 31987 2431
rect 32045 2397 32079 2431
rect 32781 2397 32815 2431
rect 38393 2397 38427 2431
rect 38853 2397 38887 2431
rect 40509 2397 40543 2431
rect 40969 2397 41003 2431
rect 42533 2397 42567 2431
rect 42993 2397 43027 2431
rect 53757 2397 53791 2431
rect 54033 2397 54067 2431
rect 54217 2397 54251 2431
rect 55505 2397 55539 2431
rect 57805 2397 57839 2431
rect 59277 2397 59311 2431
rect 61485 2397 61519 2431
rect 62221 2397 62255 2431
rect 62957 2397 62991 2431
rect 65809 2397 65843 2431
rect 66545 2397 66579 2431
rect 76481 2397 76515 2431
rect 78689 2397 78723 2431
rect 78965 2397 78999 2431
rect 81633 2397 81667 2431
rect 83841 2397 83875 2431
rect 88901 2397 88935 2431
rect 89085 2397 89119 2431
rect 90005 2397 90039 2431
rect 90741 2397 90775 2431
rect 92213 2397 92247 2431
rect 92857 2397 92891 2431
rect 93593 2397 93627 2431
rect 95525 2397 95559 2431
rect 96169 2397 96203 2431
rect 97181 2397 97215 2431
rect 99481 2397 99515 2431
rect 101321 2397 101355 2431
rect 104633 2397 104667 2431
rect 107025 2397 107059 2431
rect 109325 2397 109359 2431
rect 112177 2397 112211 2431
rect 114845 2397 114879 2431
rect 117513 2397 117547 2431
rect 118157 2397 118191 2431
rect 118801 2397 118835 2431
rect 119537 2397 119571 2431
rect 122573 2397 122607 2431
rect 124045 2397 124079 2431
rect 124965 2397 124999 2431
rect 126069 2397 126103 2431
rect 126805 2397 126839 2431
rect 128277 2397 128311 2431
rect 129013 2397 129047 2431
rect 129933 2397 129967 2431
rect 130117 2397 130151 2431
rect 130577 2397 130611 2431
rect 131497 2397 131531 2431
rect 133061 2397 133095 2431
rect 133797 2397 133831 2431
rect 134809 2397 134843 2431
rect 138857 2397 138891 2431
rect 139501 2397 139535 2431
rect 140237 2397 140271 2431
rect 140354 2397 140388 2431
rect 140513 2397 140547 2431
rect 141617 2397 141651 2431
rect 141985 2397 142019 2431
rect 143089 2397 143123 2431
rect 145389 2397 145423 2431
rect 150909 2397 150943 2431
rect 153577 2397 153611 2431
rect 154221 2397 154255 2431
rect 154865 2397 154899 2431
rect 155601 2397 155635 2431
rect 156245 2397 156279 2431
rect 156613 2397 156647 2431
rect 157717 2397 157751 2431
rect 158637 2397 158671 2431
rect 159925 2397 159959 2431
rect 160017 2397 160051 2431
rect 160201 2397 160235 2431
rect 160661 2397 160695 2431
rect 161489 2397 161523 2431
rect 163697 2397 163731 2431
rect 165077 2397 165111 2431
rect 165813 2397 165847 2431
rect 166641 2397 166675 2431
rect 167929 2397 167963 2431
rect 168021 2397 168055 2431
rect 168849 2397 168883 2431
rect 169125 2397 169159 2431
rect 176669 2397 176703 2431
rect 176945 2397 176979 2431
rect 179613 2397 179647 2431
rect 179889 2397 179923 2431
rect 181821 2397 181855 2431
rect 184765 2397 184799 2431
rect 186973 2397 187007 2431
rect 190377 2397 190411 2431
rect 191849 2397 191883 2431
rect 194701 2397 194735 2431
rect 196173 2397 196207 2431
rect 197001 2397 197035 2431
rect 197829 2397 197863 2431
rect 198565 2397 198599 2431
rect 200221 2397 200255 2431
rect 201049 2397 201083 2431
rect 201785 2397 201819 2431
rect 203165 2397 203199 2431
rect 203257 2397 203291 2431
rect 203441 2397 203475 2431
rect 203901 2397 203935 2431
rect 208317 2397 208351 2431
rect 208869 2397 208903 2431
rect 208961 2397 208995 2431
rect 209145 2397 209179 2431
rect 209513 2397 209547 2431
rect 212365 2397 212399 2431
rect 214205 2397 214239 2431
rect 215217 2397 215251 2431
rect 217701 2397 217735 2431
rect 218437 2397 218471 2431
rect 218575 2397 218609 2431
rect 218713 2397 218747 2431
rect 220553 2397 220587 2431
rect 220645 2397 220679 2431
rect 220737 2397 220771 2431
rect 221381 2397 221415 2431
rect 224049 2397 224083 2431
rect 224969 2397 225003 2431
rect 225521 2397 225555 2431
rect 226257 2397 226291 2431
rect 227177 2397 227211 2431
rect 227821 2397 227855 2431
rect 229845 2397 229879 2431
rect 231409 2397 231443 2431
rect 232237 2397 232271 2431
rect 232973 2397 233007 2431
rect 234997 2397 235031 2431
rect 235825 2397 235859 2431
rect 236009 2397 236043 2431
rect 236653 2397 236687 2431
rect 243461 2397 243495 2431
rect 243737 2397 243771 2431
rect 244749 2397 244783 2431
rect 245025 2397 245059 2431
rect 248797 2397 248831 2431
rect 251281 2397 251315 2431
rect 253581 2397 253615 2431
rect 254869 2397 254903 2431
rect 255145 2397 255179 2431
rect 256433 2397 256467 2431
rect 258733 2397 258767 2431
rect 259009 2397 259043 2431
rect 261769 2397 261803 2431
rect 261953 2397 261987 2431
rect 262413 2397 262447 2431
rect 263149 2397 263183 2431
rect 264161 2397 264195 2431
rect 265173 2397 265207 2431
rect 266737 2397 266771 2431
rect 267841 2397 267875 2431
rect 268485 2397 268519 2431
rect 268945 2397 268979 2431
rect 269129 2397 269163 2431
rect 269957 2397 269991 2431
rect 270601 2397 270635 2431
rect 32965 2329 32999 2363
rect 38485 2329 38519 2363
rect 40601 2329 40635 2363
rect 42625 2329 42659 2363
rect 60749 2329 60783 2363
rect 92397 2329 92431 2363
rect 99021 2329 99055 2363
rect 103805 2329 103839 2363
rect 112361 2329 112395 2363
rect 116685 2329 116719 2363
rect 143273 2329 143307 2363
rect 144929 2329 144963 2363
rect 157073 2329 157107 2363
rect 159005 2329 159039 2363
rect 162317 2329 162351 2363
rect 191205 2329 191239 2363
rect 210249 2329 210283 2363
rect 211905 2329 211939 2363
rect 220921 2329 220955 2363
rect 221565 2329 221599 2363
rect 230765 2329 230799 2363
rect 246313 2329 246347 2363
rect 247969 2329 248003 2363
rect 253121 2329 253155 2363
rect 260113 2329 260147 2363
rect 22937 2261 22971 2295
rect 25697 2261 25731 2295
rect 29929 2261 29963 2295
rect 32229 2261 32263 2295
rect 38117 2261 38151 2295
rect 39221 2261 39255 2295
rect 39405 2261 39439 2295
rect 40233 2261 40267 2295
rect 41337 2261 41371 2295
rect 41521 2261 41555 2295
rect 42257 2261 42291 2295
rect 43361 2261 43395 2295
rect 54401 2261 54435 2295
rect 57989 2261 58023 2295
rect 59461 2261 59495 2295
rect 60841 2261 60875 2295
rect 61669 2261 61703 2295
rect 62405 2261 62439 2295
rect 63141 2261 63175 2295
rect 65993 2261 66027 2295
rect 88533 2261 88567 2295
rect 89269 2261 89303 2295
rect 90189 2261 90223 2295
rect 90925 2261 90959 2295
rect 93041 2261 93075 2295
rect 93777 2261 93811 2295
rect 117329 2261 117363 2295
rect 117973 2261 118007 2295
rect 118617 2261 118651 2295
rect 122665 2261 122699 2295
rect 125149 2261 125183 2295
rect 126253 2261 126287 2295
rect 126989 2261 127023 2295
rect 128461 2261 128495 2295
rect 129197 2261 129231 2295
rect 130761 2261 130795 2295
rect 131681 2261 131715 2295
rect 133245 2261 133279 2295
rect 134993 2261 135027 2295
rect 142169 2261 142203 2295
rect 154037 2261 154071 2295
rect 157901 2261 157935 2295
rect 160845 2261 160879 2295
rect 161673 2261 161707 2295
rect 162409 2261 162443 2295
rect 163881 2261 163915 2295
rect 165261 2261 165295 2295
rect 165997 2261 166031 2295
rect 166825 2261 166859 2295
rect 168205 2261 168239 2295
rect 191297 2261 191331 2295
rect 194885 2261 194919 2295
rect 196357 2261 196391 2295
rect 197185 2261 197219 2295
rect 198013 2261 198047 2295
rect 201233 2261 201267 2295
rect 204085 2261 204119 2295
rect 208133 2261 208167 2295
rect 224233 2261 224267 2295
rect 224785 2261 224819 2295
rect 225705 2261 225739 2295
rect 226441 2261 226475 2295
rect 228005 2261 228039 2295
rect 230029 2261 230063 2295
rect 231593 2261 231627 2295
rect 232421 2261 232455 2295
rect 233157 2261 233191 2295
rect 235181 2261 235215 2295
rect 236193 2261 236227 2295
rect 236837 2261 236871 2295
rect 260205 2261 260239 2295
rect 263333 2261 263367 2295
rect 264345 2261 264379 2295
rect 266921 2261 266955 2295
rect 267657 2261 267691 2295
rect 269313 2261 269347 2295
rect 270785 2261 270819 2295
rect 1777 2057 1811 2091
rect 12081 2057 12115 2091
rect 12817 2057 12851 2091
rect 37933 2057 37967 2091
rect 89269 2057 89303 2091
rect 90281 2057 90315 2091
rect 91109 2057 91143 2091
rect 91937 2057 91971 2091
rect 93593 2057 93627 2091
rect 94605 2057 94639 2091
rect 96445 2057 96479 2091
rect 98745 2057 98779 2091
rect 112545 2057 112579 2091
rect 114017 2057 114051 2091
rect 116869 2057 116903 2091
rect 119353 2057 119387 2091
rect 121101 2057 121135 2091
rect 124321 2057 124355 2091
rect 126713 2057 126747 2091
rect 128369 2057 128403 2091
rect 133705 2057 133739 2091
rect 139593 2057 139627 2091
rect 142353 2057 142387 2091
rect 144653 2057 144687 2091
rect 147505 2057 147539 2091
rect 149805 2057 149839 2091
rect 152657 2057 152691 2091
rect 153117 2057 153151 2091
rect 153761 2057 153795 2091
rect 154405 2057 154439 2091
rect 155049 2057 155083 2091
rect 159465 2057 159499 2091
rect 160293 2057 160327 2091
rect 162317 2057 162351 2091
rect 163973 2057 164007 2091
rect 165629 2057 165663 2091
rect 166641 2057 166675 2091
rect 167469 2057 167503 2091
rect 190929 2057 190963 2091
rect 192217 2057 192251 2091
rect 197553 2057 197587 2091
rect 199761 2057 199795 2091
rect 216781 2057 216815 2091
rect 219633 2057 219667 2091
rect 221933 2057 221967 2091
rect 222945 2057 222979 2091
rect 224141 2057 224175 2091
rect 224509 2057 224543 2091
rect 225797 2057 225831 2091
rect 226809 2057 226843 2091
rect 228465 2057 228499 2091
rect 230949 2057 230983 2091
rect 231777 2057 231811 2091
rect 232605 2057 232639 2091
rect 233617 2057 233651 2091
rect 236101 2057 236135 2091
rect 236929 2057 236963 2091
rect 241483 2057 241517 2091
rect 260573 2057 260607 2091
rect 261677 2057 261711 2091
rect 263333 2057 263367 2091
rect 25881 1989 25915 2023
rect 39129 1989 39163 2023
rect 39405 1989 39439 2023
rect 39497 1989 39531 2023
rect 39865 1989 39899 2023
rect 40233 1989 40267 2023
rect 53297 1989 53331 2023
rect 54033 1989 54067 2023
rect 57529 1989 57563 2023
rect 59185 1989 59219 2023
rect 61669 1989 61703 2023
rect 62681 1989 62715 2023
rect 65441 1989 65475 2023
rect 89545 1989 89579 2023
rect 99481 1989 99515 2023
rect 101137 1989 101171 2023
rect 103713 1989 103747 2023
rect 107393 1989 107427 2023
rect 117237 1989 117271 2023
rect 131773 1989 131807 2023
rect 158361 1989 158395 2023
rect 201417 1989 201451 2023
rect 202705 1989 202739 2023
rect 211997 1989 212031 2023
rect 214481 1989 214515 2023
rect 226073 1989 226107 2023
rect 245025 1989 245059 2023
rect 255697 1989 255731 2023
rect 257353 1989 257387 2023
rect 1685 1921 1719 1955
rect 4077 1921 4111 1955
rect 7389 1921 7423 1955
rect 8677 1921 8711 1955
rect 11989 1921 12023 1955
rect 12725 1921 12759 1955
rect 14381 1921 14415 1955
rect 15761 1921 15795 1955
rect 17877 1921 17911 1955
rect 18061 1921 18095 1955
rect 21189 1921 21223 1955
rect 22293 1921 22327 1955
rect 23305 1921 23339 1955
rect 23489 1921 23523 1955
rect 24041 1921 24075 1955
rect 24961 1921 24995 1955
rect 27905 1921 27939 1955
rect 28733 1921 28767 1955
rect 29561 1921 29595 1955
rect 30205 1921 30239 1955
rect 31217 1921 31251 1955
rect 32505 1921 32539 1955
rect 33149 1921 33183 1955
rect 38117 1921 38151 1955
rect 45477 1921 45511 1955
rect 52745 1921 52779 1955
rect 53849 1921 53883 1955
rect 54861 1921 54895 1955
rect 55597 1921 55631 1955
rect 55689 1921 55723 1955
rect 56425 1921 56459 1955
rect 56517 1921 56551 1955
rect 57161 1921 57195 1955
rect 57345 1921 57379 1955
rect 58081 1921 58115 1955
rect 58817 1921 58851 1955
rect 59001 1921 59035 1955
rect 59737 1921 59771 1955
rect 59829 1921 59863 1955
rect 60565 1921 60599 1955
rect 60657 1921 60691 1955
rect 61301 1921 61335 1955
rect 61485 1921 61519 1955
rect 62313 1921 62347 1955
rect 62497 1921 62531 1955
rect 63417 1921 63451 1955
rect 63601 1921 63635 1955
rect 64061 1921 64095 1955
rect 64245 1921 64279 1955
rect 65257 1921 65291 1955
rect 66361 1921 66395 1955
rect 66453 1921 66487 1955
rect 66637 1921 66671 1955
rect 67097 1921 67131 1955
rect 71513 1921 71547 1955
rect 72249 1921 72283 1955
rect 73721 1921 73755 1955
rect 79701 1921 79735 1955
rect 81173 1921 81207 1955
rect 84853 1921 84887 1955
rect 86325 1921 86359 1955
rect 88165 1921 88199 1955
rect 89085 1921 89119 1955
rect 90097 1921 90131 1955
rect 90833 1921 90867 1955
rect 90925 1921 90959 1955
rect 91661 1921 91695 1955
rect 91753 1921 91787 1955
rect 92581 1921 92615 1955
rect 93225 1921 93259 1955
rect 93409 1921 93443 1955
rect 94237 1921 94271 1955
rect 94421 1921 94455 1955
rect 95433 1921 95467 1955
rect 96077 1921 96111 1955
rect 96261 1921 96295 1955
rect 96905 1921 96939 1955
rect 97843 1921 97877 1955
rect 97942 1921 97976 1955
rect 98101 1921 98135 1955
rect 101873 1921 101907 1955
rect 104909 1921 104943 1955
rect 105829 1921 105863 1955
rect 105967 1921 106001 1955
rect 106105 1921 106139 1955
rect 109601 1921 109635 1955
rect 110705 1921 110739 1955
rect 111901 1921 111935 1955
rect 113557 1921 113591 1955
rect 114201 1921 114235 1955
rect 115949 1921 115983 1955
rect 116066 1921 116100 1955
rect 116225 1921 116259 1955
rect 117513 1921 117547 1955
rect 117697 1921 117731 1955
rect 118433 1921 118467 1955
rect 120089 1921 120123 1955
rect 120733 1921 120767 1955
rect 121469 1921 121503 1955
rect 121653 1921 121687 1955
rect 122297 1921 122331 1955
rect 123309 1921 123343 1955
rect 124137 1921 124171 1955
rect 125425 1921 125459 1955
rect 125609 1921 125643 1955
rect 126345 1921 126379 1955
rect 126529 1921 126563 1955
rect 127357 1921 127391 1955
rect 128001 1921 128035 1955
rect 128185 1921 128219 1955
rect 128829 1921 128863 1955
rect 130485 1921 130519 1955
rect 130669 1921 130703 1955
rect 131405 1921 131439 1955
rect 131589 1921 131623 1955
rect 132325 1921 132359 1955
rect 132509 1921 132543 1955
rect 133337 1921 133371 1955
rect 133521 1921 133555 1955
rect 134349 1921 134383 1955
rect 135361 1921 135395 1955
rect 138489 1921 138523 1955
rect 139133 1921 139167 1955
rect 139777 1921 139811 1955
rect 140513 1921 140547 1955
rect 141433 1921 141467 1955
rect 141709 1921 141743 1955
rect 142813 1921 142847 1955
rect 143733 1921 143767 1955
rect 143871 1921 143905 1955
rect 145665 1921 145699 1955
rect 146585 1921 146619 1955
rect 147965 1921 147999 1955
rect 150817 1921 150851 1955
rect 151737 1921 151771 1955
rect 152013 1921 152047 1955
rect 153301 1921 153335 1955
rect 153945 1921 153979 1955
rect 154589 1921 154623 1955
rect 155233 1921 155267 1955
rect 155785 1921 155819 1955
rect 156429 1921 156463 1955
rect 156797 1921 156831 1955
rect 157993 1921 158027 1955
rect 159097 1921 159131 1955
rect 159281 1921 159315 1955
rect 160109 1921 160143 1955
rect 161121 1921 161155 1955
rect 161305 1921 161339 1955
rect 161949 1921 161983 1955
rect 162133 1921 162167 1955
rect 162777 1921 162811 1955
rect 162961 1921 162995 1955
rect 163605 1921 163639 1955
rect 163789 1921 163823 1955
rect 164525 1921 164559 1955
rect 164617 1921 164651 1955
rect 165261 1921 165295 1955
rect 165445 1921 165479 1955
rect 166273 1921 166307 1955
rect 166457 1921 166491 1955
rect 167101 1921 167135 1955
rect 167285 1921 167319 1955
rect 168113 1921 168147 1955
rect 168297 1921 168331 1955
rect 168757 1921 168791 1955
rect 173265 1921 173299 1955
rect 176853 1921 176887 1955
rect 179429 1921 179463 1955
rect 183293 1921 183327 1955
rect 184581 1921 184615 1955
rect 187157 1921 187191 1955
rect 188445 1921 188479 1955
rect 190285 1921 190319 1955
rect 190561 1921 190595 1955
rect 190745 1921 190779 1955
rect 192033 1921 192067 1955
rect 193045 1921 193079 1955
rect 193689 1921 193723 1955
rect 193873 1921 193907 1955
rect 194701 1921 194735 1955
rect 195345 1921 195379 1955
rect 195529 1921 195563 1955
rect 195713 1921 195747 1955
rect 196173 1921 196207 1955
rect 196357 1921 196391 1955
rect 197185 1921 197219 1955
rect 197369 1921 197403 1955
rect 199393 1921 199427 1955
rect 199577 1921 199611 1955
rect 200313 1921 200347 1955
rect 200405 1921 200439 1955
rect 201049 1921 201083 1955
rect 201233 1921 201267 1955
rect 202337 1921 202371 1955
rect 202521 1921 202555 1955
rect 203257 1921 203291 1955
rect 203349 1921 203383 1955
rect 203533 1921 203567 1955
rect 203993 1921 204027 1955
rect 207857 1921 207891 1955
rect 208501 1921 208535 1955
rect 208961 1921 208995 1955
rect 211353 1921 211387 1955
rect 211445 1921 211479 1955
rect 211629 1921 211663 1955
rect 212641 1921 212675 1955
rect 213678 1921 213712 1955
rect 213837 1921 213871 1955
rect 214941 1921 214975 1955
rect 215861 1921 215895 1955
rect 215999 1921 216033 1955
rect 218713 1921 218747 1955
rect 218989 1921 219023 1955
rect 220277 1921 220311 1955
rect 221031 1921 221065 1955
rect 221289 1921 221323 1955
rect 223129 1921 223163 1955
rect 223957 1921 223991 1955
rect 224969 1921 225003 1955
rect 225613 1921 225647 1955
rect 226625 1921 226659 1955
rect 227269 1921 227303 1955
rect 228189 1921 228223 1955
rect 228281 1921 228315 1955
rect 228925 1921 228959 1955
rect 229109 1921 229143 1955
rect 229753 1921 229787 1955
rect 229937 1921 229971 1955
rect 230673 1921 230707 1955
rect 230765 1921 230799 1955
rect 231409 1921 231443 1955
rect 231593 1921 231627 1955
rect 232237 1921 232271 1955
rect 232421 1921 232455 1955
rect 233249 1921 233283 1955
rect 233433 1921 233467 1955
rect 234077 1921 234111 1955
rect 234261 1921 234295 1955
rect 235089 1921 235123 1955
rect 235733 1921 235767 1955
rect 235917 1921 235951 1955
rect 236561 1921 236595 1955
rect 236745 1921 236779 1955
rect 237389 1921 237423 1955
rect 243829 1921 243863 1955
rect 247417 1921 247451 1955
rect 248705 1921 248739 1955
rect 254133 1921 254167 1955
rect 255513 1921 255547 1955
rect 258089 1921 258123 1955
rect 259285 1921 259319 1955
rect 260481 1921 260515 1955
rect 261493 1921 261527 1955
rect 262137 1921 262171 1955
rect 262321 1921 262355 1955
rect 262965 1921 262999 1955
rect 263149 1921 263183 1955
rect 264161 1921 264195 1955
rect 264345 1921 264379 1955
rect 264989 1921 265023 1955
rect 265173 1921 265207 1955
rect 265817 1921 265851 1955
rect 266001 1921 266035 1955
rect 266645 1921 266679 1955
rect 266829 1921 266863 1955
rect 267013 1921 267047 1955
rect 267473 1921 267507 1955
rect 267657 1921 267691 1955
rect 268301 1921 268335 1955
rect 268485 1921 268519 1955
rect 269405 1921 269439 1955
rect 269497 1921 269531 1955
rect 269681 1921 269715 1955
rect 270141 1921 270175 1955
rect 3801 1853 3835 1887
rect 5181 1853 5215 1887
rect 5457 1853 5491 1887
rect 7113 1853 7147 1887
rect 8401 1853 8435 1887
rect 9689 1853 9723 1887
rect 9965 1853 9999 1887
rect 14105 1853 14139 1887
rect 15485 1853 15519 1887
rect 22109 1853 22143 1887
rect 22845 1853 22879 1887
rect 23121 1853 23155 1887
rect 24317 1853 24351 1887
rect 27721 1853 27755 1887
rect 28549 1853 28583 1887
rect 29377 1853 29411 1887
rect 29745 1853 29779 1887
rect 30021 1853 30055 1887
rect 30757 1853 30791 1887
rect 31033 1853 31067 1887
rect 32321 1853 32355 1887
rect 53665 1853 53699 1887
rect 54677 1853 54711 1887
rect 64797 1853 64831 1887
rect 65073 1853 65107 1887
rect 75745 1853 75779 1887
rect 76021 1853 76055 1887
rect 77217 1853 77251 1887
rect 77493 1853 77527 1887
rect 79425 1853 79459 1887
rect 80897 1853 80931 1887
rect 82369 1853 82403 1887
rect 82645 1853 82679 1887
rect 84577 1853 84611 1887
rect 86049 1853 86083 1887
rect 88901 1853 88935 1887
rect 89913 1853 89947 1887
rect 92397 1853 92431 1887
rect 94973 1853 95007 1887
rect 95249 1853 95283 1887
rect 97089 1853 97123 1887
rect 99297 1853 99331 1887
rect 102057 1853 102091 1887
rect 105093 1853 105127 1887
rect 106749 1853 106783 1887
rect 107209 1853 107243 1887
rect 107669 1853 107703 1887
rect 109785 1853 109819 1887
rect 110889 1853 110923 1887
rect 111625 1853 111659 1887
rect 111763 1853 111797 1887
rect 115029 1853 115063 1887
rect 115213 1853 115247 1887
rect 118157 1853 118191 1887
rect 118550 1853 118584 1887
rect 118709 1853 118743 1887
rect 122113 1853 122147 1887
rect 122849 1853 122883 1887
rect 123125 1853 123159 1887
rect 123953 1853 123987 1887
rect 127173 1853 127207 1887
rect 129105 1853 129139 1887
rect 134165 1853 134199 1887
rect 140697 1853 140731 1887
rect 141157 1853 141191 1887
rect 141571 1853 141605 1887
rect 142997 1853 143031 1887
rect 144009 1853 144043 1887
rect 145849 1853 145883 1887
rect 146723 1853 146757 1887
rect 146861 1853 146895 1887
rect 148149 1853 148183 1887
rect 148609 1853 148643 1887
rect 148885 1853 148919 1887
rect 149002 1853 149036 1887
rect 149161 1853 149195 1887
rect 151001 1853 151035 1887
rect 151875 1853 151909 1887
rect 157073 1853 157107 1887
rect 159925 1853 159959 1887
rect 167929 1853 167963 1887
rect 172989 1853 173023 1887
rect 174461 1853 174495 1887
rect 174737 1853 174771 1887
rect 176577 1853 176611 1887
rect 177865 1853 177899 1887
rect 178141 1853 178175 1887
rect 179153 1853 179187 1887
rect 181729 1853 181763 1887
rect 182005 1853 182039 1887
rect 183017 1853 183051 1887
rect 184305 1853 184339 1887
rect 186881 1853 186915 1887
rect 188169 1853 188203 1887
rect 191849 1853 191883 1887
rect 192585 1853 192619 1887
rect 192861 1853 192895 1887
rect 194517 1853 194551 1887
rect 198105 1853 198139 1887
rect 198381 1853 198415 1887
rect 209145 1853 209179 1887
rect 209789 1853 209823 1887
rect 212825 1853 212859 1887
rect 213285 1853 213319 1887
rect 213561 1853 213595 1887
rect 215125 1853 215159 1887
rect 216137 1853 216171 1887
rect 217793 1853 217827 1887
rect 217977 1853 218011 1887
rect 218851 1853 218885 1887
rect 220093 1853 220127 1887
rect 220737 1853 220771 1887
rect 221130 1853 221164 1887
rect 223773 1853 223807 1887
rect 224785 1853 224819 1887
rect 225429 1853 225463 1887
rect 226441 1853 226475 1887
rect 234905 1853 234939 1887
rect 241253 1853 241287 1887
rect 243553 1853 243587 1887
rect 244841 1853 244875 1887
rect 246681 1853 246715 1887
rect 247141 1853 247175 1887
rect 248889 1853 248923 1887
rect 250545 1853 250579 1887
rect 251005 1853 251039 1887
rect 251281 1853 251315 1887
rect 252293 1853 252327 1887
rect 252569 1853 252603 1887
rect 253857 1853 253891 1887
rect 259009 1853 259043 1887
rect 261309 1853 261343 1887
rect 45293 1785 45327 1819
rect 71329 1785 71363 1819
rect 72065 1785 72099 1819
rect 73537 1785 73571 1819
rect 97549 1785 97583 1819
rect 105553 1785 105587 1819
rect 111349 1785 111383 1819
rect 113373 1785 113407 1819
rect 115673 1785 115707 1819
rect 138949 1785 138983 1819
rect 143457 1785 143491 1819
rect 146309 1785 146343 1819
rect 151461 1785 151495 1819
rect 207673 1785 207707 1819
rect 215585 1785 215619 1819
rect 218437 1785 218471 1819
rect 21373 1717 21407 1751
rect 22477 1717 22511 1751
rect 23765 1717 23799 1751
rect 25053 1717 25087 1751
rect 25973 1717 26007 1751
rect 28089 1717 28123 1751
rect 28917 1717 28951 1751
rect 30389 1717 30423 1751
rect 31401 1717 31435 1751
rect 32689 1717 32723 1751
rect 33333 1717 33367 1751
rect 35173 1717 35207 1751
rect 40417 1717 40451 1751
rect 52929 1717 52963 1751
rect 54309 1717 54343 1751
rect 55045 1717 55079 1751
rect 55873 1717 55907 1751
rect 56701 1717 56735 1751
rect 58265 1717 58299 1751
rect 60013 1717 60047 1751
rect 60841 1717 60875 1751
rect 63785 1717 63819 1751
rect 64429 1717 64463 1751
rect 67281 1717 67315 1751
rect 88349 1717 88383 1751
rect 92765 1717 92799 1751
rect 95617 1717 95651 1751
rect 119905 1717 119939 1751
rect 120549 1717 120583 1751
rect 121837 1717 121871 1751
rect 122481 1717 122515 1751
rect 123493 1717 123527 1751
rect 125793 1717 125827 1751
rect 127541 1717 127575 1751
rect 130853 1717 130887 1751
rect 132693 1717 132727 1751
rect 134533 1717 134567 1751
rect 135545 1717 135579 1751
rect 138305 1717 138339 1751
rect 155969 1717 156003 1751
rect 161489 1717 161523 1751
rect 163145 1717 163179 1751
rect 164801 1717 164835 1751
rect 168941 1717 168975 1751
rect 193229 1717 193263 1751
rect 194057 1717 194091 1751
rect 194885 1717 194919 1751
rect 196541 1717 196575 1751
rect 200589 1717 200623 1751
rect 204177 1717 204211 1751
rect 208317 1717 208351 1751
rect 223405 1717 223439 1751
rect 225153 1717 225187 1751
rect 227453 1717 227487 1751
rect 229293 1717 229327 1751
rect 230121 1717 230155 1751
rect 234445 1717 234479 1751
rect 235273 1717 235307 1751
rect 237573 1717 237607 1751
rect 257629 1717 257663 1751
rect 258181 1717 258215 1751
rect 262505 1717 262539 1751
rect 264529 1717 264563 1751
rect 265357 1717 265391 1751
rect 266185 1717 266219 1751
rect 267841 1717 267875 1751
rect 268669 1717 268703 1751
rect 270325 1717 270359 1751
rect 27537 1513 27571 1547
rect 58725 1513 58759 1547
rect 62405 1513 62439 1547
rect 95341 1513 95375 1547
rect 98561 1513 98595 1547
rect 117421 1513 117455 1547
rect 118525 1513 118559 1547
rect 120181 1513 120215 1547
rect 126529 1513 126563 1547
rect 129289 1513 129323 1547
rect 142169 1513 142203 1547
rect 144929 1513 144963 1547
rect 151461 1513 151495 1547
rect 156797 1513 156831 1547
rect 220369 1513 220403 1547
rect 247325 1513 247359 1547
rect 96077 1445 96111 1479
rect 97365 1445 97399 1479
rect 100309 1445 100343 1479
rect 105277 1445 105311 1479
rect 107853 1445 107887 1479
rect 109049 1445 109083 1479
rect 110429 1445 110463 1479
rect 112821 1445 112855 1479
rect 115581 1445 115615 1479
rect 133521 1445 133555 1479
rect 138121 1445 138155 1479
rect 140973 1445 141007 1479
rect 146953 1445 146987 1479
rect 148885 1445 148919 1479
rect 196633 1445 196667 1479
rect 198289 1445 198323 1479
rect 210709 1445 210743 1479
rect 22845 1377 22879 1411
rect 23673 1377 23707 1411
rect 25053 1377 25087 1411
rect 25881 1377 25915 1411
rect 27169 1377 27203 1411
rect 54309 1377 54343 1411
rect 58357 1377 58391 1411
rect 62037 1377 62071 1411
rect 65993 1377 66027 1411
rect 69121 1377 69155 1411
rect 89085 1377 89119 1411
rect 90557 1377 90591 1411
rect 94145 1377 94179 1411
rect 94973 1377 95007 1411
rect 95433 1377 95467 1411
rect 97641 1377 97675 1411
rect 99205 1377 99239 1411
rect 100585 1377 100619 1411
rect 100723 1377 100757 1411
rect 105829 1377 105863 1411
rect 108405 1377 108439 1411
rect 110705 1377 110739 1411
rect 113373 1377 113407 1411
rect 115995 1377 116029 1411
rect 126161 1377 126195 1411
rect 128921 1377 128955 1411
rect 133153 1377 133187 1411
rect 141525 1377 141559 1411
rect 143733 1377 143767 1411
rect 144285 1377 144319 1411
rect 158545 1377 158579 1411
rect 159373 1377 159407 1411
rect 162685 1377 162719 1411
rect 166917 1377 166951 1411
rect 171701 1377 171735 1411
rect 190653 1377 190687 1411
rect 190929 1377 190963 1411
rect 196265 1377 196299 1411
rect 197921 1377 197955 1411
rect 201325 1377 201359 1411
rect 202889 1377 202923 1411
rect 205833 1377 205867 1411
rect 211261 1377 211295 1411
rect 213101 1377 213135 1411
rect 213653 1377 213687 1411
rect 215861 1377 215895 1411
rect 224417 1377 224451 1411
rect 226901 1377 226935 1411
rect 227269 1377 227303 1411
rect 231317 1377 231351 1411
rect 235825 1377 235859 1411
rect 239965 1377 239999 1411
rect 246129 1377 246163 1411
rect 247509 1377 247543 1411
rect 260297 1377 260331 1411
rect 261585 1377 261619 1411
rect 269313 1377 269347 1411
rect 2605 1309 2639 1343
rect 2881 1309 2915 1343
rect 5181 1309 5215 1343
rect 5457 1309 5491 1343
rect 7757 1309 7791 1343
rect 8033 1309 8067 1343
rect 10333 1309 10367 1343
rect 10609 1309 10643 1343
rect 11713 1309 11747 1343
rect 11989 1309 12023 1343
rect 15485 1309 15519 1343
rect 15761 1309 15795 1343
rect 17049 1309 17083 1343
rect 17325 1309 17359 1343
rect 22109 1309 22143 1343
rect 23029 1309 23063 1343
rect 23213 1309 23247 1343
rect 23857 1309 23891 1343
rect 24041 1309 24075 1343
rect 25237 1309 25271 1343
rect 25421 1309 25455 1343
rect 26065 1309 26099 1343
rect 26249 1309 26283 1343
rect 27353 1309 27387 1343
rect 27997 1309 28031 1343
rect 28825 1309 28859 1343
rect 30297 1309 30331 1343
rect 31033 1309 31067 1343
rect 32321 1309 32355 1343
rect 35633 1309 35667 1343
rect 36277 1309 36311 1343
rect 36921 1309 36955 1343
rect 38209 1309 38243 1343
rect 38853 1309 38887 1343
rect 39497 1309 39531 1343
rect 40785 1309 40819 1343
rect 41429 1309 41463 1343
rect 42073 1309 42107 1343
rect 43269 1309 43303 1343
rect 44005 1309 44039 1343
rect 44649 1309 44683 1343
rect 45937 1309 45971 1343
rect 46581 1309 46615 1343
rect 47225 1309 47259 1343
rect 48421 1309 48455 1343
rect 49157 1309 49191 1343
rect 49801 1309 49835 1343
rect 50629 1309 50663 1343
rect 51365 1309 51399 1343
rect 52101 1309 52135 1343
rect 53113 1309 53147 1343
rect 54493 1309 54527 1343
rect 54677 1309 54711 1343
rect 55505 1309 55539 1343
rect 56241 1309 56275 1343
rect 56977 1309 57011 1343
rect 58541 1309 58575 1343
rect 59829 1309 59863 1343
rect 60749 1309 60783 1343
rect 62221 1309 62255 1343
rect 63693 1309 63727 1343
rect 64429 1309 64463 1343
rect 66177 1309 66211 1343
rect 66361 1309 66395 1343
rect 66821 1309 66855 1343
rect 69581 1309 69615 1343
rect 69857 1309 69891 1343
rect 70961 1309 70995 1343
rect 71237 1309 71271 1343
rect 72985 1309 73019 1343
rect 74273 1309 74307 1343
rect 74733 1309 74767 1343
rect 75009 1309 75043 1343
rect 77309 1309 77343 1343
rect 77585 1309 77619 1343
rect 79885 1309 79919 1343
rect 80161 1309 80195 1343
rect 82461 1309 82495 1343
rect 82737 1309 82771 1343
rect 85037 1309 85071 1343
rect 85313 1309 85347 1343
rect 86785 1309 86819 1343
rect 87061 1309 87095 1343
rect 88165 1309 88199 1343
rect 89269 1309 89303 1343
rect 90741 1309 90775 1343
rect 90925 1309 90959 1343
rect 91661 1309 91695 1343
rect 92397 1309 92431 1343
rect 93225 1309 93259 1343
rect 93317 1309 93351 1343
rect 93501 1309 93535 1343
rect 94329 1309 94363 1343
rect 95157 1309 95191 1343
rect 95617 1309 95651 1343
rect 96721 1309 96755 1343
rect 96905 1309 96939 1343
rect 97779 1309 97813 1343
rect 97917 1309 97951 1343
rect 98653 1309 98687 1343
rect 99389 1309 99423 1343
rect 99665 1309 99699 1343
rect 99849 1309 99883 1343
rect 100861 1309 100895 1343
rect 101505 1309 101539 1343
rect 101689 1309 101723 1343
rect 104633 1309 104667 1343
rect 104817 1309 104851 1343
rect 105553 1309 105587 1343
rect 105691 1309 105725 1343
rect 106473 1309 106507 1343
rect 107209 1309 107243 1343
rect 107393 1309 107427 1343
rect 108129 1309 108163 1343
rect 108267 1309 108301 1343
rect 109785 1309 109819 1343
rect 109969 1309 110003 1343
rect 110822 1309 110856 1343
rect 110981 1309 111015 1343
rect 111625 1309 111659 1343
rect 112177 1309 112211 1343
rect 112361 1309 112395 1343
rect 113097 1309 113131 1343
rect 113235 1309 113269 1343
rect 114937 1309 114971 1343
rect 115121 1309 115155 1343
rect 115857 1309 115891 1343
rect 116133 1309 116167 1343
rect 116777 1309 116811 1343
rect 118065 1309 118099 1343
rect 118709 1309 118743 1343
rect 119353 1309 119387 1343
rect 120365 1309 120399 1343
rect 121101 1309 121135 1343
rect 121653 1309 121687 1343
rect 122481 1309 122515 1343
rect 123217 1309 123251 1343
rect 124229 1309 124263 1343
rect 125425 1309 125459 1343
rect 126345 1309 126379 1343
rect 127633 1309 127667 1343
rect 129105 1309 129139 1343
rect 130669 1309 130703 1343
rect 131957 1309 131991 1343
rect 133337 1309 133371 1343
rect 134349 1309 134383 1343
rect 138765 1309 138799 1343
rect 139409 1309 139443 1343
rect 140329 1309 140363 1343
rect 140513 1309 140547 1343
rect 141249 1309 141283 1343
rect 141387 1309 141421 1343
rect 142537 1309 142571 1343
rect 143089 1309 143123 1343
rect 143273 1309 143307 1343
rect 144009 1309 144043 1343
rect 144126 1309 144160 1343
rect 145849 1309 145883 1343
rect 146493 1309 146527 1343
rect 147137 1309 147171 1343
rect 148241 1309 148275 1343
rect 148425 1309 148459 1343
rect 149161 1309 149195 1343
rect 149299 1309 149333 1343
rect 149437 1309 149471 1343
rect 150081 1309 150115 1343
rect 151001 1309 151035 1343
rect 151645 1309 151679 1343
rect 152289 1309 152323 1343
rect 153577 1309 153611 1343
rect 154221 1309 154255 1343
rect 154865 1309 154899 1343
rect 156429 1309 156463 1343
rect 156613 1309 156647 1343
rect 157257 1309 157291 1343
rect 157441 1309 157475 1343
rect 158729 1309 158763 1343
rect 159557 1309 159591 1343
rect 159741 1309 159775 1343
rect 160201 1309 160235 1343
rect 161121 1309 161155 1343
rect 161949 1309 161983 1343
rect 162869 1309 162903 1343
rect 163053 1309 163087 1343
rect 163697 1309 163731 1343
rect 164433 1309 164467 1343
rect 167101 1309 167135 1343
rect 167285 1309 167319 1343
rect 167745 1309 167779 1343
rect 168849 1309 168883 1343
rect 172253 1309 172287 1343
rect 172529 1309 172563 1343
rect 174001 1309 174035 1343
rect 174277 1309 174311 1343
rect 176577 1309 176611 1343
rect 176853 1309 176887 1343
rect 179153 1309 179187 1343
rect 179429 1309 179463 1343
rect 181729 1309 181763 1343
rect 182005 1309 182039 1343
rect 184305 1309 184339 1343
rect 184581 1309 184615 1343
rect 186881 1309 186915 1343
rect 187157 1309 187191 1343
rect 188629 1309 188663 1343
rect 189457 1309 189491 1343
rect 189733 1309 189767 1343
rect 191113 1309 191147 1343
rect 191297 1309 191331 1343
rect 192401 1309 192435 1343
rect 193137 1309 193171 1343
rect 194609 1309 194643 1343
rect 195437 1309 195471 1343
rect 196449 1309 196483 1343
rect 198105 1309 198139 1343
rect 199761 1309 199795 1343
rect 201509 1309 201543 1343
rect 203073 1309 203107 1343
rect 203257 1309 203291 1343
rect 203717 1309 203751 1343
rect 206569 1309 206603 1343
rect 207673 1309 207707 1343
rect 208317 1309 208351 1343
rect 208961 1309 208995 1343
rect 210065 1309 210099 1343
rect 210249 1309 210283 1343
rect 210985 1309 211019 1343
rect 211102 1309 211136 1343
rect 212457 1309 212491 1343
rect 212641 1309 212675 1343
rect 213377 1309 213411 1343
rect 213515 1309 213549 1343
rect 215217 1309 215251 1343
rect 215401 1309 215435 1343
rect 216137 1309 216171 1343
rect 216275 1309 216309 1343
rect 216413 1309 216447 1343
rect 217885 1309 217919 1343
rect 217977 1309 218011 1343
rect 218069 1309 218103 1343
rect 218897 1309 218931 1343
rect 219541 1309 219575 1343
rect 220553 1309 220587 1343
rect 221657 1309 221691 1343
rect 221749 1309 221783 1343
rect 221933 1309 221967 1343
rect 223129 1309 223163 1343
rect 224233 1309 224267 1343
rect 225521 1309 225555 1343
rect 226441 1309 226475 1343
rect 227085 1309 227119 1343
rect 228557 1309 228591 1343
rect 229293 1309 229327 1343
rect 231501 1309 231535 1343
rect 231685 1309 231719 1343
rect 232145 1309 232179 1343
rect 233709 1309 233743 1343
rect 234445 1309 234479 1343
rect 236009 1309 236043 1343
rect 236193 1309 236227 1343
rect 236653 1309 236687 1343
rect 240977 1309 241011 1343
rect 241253 1309 241287 1343
rect 243553 1309 243587 1343
rect 243829 1309 243863 1343
rect 245485 1309 245519 1343
rect 246405 1309 246439 1343
rect 247325 1309 247359 1343
rect 247601 1309 247635 1343
rect 248797 1309 248831 1343
rect 251281 1309 251315 1343
rect 251557 1309 251591 1343
rect 252753 1309 252787 1343
rect 253857 1309 253891 1343
rect 254133 1309 254167 1343
rect 255605 1309 255639 1343
rect 256433 1309 256467 1343
rect 256709 1309 256743 1343
rect 257997 1309 258031 1343
rect 258181 1309 258215 1343
rect 259009 1309 259043 1343
rect 259285 1309 259319 1343
rect 260481 1309 260515 1343
rect 260665 1309 260699 1343
rect 261769 1309 261803 1343
rect 261953 1309 261987 1343
rect 262413 1309 262447 1343
rect 263149 1309 263183 1343
rect 264161 1309 264195 1343
rect 264897 1309 264931 1343
rect 265633 1309 265667 1343
rect 266737 1309 266771 1343
rect 267473 1309 267507 1343
rect 268209 1309 268243 1343
rect 269497 1309 269531 1343
rect 269681 1309 269715 1343
rect 270141 1309 270175 1343
rect 1961 1241 1995 1275
rect 13461 1241 13495 1275
rect 18613 1241 18647 1275
rect 95801 1241 95835 1275
rect 99573 1241 99607 1275
rect 157625 1241 157659 1275
rect 158913 1241 158947 1275
rect 201693 1241 201727 1275
rect 222301 1241 222335 1275
rect 248981 1241 249015 1275
rect 250637 1241 250671 1275
rect 258365 1241 258399 1275
rect 2053 1173 2087 1207
rect 13553 1173 13587 1207
rect 18705 1173 18739 1207
rect 22293 1173 22327 1207
rect 28181 1173 28215 1207
rect 29009 1173 29043 1207
rect 30481 1173 30515 1207
rect 31217 1173 31251 1207
rect 32505 1173 32539 1207
rect 35449 1173 35483 1207
rect 36093 1173 36127 1207
rect 36737 1173 36771 1207
rect 38025 1173 38059 1207
rect 38669 1173 38703 1207
rect 39313 1173 39347 1207
rect 40601 1173 40635 1207
rect 41245 1173 41279 1207
rect 41889 1173 41923 1207
rect 43085 1173 43119 1207
rect 43821 1173 43855 1207
rect 44465 1173 44499 1207
rect 45753 1173 45787 1207
rect 46397 1173 46431 1207
rect 47041 1173 47075 1207
rect 48237 1173 48271 1207
rect 48973 1173 49007 1207
rect 49617 1173 49651 1207
rect 50445 1173 50479 1207
rect 51181 1173 51215 1207
rect 51917 1173 51951 1207
rect 52929 1173 52963 1207
rect 55689 1173 55723 1207
rect 56425 1173 56459 1207
rect 57161 1173 57195 1207
rect 60013 1173 60047 1207
rect 60933 1173 60967 1207
rect 63877 1173 63911 1207
rect 64613 1173 64647 1207
rect 67005 1173 67039 1207
rect 72801 1173 72835 1207
rect 74089 1173 74123 1207
rect 88349 1173 88383 1207
rect 89453 1173 89487 1207
rect 91845 1173 91879 1207
rect 92581 1173 92615 1207
rect 94513 1173 94547 1207
rect 98837 1173 98871 1207
rect 101873 1173 101907 1207
rect 103529 1173 103563 1207
rect 103805 1173 103839 1207
rect 109601 1173 109635 1207
rect 114017 1173 114051 1207
rect 117697 1173 117731 1207
rect 117881 1173 117915 1207
rect 119169 1173 119203 1207
rect 120917 1173 120951 1207
rect 121837 1173 121871 1207
rect 122665 1173 122699 1207
rect 123401 1173 123435 1207
rect 124413 1173 124447 1207
rect 125609 1173 125643 1207
rect 127817 1173 127851 1207
rect 130853 1173 130887 1207
rect 132141 1173 132175 1207
rect 134533 1173 134567 1207
rect 138581 1173 138615 1207
rect 139225 1173 139259 1207
rect 145665 1173 145699 1207
rect 146309 1173 146343 1207
rect 150817 1173 150851 1207
rect 152105 1173 152139 1207
rect 153393 1173 153427 1207
rect 154037 1173 154071 1207
rect 154681 1173 154715 1207
rect 160385 1173 160419 1207
rect 161305 1173 161339 1207
rect 162133 1173 162167 1207
rect 163881 1173 163915 1207
rect 164617 1173 164651 1207
rect 167929 1173 167963 1207
rect 169033 1173 169067 1207
rect 188445 1173 188479 1207
rect 192585 1173 192619 1207
rect 193321 1173 193355 1207
rect 194793 1173 194827 1207
rect 195621 1173 195655 1207
rect 199945 1173 199979 1207
rect 203901 1173 203935 1207
rect 206385 1173 206419 1207
rect 207489 1173 207523 1207
rect 208133 1173 208167 1207
rect 208777 1173 208811 1207
rect 209513 1173 209547 1207
rect 211905 1173 211939 1207
rect 214297 1173 214331 1207
rect 214665 1173 214699 1207
rect 217057 1173 217091 1207
rect 218253 1173 218287 1207
rect 218713 1173 218747 1207
rect 219357 1173 219391 1207
rect 222945 1173 222979 1207
rect 225705 1173 225739 1207
rect 226257 1173 226291 1207
rect 228741 1173 228775 1207
rect 229477 1173 229511 1207
rect 232329 1173 232363 1207
rect 233893 1173 233927 1207
rect 234629 1173 234663 1207
rect 236837 1173 236871 1207
rect 245301 1173 245335 1207
rect 247785 1173 247819 1207
rect 248061 1173 248095 1207
rect 252569 1173 252603 1207
rect 255789 1173 255823 1207
rect 262597 1173 262631 1207
rect 263333 1173 263367 1207
rect 264345 1173 264379 1207
rect 265081 1173 265115 1207
rect 265817 1173 265851 1207
rect 266921 1173 266955 1207
rect 267657 1173 267691 1207
rect 268393 1173 268427 1207
rect 270325 1173 270359 1207
<< metal1 >>
rect 82078 10820 82084 10872
rect 82136 10860 82142 10872
rect 94590 10860 94596 10872
rect 82136 10832 94596 10860
rect 82136 10820 82142 10832
rect 94590 10820 94596 10832
rect 94648 10820 94654 10872
rect 94774 10820 94780 10872
rect 94832 10860 94838 10872
rect 100754 10860 100760 10872
rect 94832 10832 100760 10860
rect 94832 10820 94838 10832
rect 100754 10820 100760 10832
rect 100812 10820 100818 10872
rect 158530 10820 158536 10872
rect 158588 10860 158594 10872
rect 166442 10860 166448 10872
rect 158588 10832 166448 10860
rect 158588 10820 158594 10832
rect 166442 10820 166448 10832
rect 166500 10820 166506 10872
rect 218716 10832 219664 10860
rect 69842 10752 69848 10804
rect 69900 10792 69906 10804
rect 81526 10792 81532 10804
rect 69900 10764 81532 10792
rect 69900 10752 69906 10764
rect 81526 10752 81532 10764
rect 81584 10752 81590 10804
rect 81710 10752 81716 10804
rect 81768 10792 81774 10804
rect 93946 10792 93952 10804
rect 81768 10764 93952 10792
rect 81768 10752 81774 10764
rect 93946 10752 93952 10764
rect 94004 10752 94010 10804
rect 99190 10752 99196 10804
rect 99248 10792 99254 10804
rect 132770 10792 132776 10804
rect 99248 10764 132776 10792
rect 99248 10752 99254 10764
rect 132770 10752 132776 10764
rect 132828 10792 132834 10804
rect 133782 10792 133788 10804
rect 132828 10764 133788 10792
rect 132828 10752 132834 10764
rect 133782 10752 133788 10764
rect 133840 10752 133846 10804
rect 146570 10752 146576 10804
rect 146628 10792 146634 10804
rect 177574 10792 177580 10804
rect 146628 10764 177580 10792
rect 146628 10752 146634 10764
rect 177574 10752 177580 10764
rect 177632 10752 177638 10804
rect 92382 10684 92388 10736
rect 92440 10724 92446 10736
rect 125870 10724 125876 10736
rect 92440 10696 125876 10724
rect 92440 10684 92446 10696
rect 125870 10684 125876 10696
rect 125928 10684 125934 10736
rect 151722 10684 151728 10736
rect 151780 10724 151786 10736
rect 162762 10724 162768 10736
rect 151780 10696 162768 10724
rect 151780 10684 151786 10696
rect 162762 10684 162768 10696
rect 162820 10684 162826 10736
rect 165062 10684 165068 10736
rect 165120 10724 165126 10736
rect 217870 10724 217876 10736
rect 165120 10696 217876 10724
rect 165120 10684 165126 10696
rect 217870 10684 217876 10696
rect 217928 10684 217934 10736
rect 60642 10616 60648 10668
rect 60700 10656 60706 10668
rect 82078 10656 82084 10668
rect 60700 10628 82084 10656
rect 60700 10616 60706 10628
rect 82078 10616 82084 10628
rect 82136 10616 82142 10668
rect 94958 10616 94964 10668
rect 95016 10656 95022 10668
rect 106182 10656 106188 10668
rect 95016 10628 106188 10656
rect 95016 10616 95022 10628
rect 106182 10616 106188 10628
rect 106240 10616 106246 10668
rect 127618 10656 127624 10668
rect 109006 10628 127624 10656
rect 96430 10588 96436 10600
rect 64846 10560 96436 10588
rect 21634 10412 21640 10464
rect 21692 10452 21698 10464
rect 30650 10452 30656 10464
rect 21692 10424 30656 10452
rect 21692 10412 21698 10424
rect 30650 10412 30656 10424
rect 30708 10412 30714 10464
rect 62022 10452 62028 10464
rect 41386 10424 62028 10452
rect 27706 10344 27712 10396
rect 27764 10384 27770 10396
rect 41386 10384 41414 10424
rect 62022 10412 62028 10424
rect 62080 10452 62086 10464
rect 64846 10452 64874 10560
rect 96430 10548 96436 10560
rect 96488 10588 96494 10600
rect 98638 10588 98644 10600
rect 96488 10560 98644 10588
rect 96488 10548 96494 10560
rect 98638 10548 98644 10560
rect 98696 10548 98702 10600
rect 100018 10548 100024 10600
rect 100076 10588 100082 10600
rect 109006 10588 109034 10628
rect 127618 10616 127624 10628
rect 127676 10616 127682 10668
rect 131114 10616 131120 10668
rect 131172 10656 131178 10668
rect 131850 10656 131856 10668
rect 131172 10628 131856 10656
rect 131172 10616 131178 10628
rect 131850 10616 131856 10628
rect 131908 10656 131914 10668
rect 158530 10656 158536 10668
rect 131908 10628 158536 10656
rect 131908 10616 131914 10628
rect 158530 10616 158536 10628
rect 158588 10616 158594 10668
rect 158622 10616 158628 10668
rect 158680 10656 158686 10668
rect 164510 10656 164516 10668
rect 158680 10628 164516 10656
rect 158680 10616 158686 10628
rect 164510 10616 164516 10628
rect 164568 10616 164574 10668
rect 202322 10616 202328 10668
rect 202380 10656 202386 10668
rect 218716 10656 218744 10832
rect 219636 10724 219664 10832
rect 220170 10820 220176 10872
rect 220228 10860 220234 10872
rect 224954 10860 224960 10872
rect 220228 10832 224960 10860
rect 220228 10820 220234 10832
rect 224954 10820 224960 10832
rect 225012 10820 225018 10872
rect 230658 10860 230664 10872
rect 225064 10832 230664 10860
rect 219894 10752 219900 10804
rect 219952 10792 219958 10804
rect 225064 10792 225092 10832
rect 230658 10820 230664 10832
rect 230716 10860 230722 10872
rect 230716 10832 241514 10860
rect 230716 10820 230722 10832
rect 219952 10764 225092 10792
rect 219952 10752 219958 10764
rect 225138 10752 225144 10804
rect 225196 10792 225202 10804
rect 233602 10792 233608 10804
rect 225196 10764 233608 10792
rect 225196 10752 225202 10764
rect 233602 10752 233608 10764
rect 233660 10752 233666 10804
rect 241486 10792 241514 10832
rect 257614 10820 257620 10872
rect 257672 10860 257678 10872
rect 266906 10860 266912 10872
rect 257672 10832 266912 10860
rect 257672 10820 257678 10832
rect 266906 10820 266912 10832
rect 266964 10820 266970 10872
rect 264698 10792 264704 10804
rect 241486 10764 264704 10792
rect 264698 10752 264704 10764
rect 264756 10752 264762 10804
rect 234706 10724 234712 10736
rect 219636 10696 234712 10724
rect 234706 10684 234712 10696
rect 234764 10684 234770 10736
rect 236638 10684 236644 10736
rect 236696 10724 236702 10736
rect 263778 10724 263784 10736
rect 236696 10696 263784 10724
rect 236696 10684 236702 10696
rect 263778 10684 263784 10696
rect 263836 10684 263842 10736
rect 202380 10628 218744 10656
rect 202380 10616 202386 10628
rect 218790 10616 218796 10668
rect 218848 10656 218854 10668
rect 226702 10656 226708 10668
rect 218848 10628 226708 10656
rect 218848 10616 218854 10628
rect 226702 10616 226708 10628
rect 226760 10616 226766 10668
rect 226978 10616 226984 10668
rect 227036 10656 227042 10668
rect 229094 10656 229100 10668
rect 227036 10628 229100 10656
rect 227036 10616 227042 10628
rect 229094 10616 229100 10628
rect 229152 10616 229158 10668
rect 258534 10616 258540 10668
rect 258592 10656 258598 10668
rect 267550 10656 267556 10668
rect 258592 10628 267556 10656
rect 258592 10616 258598 10628
rect 267550 10616 267556 10628
rect 267608 10616 267614 10668
rect 100076 10560 109034 10588
rect 100076 10548 100082 10560
rect 148686 10548 148692 10600
rect 148744 10588 148750 10600
rect 180702 10588 180708 10600
rect 148744 10560 180708 10588
rect 148744 10548 148750 10560
rect 180702 10548 180708 10560
rect 180760 10548 180766 10600
rect 200114 10548 200120 10600
rect 200172 10588 200178 10600
rect 228634 10588 228640 10600
rect 200172 10560 228640 10588
rect 200172 10548 200178 10560
rect 228634 10548 228640 10560
rect 228692 10548 228698 10600
rect 264422 10588 264428 10600
rect 228744 10560 264428 10588
rect 91002 10480 91008 10532
rect 91060 10520 91066 10532
rect 124214 10520 124220 10532
rect 91060 10492 124220 10520
rect 91060 10480 91066 10492
rect 124214 10480 124220 10492
rect 124272 10480 124278 10532
rect 124674 10480 124680 10532
rect 124732 10520 124738 10532
rect 158806 10520 158812 10532
rect 124732 10492 158812 10520
rect 124732 10480 124738 10492
rect 158806 10480 158812 10492
rect 158864 10480 158870 10532
rect 160462 10480 160468 10532
rect 160520 10520 160526 10532
rect 182082 10520 182088 10532
rect 160520 10492 182088 10520
rect 160520 10480 160526 10492
rect 182082 10480 182088 10492
rect 182140 10480 182146 10532
rect 193306 10480 193312 10532
rect 193364 10520 193370 10532
rect 220078 10520 220084 10532
rect 193364 10492 220084 10520
rect 193364 10480 193370 10492
rect 220078 10480 220084 10492
rect 220136 10480 220142 10532
rect 223482 10480 223488 10532
rect 223540 10520 223546 10532
rect 228744 10520 228772 10560
rect 264422 10548 264428 10560
rect 264480 10548 264486 10600
rect 223540 10492 228772 10520
rect 223540 10480 223546 10492
rect 228818 10480 228824 10532
rect 228876 10520 228882 10532
rect 232774 10520 232780 10532
rect 228876 10492 232780 10520
rect 228876 10480 228882 10492
rect 232774 10480 232780 10492
rect 232832 10480 232838 10532
rect 233602 10480 233608 10532
rect 233660 10520 233666 10532
rect 257614 10520 257620 10532
rect 233660 10492 257620 10520
rect 233660 10480 233666 10492
rect 257614 10480 257620 10492
rect 257672 10480 257678 10532
rect 258626 10480 258632 10532
rect 258684 10520 258690 10532
rect 266998 10520 267004 10532
rect 258684 10492 267004 10520
rect 258684 10480 258690 10492
rect 266998 10480 267004 10492
rect 267056 10480 267062 10532
rect 62080 10424 64874 10452
rect 62080 10412 62086 10424
rect 74534 10412 74540 10464
rect 74592 10452 74598 10464
rect 96614 10452 96620 10464
rect 74592 10424 96620 10452
rect 74592 10412 74598 10424
rect 96614 10412 96620 10424
rect 96672 10412 96678 10464
rect 98822 10412 98828 10464
rect 98880 10452 98886 10464
rect 122834 10452 122840 10464
rect 98880 10424 122840 10452
rect 98880 10412 98886 10424
rect 122834 10412 122840 10424
rect 122892 10412 122898 10464
rect 145374 10412 145380 10464
rect 145432 10452 145438 10464
rect 178034 10452 178040 10464
rect 145432 10424 178040 10452
rect 145432 10412 145438 10424
rect 178034 10412 178040 10424
rect 178092 10412 178098 10464
rect 223574 10412 223580 10464
rect 223632 10452 223638 10464
rect 251266 10452 251272 10464
rect 223632 10424 251272 10452
rect 223632 10412 223638 10424
rect 251266 10412 251272 10424
rect 251324 10412 251330 10464
rect 259546 10412 259552 10464
rect 259604 10452 259610 10464
rect 269022 10452 269028 10464
rect 259604 10424 269028 10452
rect 259604 10412 259610 10424
rect 269022 10412 269028 10424
rect 269080 10412 269086 10464
rect 27764 10356 41414 10384
rect 58544 10356 64874 10384
rect 27764 10344 27770 10356
rect 58544 10328 58572 10356
rect 24486 10276 24492 10328
rect 24544 10316 24550 10328
rect 58526 10316 58532 10328
rect 24544 10288 58532 10316
rect 24544 10276 24550 10288
rect 58526 10276 58532 10288
rect 58584 10276 58590 10328
rect 63218 10316 63224 10328
rect 60706 10288 63224 10316
rect 29546 10208 29552 10260
rect 29604 10248 29610 10260
rect 60706 10248 60734 10288
rect 63218 10276 63224 10288
rect 63276 10276 63282 10328
rect 64846 10316 64874 10356
rect 80606 10344 80612 10396
rect 80664 10384 80670 10396
rect 90726 10384 90732 10396
rect 80664 10356 90732 10384
rect 80664 10344 80670 10356
rect 90726 10344 90732 10356
rect 90784 10384 90790 10396
rect 91002 10384 91008 10396
rect 90784 10356 91008 10384
rect 90784 10344 90790 10356
rect 91002 10344 91008 10356
rect 91060 10344 91066 10396
rect 93302 10344 93308 10396
rect 93360 10384 93366 10396
rect 105446 10384 105452 10396
rect 93360 10356 105452 10384
rect 93360 10344 93366 10356
rect 105446 10344 105452 10356
rect 105504 10344 105510 10396
rect 126698 10344 126704 10396
rect 126756 10384 126762 10396
rect 161106 10384 161112 10396
rect 126756 10356 161112 10384
rect 126756 10344 126762 10356
rect 161106 10344 161112 10356
rect 161164 10344 161170 10396
rect 162118 10344 162124 10396
rect 162176 10384 162182 10396
rect 216582 10384 216588 10396
rect 162176 10356 216588 10384
rect 162176 10344 162182 10356
rect 216582 10344 216588 10356
rect 216640 10344 216646 10396
rect 219066 10344 219072 10396
rect 219124 10384 219130 10396
rect 244090 10384 244096 10396
rect 219124 10356 244096 10384
rect 219124 10344 219130 10356
rect 244090 10344 244096 10356
rect 244148 10344 244154 10396
rect 260190 10344 260196 10396
rect 260248 10384 260254 10396
rect 268286 10384 268292 10396
rect 260248 10356 268292 10384
rect 260248 10344 260254 10356
rect 268286 10344 268292 10356
rect 268344 10344 268350 10396
rect 92842 10316 92848 10328
rect 64846 10288 92848 10316
rect 92842 10276 92848 10288
rect 92900 10276 92906 10328
rect 92934 10276 92940 10328
rect 92992 10316 92998 10328
rect 95510 10316 95516 10328
rect 92992 10288 95516 10316
rect 92992 10276 92998 10288
rect 95510 10276 95516 10288
rect 95568 10276 95574 10328
rect 95602 10276 95608 10328
rect 95660 10316 95666 10328
rect 107010 10316 107016 10328
rect 95660 10288 107016 10316
rect 95660 10276 95666 10288
rect 107010 10276 107016 10288
rect 107068 10276 107074 10328
rect 140222 10276 140228 10328
rect 140280 10316 140286 10328
rect 174262 10316 174268 10328
rect 140280 10288 174268 10316
rect 140280 10276 140286 10288
rect 174262 10276 174268 10288
rect 174320 10276 174326 10328
rect 196158 10276 196164 10328
rect 196216 10316 196222 10328
rect 226978 10316 226984 10328
rect 196216 10288 226984 10316
rect 196216 10276 196222 10288
rect 226978 10276 226984 10288
rect 227036 10276 227042 10328
rect 227070 10276 227076 10328
rect 227128 10316 227134 10328
rect 231854 10316 231860 10328
rect 227128 10288 231860 10316
rect 227128 10276 227134 10288
rect 231854 10276 231860 10288
rect 231912 10276 231918 10328
rect 231946 10276 231952 10328
rect 232004 10316 232010 10328
rect 239306 10316 239312 10328
rect 232004 10288 239312 10316
rect 232004 10276 232010 10288
rect 239306 10276 239312 10288
rect 239364 10276 239370 10328
rect 268102 10316 268108 10328
rect 244246 10288 268108 10316
rect 29604 10220 60734 10248
rect 63236 10248 63264 10276
rect 96522 10248 96528 10260
rect 63236 10220 96528 10248
rect 29604 10208 29610 10220
rect 96522 10208 96528 10220
rect 96580 10248 96586 10260
rect 131114 10248 131120 10260
rect 96580 10220 131120 10248
rect 96580 10208 96586 10220
rect 131114 10208 131120 10220
rect 131172 10208 131178 10260
rect 133782 10208 133788 10260
rect 133840 10248 133846 10260
rect 166718 10248 166724 10260
rect 133840 10220 166724 10248
rect 133840 10208 133846 10220
rect 166718 10208 166724 10220
rect 166776 10208 166782 10260
rect 203058 10208 203064 10260
rect 203116 10248 203122 10260
rect 235994 10248 236000 10260
rect 203116 10220 236000 10248
rect 203116 10208 203122 10220
rect 235994 10208 236000 10220
rect 236052 10248 236058 10260
rect 244246 10248 244274 10288
rect 268102 10276 268108 10288
rect 268160 10276 268166 10328
rect 236052 10220 244274 10248
rect 236052 10208 236058 10220
rect 259638 10208 259644 10260
rect 259696 10248 259702 10260
rect 267090 10248 267096 10260
rect 259696 10220 267096 10248
rect 259696 10208 259702 10220
rect 267090 10208 267096 10220
rect 267148 10208 267154 10260
rect 5902 10140 5908 10192
rect 5960 10180 5966 10192
rect 39574 10180 39580 10192
rect 5960 10152 39580 10180
rect 5960 10140 5966 10152
rect 39574 10140 39580 10152
rect 39632 10140 39638 10192
rect 56318 10140 56324 10192
rect 56376 10180 56382 10192
rect 80606 10180 80612 10192
rect 56376 10152 80612 10180
rect 56376 10140 56382 10152
rect 80606 10140 80612 10152
rect 80664 10140 80670 10192
rect 81066 10140 81072 10192
rect 81124 10180 81130 10192
rect 92934 10180 92940 10192
rect 81124 10152 92940 10180
rect 81124 10140 81130 10152
rect 92934 10140 92940 10152
rect 92992 10140 92998 10192
rect 93026 10140 93032 10192
rect 93084 10180 93090 10192
rect 126698 10180 126704 10192
rect 93084 10152 126704 10180
rect 93084 10140 93090 10152
rect 126698 10140 126704 10152
rect 126756 10140 126762 10192
rect 141418 10140 141424 10192
rect 141476 10180 141482 10192
rect 175550 10180 175556 10192
rect 141476 10152 175556 10180
rect 141476 10140 141482 10152
rect 175550 10140 175556 10152
rect 175608 10140 175614 10192
rect 197078 10140 197084 10192
rect 197136 10180 197142 10192
rect 204346 10180 204352 10192
rect 197136 10152 204352 10180
rect 197136 10140 197142 10152
rect 204346 10140 204352 10152
rect 204404 10140 204410 10192
rect 211246 10140 211252 10192
rect 211304 10180 211310 10192
rect 227070 10180 227076 10192
rect 211304 10152 227076 10180
rect 211304 10140 211310 10152
rect 227070 10140 227076 10152
rect 227128 10140 227134 10192
rect 227162 10140 227168 10192
rect 227220 10180 227226 10192
rect 227220 10152 229140 10180
rect 227220 10140 227226 10152
rect 22646 10072 22652 10124
rect 22704 10112 22710 10124
rect 56870 10112 56876 10124
rect 22704 10084 56876 10112
rect 22704 10072 22710 10084
rect 56870 10072 56876 10084
rect 56928 10072 56934 10124
rect 91002 10112 91008 10124
rect 60706 10084 91008 10112
rect 22462 10004 22468 10056
rect 22520 10044 22526 10056
rect 30558 10044 30564 10056
rect 22520 10016 30564 10044
rect 22520 10004 22526 10016
rect 30558 10004 30564 10016
rect 30616 10004 30622 10056
rect 30650 10004 30656 10056
rect 30708 10044 30714 10056
rect 56410 10044 56416 10056
rect 30708 10016 56416 10044
rect 30708 10004 30714 10016
rect 56410 10004 56416 10016
rect 56468 10044 56474 10056
rect 60706 10044 60734 10084
rect 91002 10072 91008 10084
rect 91060 10112 91066 10124
rect 124674 10112 124680 10124
rect 91060 10084 124680 10112
rect 91060 10072 91066 10084
rect 124674 10072 124680 10084
rect 124732 10072 124738 10124
rect 125870 10072 125876 10124
rect 125928 10112 125934 10124
rect 125928 10084 132494 10112
rect 125928 10072 125934 10084
rect 56468 10016 60734 10044
rect 56468 10004 56474 10016
rect 61470 10004 61476 10056
rect 61528 10044 61534 10056
rect 95418 10044 95424 10056
rect 61528 10016 95424 10044
rect 61528 10004 61534 10016
rect 95418 10004 95424 10016
rect 95476 10004 95482 10056
rect 95510 10004 95516 10056
rect 95568 10044 95574 10056
rect 95786 10044 95792 10056
rect 95568 10016 95792 10044
rect 95568 10004 95574 10016
rect 95786 10004 95792 10016
rect 95844 10044 95850 10056
rect 98546 10044 98552 10056
rect 95844 10016 98552 10044
rect 95844 10004 95850 10016
rect 98546 10004 98552 10016
rect 98604 10004 98610 10056
rect 98638 10004 98644 10056
rect 98696 10044 98702 10056
rect 130102 10044 130108 10056
rect 98696 10016 130108 10044
rect 98696 10004 98702 10016
rect 130102 10004 130108 10016
rect 130160 10004 130166 10056
rect 25498 9936 25504 9988
rect 25556 9976 25562 9988
rect 59722 9976 59728 9988
rect 25556 9948 59728 9976
rect 25556 9936 25562 9948
rect 59722 9936 59728 9948
rect 59780 9936 59786 9988
rect 81526 9936 81532 9988
rect 81584 9976 81590 9988
rect 110506 9976 110512 9988
rect 81584 9948 110512 9976
rect 81584 9936 81590 9948
rect 110506 9936 110512 9948
rect 110564 9936 110570 9988
rect 130120 9976 130148 10004
rect 132466 9976 132494 10084
rect 142430 10072 142436 10124
rect 142488 10112 142494 10124
rect 152550 10112 152556 10124
rect 142488 10084 152556 10112
rect 142488 10072 142494 10084
rect 152550 10072 152556 10084
rect 152608 10072 152614 10124
rect 159634 10072 159640 10124
rect 159692 10112 159698 10124
rect 229002 10112 229008 10124
rect 159692 10084 229008 10112
rect 159692 10072 159698 10084
rect 229002 10072 229008 10084
rect 229060 10072 229066 10124
rect 159910 10044 159916 10056
rect 137986 10016 159916 10044
rect 137986 9976 138014 10016
rect 159910 10004 159916 10016
rect 159968 10004 159974 10056
rect 165338 10044 165344 10056
rect 163792 10016 165344 10044
rect 130120 9948 130332 9976
rect 132466 9948 138014 9976
rect 18046 9868 18052 9920
rect 18104 9908 18110 9920
rect 27614 9908 27620 9920
rect 18104 9880 27620 9908
rect 18104 9868 18110 9880
rect 27614 9868 27620 9880
rect 27672 9868 27678 9920
rect 30098 9868 30104 9920
rect 30156 9908 30162 9920
rect 64046 9908 64052 9920
rect 30156 9880 64052 9908
rect 30156 9868 30162 9880
rect 64046 9868 64052 9880
rect 64104 9868 64110 9920
rect 84010 9868 84016 9920
rect 84068 9908 84074 9920
rect 117038 9908 117044 9920
rect 84068 9880 117044 9908
rect 84068 9868 84074 9880
rect 117038 9868 117044 9880
rect 117096 9868 117102 9920
rect 121638 9868 121644 9920
rect 121696 9908 121702 9920
rect 130194 9908 130200 9920
rect 121696 9880 130200 9908
rect 121696 9868 121702 9880
rect 130194 9868 130200 9880
rect 130252 9868 130258 9920
rect 130304 9908 130332 9948
rect 152458 9936 152464 9988
rect 152516 9976 152522 9988
rect 161934 9976 161940 9988
rect 152516 9948 161940 9976
rect 152516 9936 152522 9948
rect 161934 9936 161940 9948
rect 161992 9936 161998 9988
rect 158622 9908 158628 9920
rect 130304 9880 158628 9908
rect 158622 9868 158628 9880
rect 158680 9868 158686 9920
rect 158714 9868 158720 9920
rect 158772 9908 158778 9920
rect 163792 9908 163820 10016
rect 165338 10004 165344 10016
rect 165396 10004 165402 10056
rect 166166 10004 166172 10056
rect 166224 10044 166230 10056
rect 219986 10044 219992 10056
rect 166224 10016 219992 10044
rect 166224 10004 166230 10016
rect 219986 10004 219992 10016
rect 220044 10004 220050 10056
rect 220446 10004 220452 10056
rect 220504 10044 220510 10056
rect 228726 10044 228732 10056
rect 220504 10016 228732 10044
rect 220504 10004 220510 10016
rect 228726 10004 228732 10016
rect 228784 10004 228790 10056
rect 229112 10044 229140 10152
rect 231854 10140 231860 10192
rect 231912 10180 231918 10192
rect 265618 10180 265624 10192
rect 231912 10152 265624 10180
rect 231912 10140 231918 10152
rect 265618 10140 265624 10152
rect 265676 10140 265682 10192
rect 229186 10072 229192 10124
rect 229244 10112 229250 10124
rect 231946 10112 231952 10124
rect 229244 10084 231952 10112
rect 229244 10072 229250 10084
rect 231946 10072 231952 10084
rect 232004 10072 232010 10124
rect 233510 10072 233516 10124
rect 233568 10112 233574 10124
rect 258534 10112 258540 10124
rect 233568 10084 258540 10112
rect 233568 10072 233574 10084
rect 258534 10072 258540 10084
rect 258592 10072 258598 10124
rect 258902 10072 258908 10124
rect 258960 10112 258966 10124
rect 266538 10112 266544 10124
rect 258960 10084 266544 10112
rect 258960 10072 258966 10084
rect 266538 10072 266544 10084
rect 266596 10072 266602 10124
rect 261570 10044 261576 10056
rect 229112 10016 261576 10044
rect 261570 10004 261576 10016
rect 261628 10004 261634 10056
rect 262674 10004 262680 10056
rect 262732 10044 262738 10056
rect 268378 10044 268384 10056
rect 262732 10016 268384 10044
rect 262732 10004 262738 10016
rect 268378 10004 268384 10016
rect 268436 10004 268442 10056
rect 163866 9936 163872 9988
rect 163924 9976 163930 9988
rect 216582 9976 216588 9988
rect 163924 9948 216588 9976
rect 163924 9936 163930 9948
rect 216582 9936 216588 9948
rect 216640 9936 216646 9988
rect 220078 9936 220084 9988
rect 220136 9976 220142 9988
rect 227162 9976 227168 9988
rect 220136 9948 227168 9976
rect 220136 9936 220142 9948
rect 227162 9936 227168 9948
rect 227220 9936 227226 9988
rect 227806 9936 227812 9988
rect 227864 9976 227870 9988
rect 262122 9976 262128 9988
rect 227864 9948 262128 9976
rect 227864 9936 227870 9948
rect 262122 9936 262128 9948
rect 262180 9936 262186 9988
rect 264790 9936 264796 9988
rect 264848 9976 264854 9988
rect 268194 9976 268200 9988
rect 264848 9948 268200 9976
rect 264848 9936 264854 9948
rect 268194 9936 268200 9948
rect 268252 9936 268258 9988
rect 158772 9880 163820 9908
rect 158772 9868 158778 9880
rect 164234 9868 164240 9920
rect 164292 9908 164298 9920
rect 176838 9908 176844 9920
rect 164292 9880 176844 9908
rect 164292 9868 164298 9880
rect 176838 9868 176844 9880
rect 176896 9868 176902 9920
rect 196342 9868 196348 9920
rect 196400 9908 196406 9920
rect 204254 9908 204260 9920
rect 196400 9880 204260 9908
rect 196400 9868 196406 9880
rect 204254 9868 204260 9880
rect 204312 9868 204318 9920
rect 204346 9868 204352 9920
rect 204404 9908 204410 9920
rect 220170 9908 220176 9920
rect 204404 9880 220176 9908
rect 204404 9868 204410 9880
rect 220170 9868 220176 9880
rect 220228 9868 220234 9920
rect 220262 9868 220268 9920
rect 220320 9908 220326 9920
rect 229646 9908 229652 9920
rect 220320 9880 229652 9908
rect 220320 9868 220326 9880
rect 229646 9868 229652 9880
rect 229704 9908 229710 9920
rect 230934 9908 230940 9920
rect 229704 9880 230940 9908
rect 229704 9868 229710 9880
rect 230934 9868 230940 9880
rect 230992 9868 230998 9920
rect 231026 9868 231032 9920
rect 231084 9908 231090 9920
rect 236638 9908 236644 9920
rect 231084 9880 236644 9908
rect 231084 9868 231090 9880
rect 236638 9868 236644 9880
rect 236696 9868 236702 9920
rect 236730 9868 236736 9920
rect 236788 9908 236794 9920
rect 258718 9908 258724 9920
rect 236788 9880 258724 9908
rect 236788 9868 236794 9880
rect 258718 9868 258724 9880
rect 258776 9868 258782 9920
rect 258810 9868 258816 9920
rect 258868 9908 258874 9920
rect 264238 9908 264244 9920
rect 258868 9880 264244 9908
rect 258868 9868 258874 9880
rect 264238 9868 264244 9880
rect 264296 9868 264302 9920
rect 265434 9868 265440 9920
rect 265492 9908 265498 9920
rect 267734 9908 267740 9920
rect 265492 9880 267740 9908
rect 265492 9868 265498 9880
rect 267734 9868 267740 9880
rect 267792 9868 267798 9920
rect 1104 9818 271651 9840
rect 1104 9766 68546 9818
rect 68598 9766 68610 9818
rect 68662 9766 68674 9818
rect 68726 9766 68738 9818
rect 68790 9766 68802 9818
rect 68854 9766 136143 9818
rect 136195 9766 136207 9818
rect 136259 9766 136271 9818
rect 136323 9766 136335 9818
rect 136387 9766 136399 9818
rect 136451 9766 203740 9818
rect 203792 9766 203804 9818
rect 203856 9766 203868 9818
rect 203920 9766 203932 9818
rect 203984 9766 203996 9818
rect 204048 9766 271337 9818
rect 271389 9766 271401 9818
rect 271453 9766 271465 9818
rect 271517 9766 271529 9818
rect 271581 9766 271593 9818
rect 271645 9766 271651 9818
rect 1104 9744 271651 9766
rect 5902 9664 5908 9716
rect 5960 9664 5966 9716
rect 6917 9707 6975 9713
rect 6917 9673 6929 9707
rect 6963 9704 6975 9707
rect 6963 9676 25820 9704
rect 6963 9673 6975 9676
rect 6917 9667 6975 9673
rect 1670 9596 1676 9648
rect 1728 9596 1734 9648
rect 2406 9596 2412 9648
rect 2464 9596 2470 9648
rect 3234 9596 3240 9648
rect 3292 9596 3298 9648
rect 4338 9596 4344 9648
rect 4396 9596 4402 9648
rect 5074 9596 5080 9648
rect 5132 9596 5138 9648
rect 5810 9596 5816 9648
rect 5868 9596 5874 9648
rect 6822 9596 6828 9648
rect 6880 9596 6886 9648
rect 7558 9596 7564 9648
rect 7616 9596 7622 9648
rect 8386 9596 8392 9648
rect 8444 9596 8450 9648
rect 9493 9639 9551 9645
rect 9493 9605 9505 9639
rect 9539 9636 9551 9639
rect 9582 9636 9588 9648
rect 9539 9608 9588 9636
rect 9539 9605 9551 9608
rect 9493 9599 9551 9605
rect 9582 9596 9588 9608
rect 9640 9596 9646 9648
rect 10226 9596 10232 9648
rect 10284 9596 10290 9648
rect 10962 9596 10968 9648
rect 11020 9596 11026 9648
rect 11974 9596 11980 9648
rect 12032 9596 12038 9648
rect 12710 9596 12716 9648
rect 12768 9596 12774 9648
rect 13541 9639 13599 9645
rect 13541 9605 13553 9639
rect 13587 9636 13599 9639
rect 13722 9636 13728 9648
rect 13587 9608 13728 9636
rect 13587 9605 13599 9608
rect 13541 9599 13599 9605
rect 13722 9596 13728 9608
rect 13780 9596 13786 9648
rect 14642 9596 14648 9648
rect 14700 9596 14706 9648
rect 15378 9596 15384 9648
rect 15436 9596 15442 9648
rect 16114 9596 16120 9648
rect 16172 9596 16178 9648
rect 17126 9596 17132 9648
rect 17184 9596 17190 9648
rect 17862 9596 17868 9648
rect 17920 9596 17926 9648
rect 18046 9596 18052 9648
rect 18104 9596 18110 9648
rect 18598 9596 18604 9648
rect 18656 9596 18662 9648
rect 24394 9636 24400 9648
rect 22066 9608 24400 9636
rect 8573 9571 8631 9577
rect 8573 9537 8585 9571
rect 8619 9568 8631 9571
rect 22066 9568 22094 9608
rect 24394 9596 24400 9608
rect 24452 9596 24458 9648
rect 8619 9540 22094 9568
rect 8619 9537 8631 9540
rect 8573 9531 8631 9537
rect 22462 9528 22468 9580
rect 22520 9528 22526 9580
rect 22557 9571 22615 9577
rect 22557 9537 22569 9571
rect 22603 9568 22615 9571
rect 23477 9571 23535 9577
rect 23477 9568 23489 9571
rect 22603 9540 23489 9568
rect 22603 9537 22615 9540
rect 22557 9531 22615 9537
rect 23477 9537 23489 9540
rect 23523 9568 23535 9571
rect 24673 9571 24731 9577
rect 24673 9568 24685 9571
rect 23523 9540 24685 9568
rect 23523 9537 23535 9540
rect 23477 9531 23535 9537
rect 24673 9537 24685 9540
rect 24719 9568 24731 9571
rect 25682 9568 25688 9580
rect 24719 9540 25688 9568
rect 24719 9537 24731 9540
rect 24673 9531 24731 9537
rect 25682 9528 25688 9540
rect 25740 9528 25746 9580
rect 12161 9503 12219 9509
rect 12161 9469 12173 9503
rect 12207 9500 12219 9503
rect 16482 9500 16488 9512
rect 12207 9472 16488 9500
rect 12207 9469 12219 9472
rect 12161 9463 12219 9469
rect 16482 9460 16488 9472
rect 16540 9460 16546 9512
rect 17218 9460 17224 9512
rect 17276 9500 17282 9512
rect 23293 9503 23351 9509
rect 17276 9472 21404 9500
rect 17276 9460 17282 9472
rect 2593 9435 2651 9441
rect 2593 9401 2605 9435
rect 2639 9432 2651 9435
rect 7558 9432 7564 9444
rect 2639 9404 7564 9432
rect 2639 9401 2651 9404
rect 2593 9395 2651 9401
rect 7558 9392 7564 9404
rect 7616 9392 7622 9444
rect 9674 9392 9680 9444
rect 9732 9392 9738 9444
rect 12894 9392 12900 9444
rect 12952 9392 12958 9444
rect 13722 9392 13728 9444
rect 13780 9392 13786 9444
rect 15562 9392 15568 9444
rect 15620 9392 15626 9444
rect 16301 9435 16359 9441
rect 16301 9401 16313 9435
rect 16347 9432 16359 9435
rect 19150 9432 19156 9444
rect 16347 9404 19156 9432
rect 16347 9401 16359 9404
rect 16301 9395 16359 9401
rect 19150 9392 19156 9404
rect 19208 9392 19214 9444
rect 21376 9432 21404 9472
rect 23293 9469 23305 9503
rect 23339 9500 23351 9503
rect 23750 9500 23756 9512
rect 23339 9472 23756 9500
rect 23339 9469 23351 9472
rect 23293 9463 23351 9469
rect 23750 9460 23756 9472
rect 23808 9460 23814 9512
rect 24302 9460 24308 9512
rect 24360 9500 24366 9512
rect 24489 9503 24547 9509
rect 24489 9500 24501 9503
rect 24360 9472 24501 9500
rect 24360 9460 24366 9472
rect 24489 9469 24501 9472
rect 24535 9469 24547 9503
rect 25498 9500 25504 9512
rect 24489 9463 24547 9469
rect 25148 9472 25504 9500
rect 24578 9432 24584 9444
rect 21376 9404 24584 9432
rect 24578 9392 24584 9404
rect 24636 9392 24642 9444
rect 25148 9376 25176 9472
rect 25498 9460 25504 9472
rect 25556 9460 25562 9512
rect 25792 9500 25820 9676
rect 25866 9664 25872 9716
rect 25924 9704 25930 9716
rect 26513 9707 26571 9713
rect 26513 9704 26525 9707
rect 25924 9676 26525 9704
rect 25924 9664 25930 9676
rect 26513 9673 26525 9676
rect 26559 9673 26571 9707
rect 26513 9667 26571 9673
rect 27338 9664 27344 9716
rect 27396 9664 27402 9716
rect 29086 9664 29092 9716
rect 29144 9664 29150 9716
rect 30282 9664 30288 9716
rect 30340 9704 30346 9716
rect 30377 9707 30435 9713
rect 30377 9704 30389 9707
rect 30340 9676 30389 9704
rect 30340 9664 30346 9676
rect 30377 9673 30389 9676
rect 30423 9673 30435 9707
rect 30377 9667 30435 9673
rect 32490 9664 32496 9716
rect 32548 9664 32554 9716
rect 38194 9664 38200 9716
rect 38252 9704 38258 9716
rect 39301 9707 39359 9713
rect 39301 9704 39313 9707
rect 38252 9676 39313 9704
rect 38252 9664 38258 9676
rect 39301 9673 39313 9676
rect 39347 9673 39359 9707
rect 39301 9667 39359 9673
rect 39666 9664 39672 9716
rect 39724 9704 39730 9716
rect 54754 9704 54760 9716
rect 39724 9676 54760 9704
rect 39724 9664 39730 9676
rect 54754 9664 54760 9676
rect 54812 9664 54818 9716
rect 54846 9664 54852 9716
rect 54904 9704 54910 9716
rect 55677 9707 55735 9713
rect 55677 9704 55689 9707
rect 54904 9676 55689 9704
rect 54904 9664 54910 9676
rect 55677 9673 55689 9676
rect 55723 9673 55735 9707
rect 55677 9667 55735 9673
rect 56502 9664 56508 9716
rect 56560 9664 56566 9716
rect 57330 9664 57336 9716
rect 57388 9664 57394 9716
rect 57790 9664 57796 9716
rect 57848 9704 57854 9716
rect 58253 9707 58311 9713
rect 58253 9704 58265 9707
rect 57848 9676 58265 9704
rect 57848 9664 57854 9676
rect 58253 9673 58265 9676
rect 58299 9673 58311 9707
rect 58253 9667 58311 9673
rect 61746 9664 61752 9716
rect 61804 9664 61810 9716
rect 62482 9664 62488 9716
rect 62540 9664 62546 9716
rect 63402 9664 63408 9716
rect 63460 9664 63466 9716
rect 83182 9704 83188 9716
rect 78692 9676 83188 9704
rect 26142 9596 26148 9648
rect 26200 9636 26206 9648
rect 54294 9636 54300 9648
rect 26200 9608 54300 9636
rect 26200 9596 26206 9608
rect 54294 9596 54300 9608
rect 54352 9596 54358 9648
rect 54570 9596 54576 9648
rect 54628 9636 54634 9648
rect 60642 9636 60648 9648
rect 54628 9608 60648 9636
rect 54628 9596 54634 9608
rect 60642 9596 60648 9608
rect 60700 9596 60706 9648
rect 60737 9639 60795 9645
rect 60737 9605 60749 9639
rect 60783 9636 60795 9639
rect 67358 9636 67364 9648
rect 60783 9608 67364 9636
rect 60783 9605 60795 9608
rect 60737 9599 60795 9605
rect 67358 9596 67364 9608
rect 67416 9636 67422 9648
rect 76374 9636 76380 9648
rect 67416 9608 76380 9636
rect 67416 9596 67422 9608
rect 76374 9596 76380 9608
rect 76432 9596 76438 9648
rect 25869 9571 25927 9577
rect 25869 9537 25881 9571
rect 25915 9568 25927 9571
rect 26329 9571 26387 9577
rect 26329 9568 26341 9571
rect 25915 9540 26341 9568
rect 25915 9537 25927 9540
rect 25869 9531 25927 9537
rect 26329 9537 26341 9540
rect 26375 9537 26387 9571
rect 26329 9531 26387 9537
rect 26510 9528 26516 9580
rect 26568 9568 26574 9580
rect 27157 9571 27215 9577
rect 27157 9568 27169 9571
rect 26568 9540 27169 9568
rect 26568 9528 26574 9540
rect 27157 9537 27169 9540
rect 27203 9537 27215 9571
rect 27157 9531 27215 9537
rect 28905 9571 28963 9577
rect 28905 9537 28917 9571
rect 28951 9568 28963 9571
rect 29822 9568 29828 9580
rect 28951 9540 29828 9568
rect 28951 9537 28963 9540
rect 28905 9531 28963 9537
rect 29822 9528 29828 9540
rect 29880 9528 29886 9580
rect 30193 9571 30251 9577
rect 30193 9537 30205 9571
rect 30239 9568 30251 9571
rect 30374 9568 30380 9580
rect 30239 9540 30380 9568
rect 30239 9537 30251 9540
rect 30193 9531 30251 9537
rect 30374 9528 30380 9540
rect 30432 9528 30438 9580
rect 32122 9528 32128 9580
rect 32180 9568 32186 9580
rect 32309 9571 32367 9577
rect 32309 9568 32321 9571
rect 32180 9540 32321 9568
rect 32180 9528 32186 9540
rect 32309 9537 32321 9540
rect 32355 9537 32367 9571
rect 32309 9531 32367 9537
rect 35618 9528 35624 9580
rect 35676 9528 35682 9580
rect 36262 9528 36268 9580
rect 36320 9528 36326 9580
rect 36906 9528 36912 9580
rect 36964 9528 36970 9580
rect 38102 9528 38108 9580
rect 38160 9528 38166 9580
rect 38838 9528 38844 9580
rect 38896 9528 38902 9580
rect 39482 9528 39488 9580
rect 39540 9528 39546 9580
rect 40770 9528 40776 9580
rect 40828 9528 40834 9580
rect 41414 9528 41420 9580
rect 41472 9528 41478 9580
rect 42058 9528 42064 9580
rect 42116 9528 42122 9580
rect 43254 9528 43260 9580
rect 43312 9528 43318 9580
rect 43990 9528 43996 9580
rect 44048 9528 44054 9580
rect 44634 9528 44640 9580
rect 44692 9528 44698 9580
rect 45922 9528 45928 9580
rect 45980 9528 45986 9580
rect 46566 9528 46572 9580
rect 46624 9528 46630 9580
rect 47210 9528 47216 9580
rect 47268 9528 47274 9580
rect 48222 9528 48228 9580
rect 48280 9568 48286 9580
rect 48409 9571 48467 9577
rect 48409 9568 48421 9571
rect 48280 9540 48421 9568
rect 48280 9528 48286 9540
rect 48409 9537 48421 9540
rect 48455 9537 48467 9571
rect 48409 9531 48467 9537
rect 49142 9528 49148 9580
rect 49200 9528 49206 9580
rect 49786 9528 49792 9580
rect 49844 9528 49850 9580
rect 50614 9528 50620 9580
rect 50672 9528 50678 9580
rect 51350 9528 51356 9580
rect 51408 9528 51414 9580
rect 52086 9528 52092 9580
rect 52144 9528 52150 9580
rect 53098 9528 53104 9580
rect 53156 9528 53162 9580
rect 54481 9571 54539 9577
rect 54481 9537 54493 9571
rect 54527 9568 54539 9571
rect 54662 9568 54668 9580
rect 54527 9540 54668 9568
rect 54527 9537 54539 9540
rect 54481 9531 54539 9537
rect 54662 9528 54668 9540
rect 54720 9528 54726 9580
rect 54938 9528 54944 9580
rect 54996 9568 55002 9580
rect 55493 9571 55551 9577
rect 55493 9568 55505 9571
rect 54996 9540 55505 9568
rect 54996 9528 55002 9540
rect 55493 9537 55505 9540
rect 55539 9537 55551 9571
rect 55493 9531 55551 9537
rect 56321 9571 56379 9577
rect 56321 9537 56333 9571
rect 56367 9568 56379 9571
rect 56594 9568 56600 9580
rect 56367 9540 56600 9568
rect 56367 9537 56379 9540
rect 56321 9531 56379 9537
rect 56594 9528 56600 9540
rect 56652 9528 56658 9580
rect 57149 9571 57207 9577
rect 57149 9537 57161 9571
rect 57195 9568 57207 9571
rect 57330 9568 57336 9580
rect 57195 9540 57336 9568
rect 57195 9537 57207 9540
rect 57149 9531 57207 9537
rect 57330 9528 57336 9540
rect 57388 9528 57394 9580
rect 58066 9528 58072 9580
rect 58124 9528 58130 9580
rect 61565 9571 61623 9577
rect 61565 9537 61577 9571
rect 61611 9568 61623 9571
rect 62206 9568 62212 9580
rect 61611 9540 62212 9568
rect 61611 9537 61623 9540
rect 61565 9531 61623 9537
rect 62206 9528 62212 9540
rect 62264 9528 62270 9580
rect 62301 9571 62359 9577
rect 62301 9537 62313 9571
rect 62347 9568 62359 9571
rect 62574 9568 62580 9580
rect 62347 9540 62580 9568
rect 62347 9537 62359 9540
rect 62301 9531 62359 9537
rect 62574 9528 62580 9540
rect 62632 9528 62638 9580
rect 62758 9528 62764 9580
rect 62816 9568 62822 9580
rect 63221 9571 63279 9577
rect 63221 9568 63233 9571
rect 62816 9540 63233 9568
rect 62816 9528 62822 9540
rect 63221 9537 63233 9540
rect 63267 9537 63279 9571
rect 63221 9531 63279 9537
rect 69106 9528 69112 9580
rect 69164 9528 69170 9580
rect 69569 9571 69627 9577
rect 69569 9537 69581 9571
rect 69615 9568 69627 9571
rect 70302 9568 70308 9580
rect 69615 9540 70308 9568
rect 69615 9537 69627 9540
rect 69569 9531 69627 9537
rect 70302 9528 70308 9540
rect 70360 9528 70366 9580
rect 71498 9528 71504 9580
rect 71556 9528 71562 9580
rect 72142 9528 72148 9580
rect 72200 9528 72206 9580
rect 74718 9528 74724 9580
rect 74776 9528 74782 9580
rect 77294 9528 77300 9580
rect 77352 9528 77358 9580
rect 30466 9500 30472 9512
rect 25792 9472 30472 9500
rect 30466 9460 30472 9472
rect 30524 9460 30530 9512
rect 30558 9460 30564 9512
rect 30616 9500 30622 9512
rect 30616 9472 51948 9500
rect 30616 9460 30622 9472
rect 25222 9392 25228 9444
rect 25280 9432 25286 9444
rect 46198 9432 46204 9444
rect 25280 9404 46204 9432
rect 25280 9392 25286 9404
rect 46198 9392 46204 9404
rect 46256 9392 46262 9444
rect 48590 9392 48596 9444
rect 48648 9432 48654 9444
rect 49605 9435 49663 9441
rect 49605 9432 49617 9435
rect 48648 9404 49617 9432
rect 48648 9392 48654 9404
rect 49605 9401 49617 9404
rect 49651 9401 49663 9435
rect 49605 9395 49663 9401
rect 51169 9435 51227 9441
rect 51169 9401 51181 9435
rect 51215 9432 51227 9435
rect 51810 9432 51816 9444
rect 51215 9404 51816 9432
rect 51215 9401 51227 9404
rect 51169 9395 51227 9401
rect 51810 9392 51816 9404
rect 51868 9392 51874 9444
rect 51920 9432 51948 9472
rect 54294 9460 54300 9512
rect 54352 9460 54358 9512
rect 54754 9460 54760 9512
rect 54812 9500 54818 9512
rect 66070 9500 66076 9512
rect 54812 9472 66076 9500
rect 54812 9460 54818 9472
rect 66070 9460 66076 9472
rect 66128 9460 66134 9512
rect 69842 9460 69848 9512
rect 69900 9460 69906 9512
rect 72421 9503 72479 9509
rect 72421 9469 72433 9503
rect 72467 9500 72479 9503
rect 74997 9503 75055 9509
rect 72467 9472 74534 9500
rect 72467 9469 72479 9472
rect 72421 9463 72479 9469
rect 56318 9432 56324 9444
rect 51920 9404 56324 9432
rect 56318 9392 56324 9404
rect 56376 9392 56382 9444
rect 59722 9392 59728 9444
rect 59780 9432 59786 9444
rect 61289 9435 61347 9441
rect 61289 9432 61301 9435
rect 59780 9404 61301 9432
rect 59780 9392 59786 9404
rect 61289 9401 61301 9404
rect 61335 9401 61347 9435
rect 73706 9432 73712 9444
rect 61289 9395 61347 9401
rect 64846 9404 73712 9432
rect 1765 9367 1823 9373
rect 1765 9333 1777 9367
rect 1811 9364 1823 9367
rect 3234 9364 3240 9376
rect 1811 9336 3240 9364
rect 1811 9333 1823 9336
rect 1765 9327 1823 9333
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 3329 9367 3387 9373
rect 3329 9333 3341 9367
rect 3375 9364 3387 9367
rect 4062 9364 4068 9376
rect 3375 9336 4068 9364
rect 3375 9333 3387 9336
rect 3329 9327 3387 9333
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 4430 9324 4436 9376
rect 4488 9324 4494 9376
rect 5166 9324 5172 9376
rect 5224 9324 5230 9376
rect 7650 9324 7656 9376
rect 7708 9324 7714 9376
rect 10318 9324 10324 9376
rect 10376 9324 10382 9376
rect 11054 9324 11060 9376
rect 11112 9324 11118 9376
rect 14734 9324 14740 9376
rect 14792 9324 14798 9376
rect 17221 9367 17279 9373
rect 17221 9333 17233 9367
rect 17267 9364 17279 9367
rect 18598 9364 18604 9376
rect 17267 9336 18604 9364
rect 17267 9333 17279 9336
rect 17221 9327 17279 9333
rect 18598 9324 18604 9336
rect 18656 9324 18662 9376
rect 18690 9324 18696 9376
rect 18748 9324 18754 9376
rect 20254 9324 20260 9376
rect 20312 9364 20318 9376
rect 22741 9367 22799 9373
rect 22741 9364 22753 9367
rect 20312 9336 22753 9364
rect 20312 9324 20318 9336
rect 22741 9333 22753 9336
rect 22787 9333 22799 9367
rect 22741 9327 22799 9333
rect 22922 9324 22928 9376
rect 22980 9364 22986 9376
rect 23661 9367 23719 9373
rect 23661 9364 23673 9367
rect 22980 9336 23673 9364
rect 22980 9324 22986 9336
rect 23661 9333 23673 9336
rect 23707 9333 23719 9367
rect 23661 9327 23719 9333
rect 24670 9324 24676 9376
rect 24728 9364 24734 9376
rect 24857 9367 24915 9373
rect 24857 9364 24869 9367
rect 24728 9336 24869 9364
rect 24728 9324 24734 9336
rect 24857 9333 24869 9336
rect 24903 9333 24915 9367
rect 24857 9327 24915 9333
rect 25130 9324 25136 9376
rect 25188 9324 25194 9376
rect 35437 9367 35495 9373
rect 35437 9333 35449 9367
rect 35483 9364 35495 9367
rect 35618 9364 35624 9376
rect 35483 9336 35624 9364
rect 35483 9333 35495 9336
rect 35437 9327 35495 9333
rect 35618 9324 35624 9336
rect 35676 9324 35682 9376
rect 35802 9324 35808 9376
rect 35860 9364 35866 9376
rect 36081 9367 36139 9373
rect 36081 9364 36093 9367
rect 35860 9336 36093 9364
rect 35860 9324 35866 9336
rect 36081 9333 36093 9336
rect 36127 9333 36139 9367
rect 36081 9327 36139 9333
rect 36630 9324 36636 9376
rect 36688 9364 36694 9376
rect 36725 9367 36783 9373
rect 36725 9364 36737 9367
rect 36688 9336 36737 9364
rect 36688 9324 36694 9336
rect 36725 9333 36737 9336
rect 36771 9333 36783 9367
rect 36725 9327 36783 9333
rect 37918 9324 37924 9376
rect 37976 9324 37982 9376
rect 38654 9324 38660 9376
rect 38712 9324 38718 9376
rect 40494 9324 40500 9376
rect 40552 9364 40558 9376
rect 40589 9367 40647 9373
rect 40589 9364 40601 9367
rect 40552 9336 40601 9364
rect 40552 9324 40558 9336
rect 40589 9333 40601 9336
rect 40635 9333 40647 9367
rect 40589 9327 40647 9333
rect 41046 9324 41052 9376
rect 41104 9364 41110 9376
rect 41233 9367 41291 9373
rect 41233 9364 41245 9367
rect 41104 9336 41245 9364
rect 41104 9324 41110 9336
rect 41233 9333 41245 9336
rect 41279 9333 41291 9367
rect 41233 9327 41291 9333
rect 41782 9324 41788 9376
rect 41840 9364 41846 9376
rect 41877 9367 41935 9373
rect 41877 9364 41889 9367
rect 41840 9336 41889 9364
rect 41840 9324 41846 9336
rect 41877 9333 41889 9336
rect 41923 9333 41935 9367
rect 41877 9327 41935 9333
rect 42886 9324 42892 9376
rect 42944 9364 42950 9376
rect 43073 9367 43131 9373
rect 43073 9364 43085 9367
rect 42944 9336 43085 9364
rect 42944 9324 42950 9336
rect 43073 9333 43085 9336
rect 43119 9333 43131 9367
rect 43073 9327 43131 9333
rect 43254 9324 43260 9376
rect 43312 9364 43318 9376
rect 43809 9367 43867 9373
rect 43809 9364 43821 9367
rect 43312 9336 43821 9364
rect 43312 9324 43318 9336
rect 43809 9333 43821 9336
rect 43855 9333 43867 9367
rect 43809 9327 43867 9333
rect 43898 9324 43904 9376
rect 43956 9364 43962 9376
rect 44453 9367 44511 9373
rect 44453 9364 44465 9367
rect 43956 9336 44465 9364
rect 43956 9324 43962 9336
rect 44453 9333 44465 9336
rect 44499 9333 44511 9367
rect 44453 9327 44511 9333
rect 45646 9324 45652 9376
rect 45704 9364 45710 9376
rect 45741 9367 45799 9373
rect 45741 9364 45753 9367
rect 45704 9336 45753 9364
rect 45704 9324 45710 9336
rect 45741 9333 45753 9336
rect 45787 9333 45799 9367
rect 45741 9327 45799 9333
rect 46014 9324 46020 9376
rect 46072 9364 46078 9376
rect 46385 9367 46443 9373
rect 46385 9364 46397 9367
rect 46072 9336 46397 9364
rect 46072 9324 46078 9336
rect 46385 9333 46397 9336
rect 46431 9333 46443 9367
rect 46385 9327 46443 9333
rect 47026 9324 47032 9376
rect 47084 9324 47090 9376
rect 48222 9324 48228 9376
rect 48280 9324 48286 9376
rect 48406 9324 48412 9376
rect 48464 9364 48470 9376
rect 48961 9367 49019 9373
rect 48961 9364 48973 9367
rect 48464 9336 48973 9364
rect 48464 9324 48470 9336
rect 48961 9333 48973 9336
rect 49007 9333 49019 9367
rect 48961 9327 49019 9333
rect 50430 9324 50436 9376
rect 50488 9324 50494 9376
rect 51258 9324 51264 9376
rect 51316 9364 51322 9376
rect 51905 9367 51963 9373
rect 51905 9364 51917 9367
rect 51316 9336 51917 9364
rect 51316 9324 51322 9336
rect 51905 9333 51917 9336
rect 51951 9333 51963 9367
rect 51905 9327 51963 9333
rect 52270 9324 52276 9376
rect 52328 9364 52334 9376
rect 52917 9367 52975 9373
rect 52917 9364 52929 9367
rect 52328 9336 52929 9364
rect 52328 9324 52334 9336
rect 52917 9333 52929 9336
rect 52963 9333 52975 9367
rect 52917 9327 52975 9333
rect 53098 9324 53104 9376
rect 53156 9364 53162 9376
rect 54665 9367 54723 9373
rect 54665 9364 54677 9367
rect 53156 9336 54677 9364
rect 53156 9324 53162 9336
rect 54665 9333 54677 9336
rect 54711 9333 54723 9367
rect 54665 9327 54723 9333
rect 59906 9324 59912 9376
rect 59964 9364 59970 9376
rect 60829 9367 60887 9373
rect 60829 9364 60841 9367
rect 59964 9336 60841 9364
rect 59964 9324 59970 9336
rect 60829 9333 60841 9336
rect 60875 9333 60887 9367
rect 61304 9364 61332 9395
rect 64846 9364 64874 9404
rect 73706 9392 73712 9404
rect 73764 9392 73770 9444
rect 74506 9432 74534 9472
rect 74997 9469 75009 9503
rect 75043 9500 75055 9503
rect 75822 9500 75828 9512
rect 75043 9472 75828 9500
rect 75043 9469 75055 9472
rect 74997 9463 75055 9469
rect 75822 9460 75828 9472
rect 75880 9460 75886 9512
rect 77570 9460 77576 9512
rect 77628 9460 77634 9512
rect 78692 9432 78720 9676
rect 83182 9664 83188 9676
rect 83240 9664 83246 9716
rect 84010 9664 84016 9716
rect 84068 9664 84074 9716
rect 87003 9707 87061 9713
rect 87003 9673 87015 9707
rect 87049 9704 87061 9707
rect 87049 9676 92704 9704
rect 87049 9673 87061 9676
rect 87003 9667 87061 9673
rect 79226 9596 79232 9648
rect 79284 9596 79290 9648
rect 79413 9639 79471 9645
rect 79413 9605 79425 9639
rect 79459 9636 79471 9639
rect 79459 9608 83044 9636
rect 79459 9605 79471 9608
rect 79413 9599 79471 9605
rect 79873 9571 79931 9577
rect 79873 9537 79885 9571
rect 79919 9568 79931 9571
rect 79962 9568 79968 9580
rect 79919 9540 79968 9568
rect 79919 9537 79931 9540
rect 79873 9531 79931 9537
rect 79962 9528 79968 9540
rect 80020 9528 80026 9580
rect 81618 9528 81624 9580
rect 81676 9528 81682 9580
rect 83016 9568 83044 9608
rect 83090 9596 83096 9648
rect 83148 9596 83154 9648
rect 83918 9596 83924 9648
rect 83976 9596 83982 9648
rect 84654 9596 84660 9648
rect 84712 9596 84718 9648
rect 85390 9596 85396 9648
rect 85448 9596 85454 9648
rect 92676 9636 92704 9676
rect 92750 9664 92756 9716
rect 92808 9664 92814 9716
rect 93486 9664 93492 9716
rect 93544 9664 93550 9716
rect 94590 9664 94596 9716
rect 94648 9704 94654 9716
rect 95970 9704 95976 9716
rect 94648 9676 95976 9704
rect 94648 9664 94654 9676
rect 95970 9664 95976 9676
rect 96028 9664 96034 9716
rect 96062 9664 96068 9716
rect 96120 9664 96126 9716
rect 96338 9664 96344 9716
rect 96396 9704 96402 9716
rect 96893 9707 96951 9713
rect 96893 9704 96905 9707
rect 96396 9676 96905 9704
rect 96396 9664 96402 9676
rect 96893 9673 96905 9676
rect 96939 9673 96951 9707
rect 96893 9667 96951 9673
rect 99374 9664 99380 9716
rect 99432 9704 99438 9716
rect 99469 9707 99527 9713
rect 99469 9704 99481 9707
rect 99432 9676 99481 9704
rect 99432 9664 99438 9676
rect 99469 9673 99481 9676
rect 99515 9673 99527 9707
rect 99469 9667 99527 9673
rect 100478 9664 100484 9716
rect 100536 9664 100542 9716
rect 100662 9664 100668 9716
rect 100720 9704 100726 9716
rect 104713 9707 104771 9713
rect 104713 9704 104725 9707
rect 100720 9676 104725 9704
rect 100720 9664 100726 9676
rect 104713 9673 104725 9676
rect 104759 9673 104771 9707
rect 104713 9667 104771 9673
rect 105446 9664 105452 9716
rect 105504 9664 105510 9716
rect 106182 9664 106188 9716
rect 106240 9664 106246 9716
rect 107565 9707 107623 9713
rect 107565 9673 107577 9707
rect 107611 9673 107623 9707
rect 107565 9667 107623 9673
rect 85500 9608 91876 9636
rect 92676 9608 99512 9636
rect 85500 9568 85528 9608
rect 83016 9540 85528 9568
rect 86770 9528 86776 9580
rect 86828 9528 86834 9580
rect 89349 9571 89407 9577
rect 86926 9540 89300 9568
rect 80146 9460 80152 9512
rect 80204 9460 80210 9512
rect 81897 9503 81955 9509
rect 81897 9469 81909 9503
rect 81943 9500 81955 9503
rect 86926 9500 86954 9540
rect 81943 9472 86954 9500
rect 81943 9469 81955 9472
rect 81897 9463 81955 9469
rect 88978 9460 88984 9512
rect 89036 9500 89042 9512
rect 89165 9503 89223 9509
rect 89165 9500 89177 9503
rect 89036 9472 89177 9500
rect 89036 9460 89042 9472
rect 89165 9469 89177 9472
rect 89211 9469 89223 9503
rect 89272 9500 89300 9540
rect 89349 9537 89361 9571
rect 89395 9568 89407 9571
rect 89438 9568 89444 9580
rect 89395 9540 89444 9568
rect 89395 9537 89407 9540
rect 89349 9531 89407 9537
rect 89438 9528 89444 9540
rect 89496 9528 89502 9580
rect 90082 9528 90088 9580
rect 90140 9568 90146 9580
rect 90177 9571 90235 9577
rect 90177 9568 90189 9571
rect 90140 9540 90189 9568
rect 90140 9528 90146 9540
rect 90177 9537 90189 9540
rect 90223 9537 90235 9571
rect 90177 9531 90235 9537
rect 91554 9528 91560 9580
rect 91612 9528 91618 9580
rect 91646 9528 91652 9580
rect 91704 9568 91710 9580
rect 91704 9540 91784 9568
rect 91704 9528 91710 9540
rect 89272 9472 89668 9500
rect 89165 9463 89223 9469
rect 74506 9404 78720 9432
rect 79244 9404 80054 9432
rect 61304 9336 64874 9364
rect 71317 9367 71375 9373
rect 60829 9327 60887 9333
rect 71317 9333 71329 9367
rect 71363 9364 71375 9367
rect 79244 9364 79272 9404
rect 71363 9336 79272 9364
rect 80026 9364 80054 9404
rect 83274 9392 83280 9444
rect 83332 9392 83338 9444
rect 84841 9435 84899 9441
rect 84841 9401 84853 9435
rect 84887 9432 84899 9435
rect 85482 9432 85488 9444
rect 84887 9404 85488 9432
rect 84887 9401 84899 9404
rect 84841 9395 84899 9401
rect 85482 9392 85488 9404
rect 85540 9392 85546 9444
rect 85577 9435 85635 9441
rect 85577 9401 85589 9435
rect 85623 9432 85635 9435
rect 89346 9432 89352 9444
rect 85623 9404 89352 9432
rect 85623 9401 85635 9404
rect 85577 9395 85635 9401
rect 89346 9392 89352 9404
rect 89404 9392 89410 9444
rect 89533 9435 89591 9441
rect 89533 9432 89545 9435
rect 89456 9404 89545 9432
rect 88334 9364 88340 9376
rect 80026 9336 88340 9364
rect 71363 9333 71375 9336
rect 71317 9327 71375 9333
rect 88334 9324 88340 9336
rect 88392 9324 88398 9376
rect 88794 9324 88800 9376
rect 88852 9364 88858 9376
rect 89456 9364 89484 9404
rect 89533 9401 89545 9404
rect 89579 9401 89591 9435
rect 89533 9395 89591 9401
rect 88852 9336 89484 9364
rect 89640 9364 89668 9472
rect 90358 9392 90364 9444
rect 90416 9392 90422 9444
rect 91756 9441 91784 9540
rect 91848 9500 91876 9608
rect 92566 9528 92572 9580
rect 92624 9528 92630 9580
rect 93305 9571 93363 9577
rect 93305 9537 93317 9571
rect 93351 9568 93363 9571
rect 93670 9568 93676 9580
rect 93351 9540 93676 9568
rect 93351 9537 93363 9540
rect 93305 9531 93363 9537
rect 93670 9528 93676 9540
rect 93728 9528 93734 9580
rect 94774 9528 94780 9580
rect 94832 9528 94838 9580
rect 94866 9528 94872 9580
rect 94924 9568 94930 9580
rect 94961 9571 95019 9577
rect 94961 9568 94973 9571
rect 94924 9540 94973 9568
rect 94924 9528 94930 9540
rect 94961 9537 94973 9540
rect 95007 9537 95019 9571
rect 94961 9531 95019 9537
rect 95881 9571 95939 9577
rect 95881 9537 95893 9571
rect 95927 9568 95939 9571
rect 96154 9568 96160 9580
rect 95927 9540 96160 9568
rect 95927 9537 95939 9540
rect 95881 9531 95939 9537
rect 96154 9528 96160 9540
rect 96212 9528 96218 9580
rect 96709 9571 96767 9577
rect 96709 9537 96721 9571
rect 96755 9568 96767 9571
rect 96890 9568 96896 9580
rect 96755 9540 96896 9568
rect 96755 9537 96767 9540
rect 96709 9531 96767 9537
rect 96890 9528 96896 9540
rect 96948 9528 96954 9580
rect 98914 9528 98920 9580
rect 98972 9568 98978 9580
rect 99285 9571 99343 9577
rect 99285 9568 99297 9571
rect 98972 9540 99297 9568
rect 98972 9528 98978 9540
rect 99285 9537 99297 9540
rect 99331 9537 99343 9571
rect 99484 9568 99512 9608
rect 103054 9596 103060 9648
rect 103112 9636 103118 9648
rect 107580 9636 107608 9667
rect 108114 9664 108120 9716
rect 108172 9704 108178 9716
rect 108172 9676 113772 9704
rect 108172 9664 108178 9676
rect 103112 9608 107608 9636
rect 113744 9636 113772 9676
rect 113818 9664 113824 9716
rect 113876 9704 113882 9716
rect 121638 9704 121644 9716
rect 113876 9676 121644 9704
rect 113876 9664 113882 9676
rect 121638 9664 121644 9676
rect 121696 9664 121702 9716
rect 121730 9664 121736 9716
rect 121788 9664 121794 9716
rect 125226 9664 125232 9716
rect 125284 9664 125290 9716
rect 126330 9664 126336 9716
rect 126388 9664 126394 9716
rect 129553 9707 129611 9713
rect 129553 9673 129565 9707
rect 129599 9704 129611 9707
rect 129642 9704 129648 9716
rect 129599 9676 129648 9704
rect 129599 9673 129611 9676
rect 129553 9667 129611 9673
rect 129642 9664 129648 9676
rect 129700 9664 129706 9716
rect 130746 9664 130752 9716
rect 130804 9664 130810 9716
rect 131482 9664 131488 9716
rect 131540 9664 131546 9716
rect 133414 9664 133420 9716
rect 133472 9664 133478 9716
rect 134150 9664 134156 9716
rect 134208 9664 134214 9716
rect 158714 9704 158720 9716
rect 137986 9676 158720 9704
rect 117314 9636 117320 9648
rect 113744 9608 117320 9636
rect 103112 9596 103118 9608
rect 117314 9596 117320 9608
rect 117372 9596 117378 9648
rect 123294 9596 123300 9648
rect 123352 9636 123358 9648
rect 131114 9636 131120 9648
rect 123352 9608 131120 9636
rect 123352 9596 123358 9608
rect 131114 9596 131120 9608
rect 131172 9636 131178 9648
rect 137986 9636 138014 9676
rect 158714 9664 158720 9676
rect 158772 9664 158778 9716
rect 164326 9704 164332 9716
rect 158916 9676 164332 9704
rect 131172 9608 138014 9636
rect 131172 9596 131178 9608
rect 147858 9596 147864 9648
rect 147916 9636 147922 9648
rect 155678 9636 155684 9648
rect 147916 9608 155684 9636
rect 147916 9596 147922 9608
rect 155678 9596 155684 9608
rect 155736 9596 155742 9648
rect 158916 9636 158944 9676
rect 164326 9664 164332 9676
rect 164384 9664 164390 9716
rect 166644 9676 167500 9704
rect 155880 9608 158944 9636
rect 159008 9608 161336 9636
rect 100202 9568 100208 9580
rect 99484 9540 100208 9568
rect 99285 9531 99343 9537
rect 100202 9528 100208 9540
rect 100260 9528 100266 9580
rect 100297 9571 100355 9577
rect 100297 9537 100309 9571
rect 100343 9568 100355 9571
rect 100570 9568 100576 9580
rect 100343 9540 100576 9568
rect 100343 9537 100355 9540
rect 100297 9531 100355 9537
rect 100570 9528 100576 9540
rect 100628 9528 100634 9580
rect 100846 9528 100852 9580
rect 100904 9568 100910 9580
rect 100904 9540 101628 9568
rect 100904 9528 100910 9540
rect 101490 9500 101496 9512
rect 91848 9472 101496 9500
rect 101490 9460 101496 9472
rect 101548 9460 101554 9512
rect 101600 9500 101628 9540
rect 103238 9528 103244 9580
rect 103296 9528 103302 9580
rect 103882 9528 103888 9580
rect 103940 9528 103946 9580
rect 104710 9528 104716 9580
rect 104768 9568 104774 9580
rect 104897 9571 104955 9577
rect 104897 9568 104909 9571
rect 104768 9540 104909 9568
rect 104768 9528 104774 9540
rect 104897 9537 104909 9540
rect 104943 9537 104955 9571
rect 104897 9531 104955 9537
rect 105630 9528 105636 9580
rect 105688 9528 105694 9580
rect 106274 9528 106280 9580
rect 106332 9568 106338 9580
rect 106369 9571 106427 9577
rect 106369 9568 106381 9571
rect 106332 9540 106381 9568
rect 106332 9528 106338 9540
rect 106369 9537 106381 9540
rect 106415 9537 106427 9571
rect 106369 9531 106427 9537
rect 107746 9528 107752 9580
rect 107804 9528 107810 9580
rect 108390 9528 108396 9580
rect 108448 9528 108454 9580
rect 109034 9528 109040 9580
rect 109092 9528 109098 9580
rect 110046 9528 110052 9580
rect 110104 9528 110110 9580
rect 110782 9528 110788 9580
rect 110840 9528 110846 9580
rect 111518 9528 111524 9580
rect 111576 9528 111582 9580
rect 112898 9528 112904 9580
rect 112956 9528 112962 9580
rect 113542 9528 113548 9580
rect 113600 9528 113606 9580
rect 114186 9528 114192 9580
rect 114244 9528 114250 9580
rect 115198 9528 115204 9580
rect 115256 9528 115262 9580
rect 115750 9528 115756 9580
rect 115808 9568 115814 9580
rect 115937 9571 115995 9577
rect 115937 9568 115949 9571
rect 115808 9540 115949 9568
rect 115808 9528 115814 9540
rect 115937 9537 115949 9540
rect 115983 9537 115995 9571
rect 115937 9531 115995 9537
rect 116670 9528 116676 9580
rect 116728 9528 116734 9580
rect 118050 9528 118056 9580
rect 118108 9528 118114 9580
rect 118694 9528 118700 9580
rect 118752 9528 118758 9580
rect 119338 9528 119344 9580
rect 119396 9528 119402 9580
rect 120350 9528 120356 9580
rect 120408 9528 120414 9580
rect 121086 9528 121092 9580
rect 121144 9528 121150 9580
rect 121549 9571 121607 9577
rect 121549 9537 121561 9571
rect 121595 9568 121607 9571
rect 121638 9568 121644 9580
rect 121595 9540 121644 9568
rect 121595 9537 121607 9540
rect 121549 9531 121607 9537
rect 121638 9528 121644 9540
rect 121696 9528 121702 9580
rect 124398 9528 124404 9580
rect 124456 9568 124462 9580
rect 125045 9571 125103 9577
rect 125045 9568 125057 9571
rect 124456 9540 125057 9568
rect 124456 9528 124462 9540
rect 125045 9537 125057 9540
rect 125091 9537 125103 9571
rect 125045 9531 125103 9537
rect 126149 9571 126207 9577
rect 126149 9537 126161 9571
rect 126195 9568 126207 9571
rect 126238 9568 126244 9580
rect 126195 9540 126244 9568
rect 126195 9537 126207 9540
rect 126149 9531 126207 9537
rect 126238 9528 126244 9540
rect 126296 9528 126302 9580
rect 128449 9571 128507 9577
rect 128449 9537 128461 9571
rect 128495 9568 128507 9571
rect 128814 9568 128820 9580
rect 128495 9540 128820 9568
rect 128495 9537 128507 9540
rect 128449 9531 128507 9537
rect 128814 9528 128820 9540
rect 128872 9528 128878 9580
rect 129366 9528 129372 9580
rect 129424 9528 129430 9580
rect 130562 9528 130568 9580
rect 130620 9528 130626 9580
rect 131301 9571 131359 9577
rect 131301 9537 131313 9571
rect 131347 9568 131359 9571
rect 131390 9568 131396 9580
rect 131347 9540 131396 9568
rect 131347 9537 131359 9540
rect 131301 9531 131359 9537
rect 131390 9528 131396 9540
rect 131448 9528 131454 9580
rect 133046 9528 133052 9580
rect 133104 9568 133110 9580
rect 133233 9571 133291 9577
rect 133233 9568 133245 9571
rect 133104 9540 133245 9568
rect 133104 9528 133110 9540
rect 133233 9537 133245 9540
rect 133279 9537 133291 9571
rect 133233 9531 133291 9537
rect 133969 9571 134027 9577
rect 133969 9537 133981 9571
rect 134015 9568 134027 9571
rect 134058 9568 134064 9580
rect 134015 9540 134064 9568
rect 134015 9537 134027 9540
rect 133969 9531 134027 9537
rect 134058 9528 134064 9540
rect 134116 9528 134122 9580
rect 138014 9528 138020 9580
rect 138072 9568 138078 9580
rect 138109 9571 138167 9577
rect 138109 9568 138121 9571
rect 138072 9540 138121 9568
rect 138072 9528 138078 9540
rect 138109 9537 138121 9540
rect 138155 9537 138167 9571
rect 138109 9531 138167 9537
rect 138750 9528 138756 9580
rect 138808 9528 138814 9580
rect 139394 9528 139400 9580
rect 139452 9528 139458 9580
rect 140682 9528 140688 9580
rect 140740 9528 140746 9580
rect 141326 9528 141332 9580
rect 141384 9528 141390 9580
rect 141970 9528 141976 9580
rect 142028 9528 142034 9580
rect 143258 9528 143264 9580
rect 143316 9528 143322 9580
rect 143534 9528 143540 9580
rect 143592 9568 143598 9580
rect 143905 9571 143963 9577
rect 143905 9568 143917 9571
rect 143592 9540 143917 9568
rect 143592 9528 143598 9540
rect 143905 9537 143917 9540
rect 143951 9537 143963 9571
rect 143905 9531 143963 9537
rect 144546 9528 144552 9580
rect 144604 9528 144610 9580
rect 145834 9528 145840 9580
rect 145892 9528 145898 9580
rect 146294 9528 146300 9580
rect 146352 9568 146358 9580
rect 146481 9571 146539 9577
rect 146481 9568 146493 9571
rect 146352 9540 146493 9568
rect 146352 9528 146358 9540
rect 146481 9537 146493 9540
rect 146527 9537 146539 9571
rect 146481 9531 146539 9537
rect 147122 9528 147128 9580
rect 147180 9528 147186 9580
rect 148410 9528 148416 9580
rect 148468 9528 148474 9580
rect 149054 9528 149060 9580
rect 149112 9528 149118 9580
rect 149698 9528 149704 9580
rect 149756 9528 149762 9580
rect 150986 9528 150992 9580
rect 151044 9528 151050 9580
rect 151630 9528 151636 9580
rect 151688 9528 151694 9580
rect 152274 9528 152280 9580
rect 152332 9528 152338 9580
rect 152826 9528 152832 9580
rect 152884 9568 152890 9580
rect 153565 9571 153623 9577
rect 153565 9568 153577 9571
rect 152884 9540 153577 9568
rect 152884 9528 152890 9540
rect 153565 9537 153577 9540
rect 153611 9537 153623 9571
rect 153565 9531 153623 9537
rect 154206 9528 154212 9580
rect 154264 9528 154270 9580
rect 154298 9528 154304 9580
rect 154356 9568 154362 9580
rect 154853 9571 154911 9577
rect 154853 9568 154865 9571
rect 154356 9540 154865 9568
rect 154356 9528 154362 9540
rect 154853 9537 154865 9540
rect 154899 9537 154911 9571
rect 154853 9531 154911 9537
rect 127897 9503 127955 9509
rect 127897 9500 127909 9503
rect 101600 9472 108896 9500
rect 91741 9435 91799 9441
rect 91741 9401 91753 9435
rect 91787 9401 91799 9435
rect 91741 9395 91799 9401
rect 92014 9392 92020 9444
rect 92072 9432 92078 9444
rect 108114 9432 108120 9444
rect 92072 9404 108120 9432
rect 92072 9392 92078 9404
rect 108114 9392 108120 9404
rect 108172 9392 108178 9444
rect 108868 9441 108896 9472
rect 109052 9472 127909 9500
rect 109052 9444 109080 9472
rect 127897 9469 127909 9472
rect 127943 9500 127955 9503
rect 127986 9500 127992 9512
rect 127943 9472 127992 9500
rect 127943 9469 127955 9472
rect 127897 9463 127955 9469
rect 127986 9460 127992 9472
rect 128044 9500 128050 9512
rect 128265 9503 128323 9509
rect 128265 9500 128277 9503
rect 128044 9472 128277 9500
rect 128044 9460 128050 9472
rect 128265 9469 128277 9472
rect 128311 9500 128323 9503
rect 152458 9500 152464 9512
rect 128311 9472 152464 9500
rect 128311 9469 128323 9472
rect 128265 9463 128323 9469
rect 152458 9460 152464 9472
rect 152516 9460 152522 9512
rect 155880 9500 155908 9608
rect 156509 9571 156567 9577
rect 156509 9537 156521 9571
rect 156555 9568 156567 9571
rect 157334 9568 157340 9580
rect 156555 9540 157340 9568
rect 156555 9537 156567 9540
rect 156509 9531 156567 9537
rect 157334 9528 157340 9540
rect 157392 9528 157398 9580
rect 157429 9571 157487 9577
rect 157429 9537 157441 9571
rect 157475 9568 157487 9571
rect 157518 9568 157524 9580
rect 157475 9540 157524 9568
rect 157475 9537 157487 9540
rect 157429 9531 157487 9537
rect 157518 9528 157524 9540
rect 157576 9568 157582 9580
rect 159008 9577 159036 9608
rect 161308 9580 161336 9608
rect 158993 9571 159051 9577
rect 158993 9568 159005 9571
rect 157576 9540 159005 9568
rect 157576 9528 157582 9540
rect 158993 9537 159005 9540
rect 159039 9537 159051 9571
rect 158993 9531 159051 9537
rect 159729 9571 159787 9577
rect 159729 9537 159741 9571
rect 159775 9568 159787 9571
rect 161198 9568 161204 9580
rect 159775 9540 161204 9568
rect 159775 9537 159787 9540
rect 159729 9531 159787 9537
rect 161198 9528 161204 9540
rect 161256 9528 161262 9580
rect 161290 9528 161296 9580
rect 161348 9568 161354 9580
rect 162121 9571 162179 9577
rect 162121 9568 162133 9571
rect 161348 9540 162133 9568
rect 161348 9528 161354 9540
rect 162121 9537 162133 9540
rect 162167 9537 162179 9571
rect 162121 9531 162179 9537
rect 162762 9528 162768 9580
rect 162820 9528 162826 9580
rect 162949 9571 163007 9577
rect 162949 9537 162961 9571
rect 162995 9568 163007 9571
rect 163869 9571 163927 9577
rect 163869 9568 163881 9571
rect 162995 9540 163881 9568
rect 162995 9537 163007 9540
rect 162949 9531 163007 9537
rect 163869 9537 163881 9540
rect 163915 9568 163927 9571
rect 164697 9571 164755 9577
rect 164697 9568 164709 9571
rect 163915 9540 164709 9568
rect 163915 9537 163927 9540
rect 163869 9531 163927 9537
rect 164697 9537 164709 9540
rect 164743 9568 164755 9571
rect 165525 9571 165583 9577
rect 165525 9568 165537 9571
rect 164743 9540 165537 9568
rect 164743 9537 164755 9540
rect 164697 9531 164755 9537
rect 165525 9537 165537 9540
rect 165571 9568 165583 9571
rect 166534 9568 166540 9580
rect 165571 9540 166540 9568
rect 165571 9537 165583 9540
rect 165525 9531 165583 9537
rect 166534 9528 166540 9540
rect 166592 9568 166598 9580
rect 166644 9577 166672 9676
rect 166629 9571 166687 9577
rect 166629 9568 166641 9571
rect 166592 9540 166641 9568
rect 166592 9528 166598 9540
rect 166629 9537 166641 9540
rect 166675 9537 166687 9571
rect 166629 9531 166687 9537
rect 166718 9528 166724 9580
rect 166776 9568 166782 9580
rect 166902 9568 166908 9580
rect 166776 9540 166908 9568
rect 166776 9528 166782 9540
rect 166902 9528 166908 9540
rect 166960 9568 166966 9580
rect 167472 9577 167500 9676
rect 168374 9664 168380 9716
rect 168432 9704 168438 9716
rect 169021 9707 169079 9713
rect 169021 9704 169033 9707
rect 168432 9676 169033 9704
rect 168432 9664 168438 9676
rect 169021 9673 169033 9676
rect 169067 9673 169079 9707
rect 215202 9704 215208 9716
rect 169021 9667 169079 9673
rect 169772 9676 215208 9704
rect 168742 9596 168748 9648
rect 168800 9636 168806 9648
rect 169772 9636 169800 9676
rect 215202 9664 215208 9676
rect 215260 9664 215266 9716
rect 215849 9707 215907 9713
rect 215849 9673 215861 9707
rect 215895 9704 215907 9707
rect 218514 9704 218520 9716
rect 215895 9676 218520 9704
rect 215895 9673 215907 9676
rect 215849 9667 215907 9673
rect 218514 9664 218520 9676
rect 218572 9664 218578 9716
rect 220078 9664 220084 9716
rect 220136 9704 220142 9716
rect 224770 9704 224776 9716
rect 220136 9676 224776 9704
rect 220136 9664 220142 9676
rect 224770 9664 224776 9676
rect 224828 9664 224834 9716
rect 225046 9664 225052 9716
rect 225104 9704 225110 9716
rect 258810 9704 258816 9716
rect 225104 9676 258816 9704
rect 225104 9664 225110 9676
rect 258810 9664 258816 9676
rect 258868 9664 258874 9716
rect 259178 9664 259184 9716
rect 259236 9664 259242 9716
rect 260009 9707 260067 9713
rect 260009 9673 260021 9707
rect 260055 9673 260067 9707
rect 260009 9667 260067 9673
rect 168800 9608 169800 9636
rect 168800 9596 168806 9608
rect 171226 9596 171232 9648
rect 171284 9636 171290 9648
rect 171284 9608 174124 9636
rect 171284 9596 171290 9608
rect 167273 9571 167331 9577
rect 167273 9568 167285 9571
rect 166960 9540 167285 9568
rect 166960 9528 166966 9540
rect 167273 9537 167285 9540
rect 167319 9537 167331 9571
rect 167273 9531 167331 9537
rect 167457 9571 167515 9577
rect 167457 9537 167469 9571
rect 167503 9537 167515 9571
rect 167457 9531 167515 9537
rect 167641 9571 167699 9577
rect 167641 9537 167653 9571
rect 167687 9568 167699 9571
rect 168837 9571 168895 9577
rect 168837 9568 168849 9571
rect 167687 9540 168849 9568
rect 167687 9537 167699 9540
rect 167641 9531 167699 9537
rect 168837 9537 168849 9540
rect 168883 9537 168895 9571
rect 168837 9531 168895 9537
rect 169202 9528 169208 9580
rect 169260 9568 169266 9580
rect 169573 9571 169631 9577
rect 169573 9568 169585 9571
rect 169260 9540 169585 9568
rect 169260 9528 169266 9540
rect 169573 9537 169585 9540
rect 169619 9537 169631 9571
rect 169573 9531 169631 9537
rect 171686 9528 171692 9580
rect 171744 9528 171750 9580
rect 172238 9528 172244 9580
rect 172296 9528 172302 9580
rect 173986 9528 173992 9580
rect 174044 9528 174050 9580
rect 174096 9568 174124 9608
rect 174446 9596 174452 9648
rect 174504 9636 174510 9648
rect 175369 9639 175427 9645
rect 175369 9636 175381 9639
rect 174504 9608 175381 9636
rect 174504 9596 174510 9608
rect 175369 9605 175381 9608
rect 175415 9605 175427 9639
rect 175369 9599 175427 9605
rect 175550 9596 175556 9648
rect 175608 9596 175614 9648
rect 220170 9636 220176 9648
rect 175660 9608 220176 9636
rect 175660 9568 175688 9608
rect 220170 9596 220176 9608
rect 220228 9596 220234 9648
rect 220354 9596 220360 9648
rect 220412 9636 220418 9648
rect 220412 9608 221228 9636
rect 220412 9596 220418 9608
rect 174096 9540 175688 9568
rect 175918 9528 175924 9580
rect 175976 9568 175982 9580
rect 176657 9571 176715 9577
rect 176657 9568 176669 9571
rect 175976 9540 176669 9568
rect 175976 9528 175982 9540
rect 176657 9537 176669 9540
rect 176703 9537 176715 9571
rect 176657 9531 176715 9537
rect 177761 9571 177819 9577
rect 177761 9537 177773 9571
rect 177807 9568 177819 9571
rect 177942 9568 177948 9580
rect 177807 9540 177948 9568
rect 177807 9537 177819 9540
rect 177761 9531 177819 9537
rect 177942 9528 177948 9540
rect 178000 9528 178006 9580
rect 178034 9528 178040 9580
rect 178092 9528 178098 9580
rect 179138 9528 179144 9580
rect 179196 9528 179202 9580
rect 179248 9540 179552 9568
rect 154684 9472 155908 9500
rect 108853 9435 108911 9441
rect 108853 9401 108865 9435
rect 108899 9401 108911 9435
rect 108853 9395 108911 9401
rect 109034 9392 109040 9444
rect 109092 9392 109098 9444
rect 109678 9392 109684 9444
rect 109736 9432 109742 9444
rect 111337 9435 111395 9441
rect 111337 9432 111349 9435
rect 109736 9404 111349 9432
rect 109736 9392 109742 9404
rect 111337 9401 111349 9404
rect 111383 9401 111395 9435
rect 111337 9395 111395 9401
rect 112070 9392 112076 9444
rect 112128 9432 112134 9444
rect 114005 9435 114063 9441
rect 114005 9432 114017 9435
rect 112128 9404 114017 9432
rect 112128 9392 112134 9404
rect 114005 9401 114017 9404
rect 114051 9401 114063 9435
rect 114005 9395 114063 9401
rect 116026 9392 116032 9444
rect 116084 9432 116090 9444
rect 120169 9435 120227 9441
rect 120169 9432 120181 9435
rect 116084 9404 120181 9432
rect 116084 9392 116090 9404
rect 120169 9401 120181 9404
rect 120215 9401 120227 9435
rect 120169 9395 120227 9401
rect 121546 9392 121552 9444
rect 121604 9432 121610 9444
rect 132678 9432 132684 9444
rect 121604 9404 132684 9432
rect 121604 9392 121610 9404
rect 132678 9392 132684 9404
rect 132736 9392 132742 9444
rect 142798 9432 142804 9444
rect 137296 9404 142804 9432
rect 103422 9364 103428 9376
rect 89640 9336 103428 9364
rect 88852 9324 88858 9336
rect 103422 9324 103428 9336
rect 103480 9324 103486 9376
rect 103698 9324 103704 9376
rect 103756 9324 103762 9376
rect 104066 9324 104072 9376
rect 104124 9364 104130 9376
rect 108209 9367 108267 9373
rect 108209 9364 108221 9367
rect 104124 9336 108221 9364
rect 104124 9324 104130 9336
rect 108209 9333 108221 9336
rect 108255 9333 108267 9367
rect 108209 9327 108267 9333
rect 108942 9324 108948 9376
rect 109000 9364 109006 9376
rect 109865 9367 109923 9373
rect 109865 9364 109877 9367
rect 109000 9336 109877 9364
rect 109000 9324 109006 9336
rect 109865 9333 109877 9336
rect 109911 9333 109923 9367
rect 109865 9327 109923 9333
rect 110598 9324 110604 9376
rect 110656 9324 110662 9376
rect 112622 9324 112628 9376
rect 112680 9364 112686 9376
rect 112717 9367 112775 9373
rect 112717 9364 112729 9367
rect 112680 9336 112729 9364
rect 112680 9324 112686 9336
rect 112717 9333 112729 9336
rect 112763 9333 112775 9367
rect 112717 9327 112775 9333
rect 113174 9324 113180 9376
rect 113232 9364 113238 9376
rect 113361 9367 113419 9373
rect 113361 9364 113373 9367
rect 113232 9336 113373 9364
rect 113232 9324 113238 9336
rect 113361 9333 113373 9336
rect 113407 9333 113419 9367
rect 113361 9327 113419 9333
rect 115014 9324 115020 9376
rect 115072 9324 115078 9376
rect 115750 9324 115756 9376
rect 115808 9324 115814 9376
rect 115842 9324 115848 9376
rect 115900 9364 115906 9376
rect 116489 9367 116547 9373
rect 116489 9364 116501 9367
rect 115900 9336 116501 9364
rect 115900 9324 115906 9336
rect 116489 9333 116501 9336
rect 116535 9333 116547 9367
rect 116489 9327 116547 9333
rect 117869 9367 117927 9373
rect 117869 9333 117881 9367
rect 117915 9364 117927 9367
rect 117958 9364 117964 9376
rect 117915 9336 117964 9364
rect 117915 9333 117927 9336
rect 117869 9327 117927 9333
rect 117958 9324 117964 9336
rect 118016 9324 118022 9376
rect 118326 9324 118332 9376
rect 118384 9364 118390 9376
rect 118513 9367 118571 9373
rect 118513 9364 118525 9367
rect 118384 9336 118525 9364
rect 118384 9324 118390 9336
rect 118513 9333 118525 9336
rect 118559 9333 118571 9367
rect 118513 9327 118571 9333
rect 119154 9324 119160 9376
rect 119212 9324 119218 9376
rect 120902 9324 120908 9376
rect 120960 9324 120966 9376
rect 128078 9324 128084 9376
rect 128136 9364 128142 9376
rect 128633 9367 128691 9373
rect 128633 9364 128645 9367
rect 128136 9336 128645 9364
rect 128136 9324 128142 9336
rect 128633 9333 128645 9336
rect 128679 9333 128691 9367
rect 128633 9327 128691 9333
rect 128722 9324 128728 9376
rect 128780 9364 128786 9376
rect 137296 9364 137324 9404
rect 142798 9392 142804 9404
rect 142856 9392 142862 9444
rect 143721 9435 143779 9441
rect 143721 9401 143733 9435
rect 143767 9432 143779 9435
rect 145190 9432 145196 9444
rect 143767 9404 145196 9432
rect 143767 9401 143779 9404
rect 143721 9395 143779 9401
rect 145190 9392 145196 9404
rect 145248 9392 145254 9444
rect 146297 9435 146355 9441
rect 146297 9401 146309 9435
rect 146343 9432 146355 9435
rect 148042 9432 148048 9444
rect 146343 9404 148048 9432
rect 146343 9401 146355 9404
rect 146297 9395 146355 9401
rect 148042 9392 148048 9404
rect 148100 9392 148106 9444
rect 150710 9432 150716 9444
rect 148152 9404 150716 9432
rect 128780 9336 137324 9364
rect 128780 9324 128786 9336
rect 138566 9324 138572 9376
rect 138624 9324 138630 9376
rect 139213 9367 139271 9373
rect 139213 9333 139225 9367
rect 139259 9364 139271 9367
rect 140406 9364 140412 9376
rect 139259 9336 140412 9364
rect 139259 9333 139271 9336
rect 139213 9327 139271 9333
rect 140406 9324 140412 9336
rect 140464 9324 140470 9376
rect 140498 9324 140504 9376
rect 140556 9324 140562 9376
rect 140590 9324 140596 9376
rect 140648 9364 140654 9376
rect 141145 9367 141203 9373
rect 141145 9364 141157 9367
rect 140648 9336 141157 9364
rect 140648 9324 140654 9336
rect 141145 9333 141157 9336
rect 141191 9333 141203 9367
rect 141145 9327 141203 9333
rect 141789 9367 141847 9373
rect 141789 9333 141801 9367
rect 141835 9364 141847 9367
rect 142706 9364 142712 9376
rect 141835 9336 142712 9364
rect 141835 9333 141847 9336
rect 141789 9327 141847 9333
rect 142706 9324 142712 9336
rect 142764 9324 142770 9376
rect 143074 9324 143080 9376
rect 143132 9324 143138 9376
rect 144362 9324 144368 9376
rect 144420 9324 144426 9376
rect 145653 9367 145711 9373
rect 145653 9333 145665 9367
rect 145699 9364 145711 9367
rect 145742 9364 145748 9376
rect 145699 9336 145748 9364
rect 145699 9333 145711 9336
rect 145653 9327 145711 9333
rect 145742 9324 145748 9336
rect 145800 9324 145806 9376
rect 146941 9367 146999 9373
rect 146941 9333 146953 9367
rect 146987 9364 146999 9367
rect 148152 9364 148180 9404
rect 150710 9392 150716 9404
rect 150768 9392 150774 9444
rect 151449 9435 151507 9441
rect 151449 9401 151461 9435
rect 151495 9432 151507 9435
rect 153194 9432 153200 9444
rect 151495 9404 153200 9432
rect 151495 9401 151507 9404
rect 151449 9395 151507 9401
rect 153194 9392 153200 9404
rect 153252 9392 153258 9444
rect 154684 9441 154712 9472
rect 156966 9460 156972 9512
rect 157024 9500 157030 9512
rect 157245 9503 157303 9509
rect 157245 9500 157257 9503
rect 157024 9472 157257 9500
rect 157024 9460 157030 9472
rect 157245 9469 157257 9472
rect 157291 9469 157303 9503
rect 157245 9463 157303 9469
rect 158806 9460 158812 9512
rect 158864 9500 158870 9512
rect 159542 9500 159548 9512
rect 158864 9472 159548 9500
rect 158864 9460 158870 9472
rect 159542 9460 159548 9472
rect 159600 9460 159606 9512
rect 159910 9460 159916 9512
rect 159968 9500 159974 9512
rect 160005 9503 160063 9509
rect 160005 9500 160017 9503
rect 159968 9472 160017 9500
rect 159968 9460 159974 9472
rect 160005 9469 160017 9472
rect 160051 9469 160063 9503
rect 160005 9463 160063 9469
rect 161109 9503 161167 9509
rect 161109 9469 161121 9503
rect 161155 9500 161167 9503
rect 161658 9500 161664 9512
rect 161155 9472 161664 9500
rect 161155 9469 161167 9472
rect 161109 9463 161167 9469
rect 161658 9460 161664 9472
rect 161716 9460 161722 9512
rect 161934 9460 161940 9512
rect 161992 9500 161998 9512
rect 162670 9500 162676 9512
rect 161992 9472 162676 9500
rect 161992 9460 161998 9472
rect 162670 9460 162676 9472
rect 162728 9460 162734 9512
rect 163590 9460 163596 9512
rect 163648 9500 163654 9512
rect 163685 9503 163743 9509
rect 163685 9500 163697 9503
rect 163648 9472 163697 9500
rect 163648 9460 163654 9472
rect 163685 9469 163697 9472
rect 163731 9469 163743 9503
rect 163685 9463 163743 9469
rect 164510 9460 164516 9512
rect 164568 9460 164574 9512
rect 165338 9460 165344 9512
rect 165396 9460 165402 9512
rect 165798 9460 165804 9512
rect 165856 9500 165862 9512
rect 166445 9503 166503 9509
rect 166445 9500 166457 9503
rect 165856 9472 166457 9500
rect 165856 9460 165862 9472
rect 166445 9469 166457 9472
rect 166491 9500 166503 9503
rect 167086 9500 167092 9512
rect 166491 9472 167092 9500
rect 166491 9469 166503 9472
rect 166445 9463 166503 9469
rect 167086 9460 167092 9472
rect 167144 9460 167150 9512
rect 169478 9460 169484 9512
rect 169536 9500 169542 9512
rect 169536 9472 169800 9500
rect 169536 9460 169542 9472
rect 153381 9435 153439 9441
rect 153381 9401 153393 9435
rect 153427 9432 153439 9435
rect 154669 9435 154727 9441
rect 153427 9404 154620 9432
rect 153427 9401 153439 9404
rect 153381 9395 153439 9401
rect 146987 9336 148180 9364
rect 146987 9333 146999 9336
rect 146941 9327 146999 9333
rect 148226 9324 148232 9376
rect 148284 9324 148290 9376
rect 148870 9324 148876 9376
rect 148928 9324 148934 9376
rect 149517 9367 149575 9373
rect 149517 9333 149529 9367
rect 149563 9364 149575 9367
rect 150526 9364 150532 9376
rect 149563 9336 150532 9364
rect 149563 9333 149575 9336
rect 149517 9327 149575 9333
rect 150526 9324 150532 9336
rect 150584 9324 150590 9376
rect 150802 9324 150808 9376
rect 150860 9324 150866 9376
rect 152093 9367 152151 9373
rect 152093 9333 152105 9367
rect 152139 9364 152151 9367
rect 153286 9364 153292 9376
rect 152139 9336 153292 9364
rect 152139 9333 152151 9336
rect 152093 9327 152151 9333
rect 153286 9324 153292 9336
rect 153344 9324 153350 9376
rect 154022 9324 154028 9376
rect 154080 9324 154086 9376
rect 154592 9364 154620 9404
rect 154669 9401 154681 9435
rect 154715 9401 154727 9435
rect 154669 9395 154727 9401
rect 156690 9392 156696 9444
rect 156748 9392 156754 9444
rect 169570 9432 169576 9444
rect 157306 9404 169576 9432
rect 155586 9364 155592 9376
rect 154592 9336 155592 9364
rect 155586 9324 155592 9336
rect 155644 9324 155650 9376
rect 155678 9324 155684 9376
rect 155736 9364 155742 9376
rect 157306 9364 157334 9404
rect 169570 9392 169576 9404
rect 169628 9392 169634 9444
rect 169772 9441 169800 9472
rect 171134 9460 171140 9512
rect 171192 9500 171198 9512
rect 172517 9503 172575 9509
rect 172517 9500 172529 9503
rect 171192 9472 172529 9500
rect 171192 9460 171198 9472
rect 172517 9469 172529 9472
rect 172563 9469 172575 9503
rect 172517 9463 172575 9469
rect 172606 9460 172612 9512
rect 172664 9500 172670 9512
rect 179248 9500 179276 9540
rect 172664 9472 179276 9500
rect 179417 9503 179475 9509
rect 172664 9460 172670 9472
rect 179417 9469 179429 9503
rect 179463 9469 179475 9503
rect 179524 9500 179552 9540
rect 180518 9528 180524 9580
rect 180576 9528 180582 9580
rect 180702 9528 180708 9580
rect 180760 9528 180766 9580
rect 181806 9528 181812 9580
rect 181864 9528 181870 9580
rect 182542 9528 182548 9580
rect 182600 9528 182606 9580
rect 183278 9528 183284 9580
rect 183336 9568 183342 9580
rect 184293 9571 184351 9577
rect 184293 9568 184305 9571
rect 183336 9540 184305 9568
rect 183336 9528 183342 9540
rect 184293 9537 184305 9540
rect 184339 9537 184351 9571
rect 184293 9531 184351 9537
rect 185486 9528 185492 9580
rect 185544 9568 185550 9580
rect 186869 9571 186927 9577
rect 186869 9568 186881 9571
rect 185544 9540 186881 9568
rect 185544 9528 185550 9540
rect 186869 9537 186881 9540
rect 186915 9537 186927 9571
rect 186869 9531 186927 9537
rect 188614 9528 188620 9580
rect 188672 9528 188678 9580
rect 190178 9528 190184 9580
rect 190236 9568 190242 9580
rect 190822 9568 190828 9580
rect 190236 9540 190828 9568
rect 190236 9528 190242 9540
rect 190822 9528 190828 9540
rect 190880 9528 190886 9580
rect 192018 9528 192024 9580
rect 192076 9528 192082 9580
rect 192662 9528 192668 9580
rect 192720 9568 192726 9580
rect 192757 9571 192815 9577
rect 192757 9568 192769 9571
rect 192720 9540 192769 9568
rect 192720 9528 192726 9540
rect 192757 9537 192769 9540
rect 192803 9537 192815 9571
rect 192757 9531 192815 9537
rect 194594 9528 194600 9580
rect 194652 9528 194658 9580
rect 195333 9571 195391 9577
rect 195333 9537 195345 9571
rect 195379 9568 195391 9571
rect 195606 9568 195612 9580
rect 195379 9540 195612 9568
rect 195379 9537 195391 9540
rect 195333 9531 195391 9537
rect 195606 9528 195612 9540
rect 195664 9528 195670 9580
rect 196345 9571 196403 9577
rect 196345 9537 196357 9571
rect 196391 9568 196403 9571
rect 197538 9568 197544 9580
rect 196391 9540 197544 9568
rect 196391 9537 196403 9540
rect 196345 9531 196403 9537
rect 197538 9528 197544 9540
rect 197596 9528 197602 9580
rect 197633 9571 197691 9577
rect 197633 9537 197645 9571
rect 197679 9568 197691 9571
rect 197722 9568 197728 9580
rect 197679 9540 197728 9568
rect 197679 9537 197691 9540
rect 197633 9531 197691 9537
rect 197722 9528 197728 9540
rect 197780 9528 197786 9580
rect 197817 9571 197875 9577
rect 197817 9537 197829 9571
rect 197863 9568 197875 9571
rect 198277 9571 198335 9577
rect 198277 9568 198289 9571
rect 197863 9540 198289 9568
rect 197863 9537 197875 9540
rect 197817 9531 197875 9537
rect 198277 9537 198289 9540
rect 198323 9537 198335 9571
rect 198277 9531 198335 9537
rect 202325 9571 202383 9577
rect 202325 9537 202337 9571
rect 202371 9568 202383 9571
rect 202690 9568 202696 9580
rect 202371 9540 202696 9568
rect 202371 9537 202383 9540
rect 202325 9531 202383 9537
rect 202690 9528 202696 9540
rect 202748 9528 202754 9580
rect 203061 9571 203119 9577
rect 203061 9537 203073 9571
rect 203107 9568 203119 9571
rect 203426 9568 203432 9580
rect 203107 9540 203432 9568
rect 203107 9537 203119 9540
rect 203061 9531 203119 9537
rect 203426 9528 203432 9540
rect 203484 9528 203490 9580
rect 205818 9528 205824 9580
rect 205876 9528 205882 9580
rect 206554 9528 206560 9580
rect 206612 9528 206618 9580
rect 207658 9528 207664 9580
rect 207716 9528 207722 9580
rect 208302 9528 208308 9580
rect 208360 9528 208366 9580
rect 208946 9528 208952 9580
rect 209004 9528 209010 9580
rect 209314 9528 209320 9580
rect 209372 9568 209378 9580
rect 210237 9571 210295 9577
rect 210237 9568 210249 9571
rect 209372 9540 210249 9568
rect 209372 9528 209378 9540
rect 210237 9537 210249 9540
rect 210283 9537 210295 9571
rect 210237 9531 210295 9537
rect 210878 9528 210884 9580
rect 210936 9528 210942 9580
rect 211154 9528 211160 9580
rect 211212 9568 211218 9580
rect 211525 9571 211583 9577
rect 211525 9568 211537 9571
rect 211212 9540 211537 9568
rect 211212 9528 211218 9540
rect 211525 9537 211537 9540
rect 211571 9537 211583 9571
rect 211525 9531 211583 9537
rect 212534 9528 212540 9580
rect 212592 9568 212598 9580
rect 212813 9571 212871 9577
rect 212813 9568 212825 9571
rect 212592 9540 212825 9568
rect 212592 9528 212598 9540
rect 212813 9537 212825 9540
rect 212859 9537 212871 9571
rect 212813 9531 212871 9537
rect 213454 9528 213460 9580
rect 213512 9528 213518 9580
rect 213914 9528 213920 9580
rect 213972 9568 213978 9580
rect 214101 9571 214159 9577
rect 214101 9568 214113 9571
rect 213972 9540 214113 9568
rect 213972 9528 213978 9540
rect 214101 9537 214113 9540
rect 214147 9537 214159 9571
rect 214101 9531 214159 9537
rect 214466 9528 214472 9580
rect 214524 9568 214530 9580
rect 215389 9571 215447 9577
rect 215389 9568 215401 9571
rect 214524 9540 215401 9568
rect 214524 9528 214530 9540
rect 215389 9537 215401 9540
rect 215435 9537 215447 9571
rect 215389 9531 215447 9537
rect 215478 9528 215484 9580
rect 215536 9568 215542 9580
rect 216033 9571 216091 9577
rect 216033 9568 216045 9571
rect 215536 9540 216045 9568
rect 215536 9528 215542 9540
rect 216033 9537 216045 9540
rect 216079 9537 216091 9571
rect 216033 9531 216091 9537
rect 216674 9528 216680 9580
rect 216732 9528 216738 9580
rect 217962 9528 217968 9580
rect 218020 9528 218026 9580
rect 218606 9528 218612 9580
rect 218664 9528 218670 9580
rect 219250 9528 219256 9580
rect 219308 9528 219314 9580
rect 220538 9528 220544 9580
rect 220596 9528 220602 9580
rect 221200 9577 221228 9608
rect 229002 9596 229008 9648
rect 229060 9636 229066 9648
rect 229060 9608 255176 9636
rect 229060 9596 229066 9608
rect 221185 9571 221243 9577
rect 221185 9537 221197 9571
rect 221231 9537 221243 9571
rect 221185 9531 221243 9537
rect 221826 9528 221832 9580
rect 221884 9528 221890 9580
rect 223114 9528 223120 9580
rect 223172 9528 223178 9580
rect 223758 9528 223764 9580
rect 223816 9568 223822 9580
rect 223853 9571 223911 9577
rect 223853 9568 223865 9571
rect 223816 9540 223865 9568
rect 223816 9528 223822 9540
rect 223853 9537 223865 9540
rect 223899 9537 223911 9571
rect 223853 9531 223911 9537
rect 223942 9528 223948 9580
rect 224000 9568 224006 9580
rect 224773 9575 224831 9581
rect 224773 9574 224785 9575
rect 224696 9568 224785 9574
rect 224000 9546 224785 9568
rect 224000 9540 224724 9546
rect 224773 9541 224785 9546
rect 224819 9541 224831 9575
rect 224000 9528 224006 9540
rect 224773 9535 224831 9541
rect 224862 9528 224868 9580
rect 224920 9568 224926 9580
rect 227806 9568 227812 9580
rect 224920 9540 227812 9568
rect 224920 9528 224926 9540
rect 227806 9528 227812 9540
rect 227864 9528 227870 9580
rect 228085 9571 228143 9577
rect 228085 9537 228097 9571
rect 228131 9568 228143 9571
rect 228358 9568 228364 9580
rect 228131 9540 228364 9568
rect 228131 9537 228143 9540
rect 228085 9531 228143 9537
rect 228358 9528 228364 9540
rect 228416 9528 228422 9580
rect 228450 9528 228456 9580
rect 228508 9568 228514 9580
rect 228821 9571 228879 9577
rect 228821 9568 228833 9571
rect 228508 9540 228833 9568
rect 228508 9528 228514 9540
rect 228821 9537 228833 9540
rect 228867 9537 228879 9571
rect 228821 9531 228879 9537
rect 229649 9571 229707 9577
rect 229649 9537 229661 9571
rect 229695 9568 229707 9571
rect 230014 9568 230020 9580
rect 229695 9540 230020 9568
rect 229695 9537 229707 9540
rect 229649 9531 229707 9537
rect 230014 9528 230020 9540
rect 230072 9528 230078 9580
rect 230658 9528 230664 9580
rect 230716 9528 230722 9580
rect 230842 9528 230848 9580
rect 230900 9528 230906 9580
rect 231765 9571 231823 9577
rect 231765 9537 231777 9571
rect 231811 9568 231823 9571
rect 232314 9568 232320 9580
rect 231811 9540 232320 9568
rect 231811 9537 231823 9540
rect 231765 9531 231823 9537
rect 232314 9528 232320 9540
rect 232372 9528 232378 9580
rect 233237 9571 233295 9577
rect 233237 9537 233249 9571
rect 233283 9568 233295 9571
rect 233970 9568 233976 9580
rect 233283 9540 233976 9568
rect 233283 9537 233295 9540
rect 233237 9531 233295 9537
rect 233970 9528 233976 9540
rect 234028 9528 234034 9580
rect 234798 9528 234804 9580
rect 234856 9528 234862 9580
rect 234985 9571 235043 9577
rect 234985 9537 234997 9571
rect 235031 9568 235043 9571
rect 235813 9571 235871 9577
rect 235813 9568 235825 9571
rect 235031 9540 235825 9568
rect 235031 9537 235043 9540
rect 234985 9531 235043 9537
rect 235813 9537 235825 9540
rect 235859 9537 235871 9571
rect 235813 9531 235871 9537
rect 239950 9528 239956 9580
rect 240008 9528 240014 9580
rect 240962 9528 240968 9580
rect 241020 9528 241026 9580
rect 242342 9528 242348 9580
rect 242400 9528 242406 9580
rect 242894 9528 242900 9580
rect 242952 9568 242958 9580
rect 243633 9571 243691 9577
rect 243633 9568 243645 9571
rect 242952 9540 243645 9568
rect 242952 9528 242958 9540
rect 243633 9537 243645 9540
rect 243679 9537 243691 9571
rect 244369 9571 244427 9577
rect 244369 9568 244381 9571
rect 243633 9531 243691 9537
rect 243924 9540 244381 9568
rect 181993 9503 182051 9509
rect 181993 9500 182005 9503
rect 179524 9472 182005 9500
rect 179417 9463 179475 9469
rect 181993 9469 182005 9472
rect 182039 9469 182051 9503
rect 181993 9463 182051 9469
rect 182821 9503 182879 9509
rect 182821 9469 182833 9503
rect 182867 9469 182879 9503
rect 182821 9463 182879 9469
rect 169757 9435 169815 9441
rect 169757 9401 169769 9435
rect 169803 9401 169815 9435
rect 169757 9395 169815 9401
rect 169846 9392 169852 9444
rect 169904 9432 169910 9444
rect 179432 9432 179460 9463
rect 169904 9404 179460 9432
rect 169904 9392 169910 9404
rect 155736 9336 157334 9364
rect 157613 9367 157671 9373
rect 155736 9324 155742 9336
rect 157613 9333 157625 9367
rect 157659 9364 157671 9367
rect 158530 9364 158536 9376
rect 157659 9336 158536 9364
rect 157659 9333 157671 9336
rect 157613 9327 157671 9333
rect 158530 9324 158536 9336
rect 158588 9324 158594 9376
rect 159177 9367 159235 9373
rect 159177 9333 159189 9367
rect 159223 9364 159235 9367
rect 160002 9364 160008 9376
rect 159223 9336 160008 9364
rect 159223 9333 159235 9336
rect 159177 9327 159235 9333
rect 160002 9324 160008 9336
rect 160060 9324 160066 9376
rect 161477 9367 161535 9373
rect 161477 9333 161489 9367
rect 161523 9364 161535 9367
rect 162210 9364 162216 9376
rect 161523 9336 162216 9364
rect 161523 9333 161535 9336
rect 161477 9327 161535 9333
rect 162210 9324 162216 9336
rect 162268 9324 162274 9376
rect 162305 9367 162363 9373
rect 162305 9333 162317 9367
rect 162351 9364 162363 9367
rect 162946 9364 162952 9376
rect 162351 9336 162952 9364
rect 162351 9333 162363 9336
rect 162305 9327 162363 9333
rect 162946 9324 162952 9336
rect 163004 9324 163010 9376
rect 163133 9367 163191 9373
rect 163133 9333 163145 9367
rect 163179 9364 163191 9367
rect 163682 9364 163688 9376
rect 163179 9336 163688 9364
rect 163179 9333 163191 9336
rect 163133 9327 163191 9333
rect 163682 9324 163688 9336
rect 163740 9324 163746 9376
rect 164053 9367 164111 9373
rect 164053 9333 164065 9367
rect 164099 9364 164111 9367
rect 164418 9364 164424 9376
rect 164099 9336 164424 9364
rect 164099 9333 164111 9336
rect 164053 9327 164111 9333
rect 164418 9324 164424 9336
rect 164476 9324 164482 9376
rect 164881 9367 164939 9373
rect 164881 9333 164893 9367
rect 164927 9364 164939 9367
rect 165154 9364 165160 9376
rect 164927 9336 165160 9364
rect 164927 9333 164939 9336
rect 164881 9327 164939 9333
rect 165154 9324 165160 9336
rect 165212 9324 165218 9376
rect 165709 9367 165767 9373
rect 165709 9333 165721 9367
rect 165755 9364 165767 9367
rect 165890 9364 165896 9376
rect 165755 9336 165896 9364
rect 165755 9333 165767 9336
rect 165709 9327 165767 9333
rect 165890 9324 165896 9336
rect 165948 9324 165954 9376
rect 166718 9324 166724 9376
rect 166776 9364 166782 9376
rect 166813 9367 166871 9373
rect 166813 9364 166825 9367
rect 166776 9336 166825 9364
rect 166776 9324 166782 9336
rect 166813 9333 166825 9336
rect 166859 9333 166871 9367
rect 166813 9327 166871 9333
rect 169662 9324 169668 9376
rect 169720 9364 169726 9376
rect 174219 9367 174277 9373
rect 174219 9364 174231 9367
rect 169720 9336 174231 9364
rect 169720 9324 169726 9336
rect 174219 9333 174231 9336
rect 174265 9333 174277 9367
rect 174219 9327 174277 9333
rect 175550 9324 175556 9376
rect 175608 9364 175614 9376
rect 176749 9367 176807 9373
rect 176749 9364 176761 9367
rect 175608 9336 176761 9364
rect 175608 9324 175614 9336
rect 176749 9333 176761 9336
rect 176795 9333 176807 9367
rect 176749 9327 176807 9333
rect 178402 9324 178408 9376
rect 178460 9364 178466 9376
rect 182836 9364 182864 9463
rect 184566 9460 184572 9512
rect 184624 9460 184630 9512
rect 186406 9460 186412 9512
rect 186464 9500 186470 9512
rect 187145 9503 187203 9509
rect 187145 9500 187157 9503
rect 186464 9472 187157 9500
rect 186464 9460 186470 9472
rect 187145 9469 187157 9472
rect 187191 9469 187203 9503
rect 187145 9463 187203 9469
rect 187694 9460 187700 9512
rect 187752 9500 187758 9512
rect 189445 9503 189503 9509
rect 189445 9500 189457 9503
rect 187752 9472 189457 9500
rect 187752 9460 187758 9472
rect 189445 9469 189457 9472
rect 189491 9469 189503 9503
rect 189445 9463 189503 9469
rect 189721 9503 189779 9509
rect 189721 9469 189733 9503
rect 189767 9469 189779 9503
rect 189721 9463 189779 9469
rect 197449 9503 197507 9509
rect 197449 9469 197461 9503
rect 197495 9500 197507 9503
rect 197906 9500 197912 9512
rect 197495 9472 197912 9500
rect 197495 9469 197507 9472
rect 197449 9463 197507 9469
rect 184842 9392 184848 9444
rect 184900 9432 184906 9444
rect 189736 9432 189764 9463
rect 197906 9460 197912 9472
rect 197964 9500 197970 9512
rect 219894 9500 219900 9512
rect 197964 9472 219900 9500
rect 197964 9460 197970 9472
rect 219894 9460 219900 9472
rect 219952 9460 219958 9512
rect 219986 9460 219992 9512
rect 220044 9500 220050 9512
rect 220044 9472 229968 9500
rect 220044 9460 220050 9472
rect 184900 9404 189764 9432
rect 184900 9392 184906 9404
rect 191374 9392 191380 9444
rect 191432 9432 191438 9444
rect 192205 9435 192263 9441
rect 192205 9432 192217 9435
rect 191432 9404 192217 9432
rect 191432 9392 191438 9404
rect 192205 9401 192217 9404
rect 192251 9401 192263 9435
rect 192205 9395 192263 9401
rect 192938 9392 192944 9444
rect 192996 9392 193002 9444
rect 194318 9392 194324 9444
rect 194376 9432 194382 9444
rect 194781 9435 194839 9441
rect 194781 9432 194793 9435
rect 194376 9404 194793 9432
rect 194376 9392 194382 9404
rect 194781 9401 194793 9404
rect 194827 9401 194839 9435
rect 194781 9395 194839 9401
rect 195514 9392 195520 9444
rect 195572 9392 195578 9444
rect 196526 9392 196532 9444
rect 196584 9392 196590 9444
rect 197262 9392 197268 9444
rect 197320 9432 197326 9444
rect 198461 9435 198519 9441
rect 198461 9432 198473 9435
rect 197320 9404 198473 9432
rect 197320 9392 197326 9404
rect 198461 9401 198473 9404
rect 198507 9401 198519 9435
rect 198461 9395 198519 9401
rect 202506 9392 202512 9444
rect 202564 9392 202570 9444
rect 207014 9392 207020 9444
rect 207072 9432 207078 9444
rect 208121 9435 208179 9441
rect 208121 9432 208133 9435
rect 207072 9404 208133 9432
rect 207072 9392 207078 9404
rect 208121 9401 208133 9404
rect 208167 9401 208179 9435
rect 208121 9395 208179 9401
rect 213917 9435 213975 9441
rect 213917 9401 213929 9435
rect 213963 9432 213975 9435
rect 215018 9432 215024 9444
rect 213963 9404 215024 9432
rect 213963 9401 213975 9404
rect 213917 9395 213975 9401
rect 215018 9392 215024 9404
rect 215076 9392 215082 9444
rect 215110 9392 215116 9444
rect 215168 9432 215174 9444
rect 215168 9404 227024 9432
rect 215168 9392 215174 9404
rect 178460 9336 182864 9364
rect 178460 9324 178466 9336
rect 186314 9324 186320 9376
rect 186372 9364 186378 9376
rect 188433 9367 188491 9373
rect 188433 9364 188445 9367
rect 186372 9336 188445 9364
rect 186372 9324 186378 9336
rect 188433 9333 188445 9336
rect 188479 9333 188491 9367
rect 188433 9327 188491 9333
rect 190914 9324 190920 9376
rect 190972 9324 190978 9376
rect 194502 9324 194508 9376
rect 194560 9364 194566 9376
rect 197170 9364 197176 9376
rect 194560 9336 197176 9364
rect 194560 9324 194566 9336
rect 197170 9324 197176 9336
rect 197228 9324 197234 9376
rect 202414 9324 202420 9376
rect 202472 9364 202478 9376
rect 203245 9367 203303 9373
rect 203245 9364 203257 9367
rect 202472 9336 203257 9364
rect 202472 9324 202478 9336
rect 203245 9333 203257 9336
rect 203291 9333 203303 9367
rect 203245 9327 203303 9333
rect 206373 9367 206431 9373
rect 206373 9333 206385 9367
rect 206419 9364 206431 9367
rect 206830 9364 206836 9376
rect 206419 9336 206836 9364
rect 206419 9333 206431 9336
rect 206373 9327 206431 9333
rect 206830 9324 206836 9336
rect 206888 9324 206894 9376
rect 207474 9324 207480 9376
rect 207532 9324 207538 9376
rect 208762 9324 208768 9376
rect 208820 9324 208826 9376
rect 210050 9324 210056 9376
rect 210108 9324 210114 9376
rect 210694 9324 210700 9376
rect 210752 9324 210758 9376
rect 211341 9367 211399 9373
rect 211341 9333 211353 9367
rect 211387 9364 211399 9367
rect 212442 9364 212448 9376
rect 211387 9336 212448 9364
rect 211387 9333 211399 9336
rect 211341 9327 211399 9333
rect 212442 9324 212448 9336
rect 212500 9324 212506 9376
rect 212626 9324 212632 9376
rect 212684 9324 212690 9376
rect 213270 9324 213276 9376
rect 213328 9324 213334 9376
rect 214834 9324 214840 9376
rect 214892 9364 214898 9376
rect 215205 9367 215263 9373
rect 215205 9364 215217 9367
rect 214892 9336 215217 9364
rect 214892 9324 214898 9336
rect 215205 9333 215217 9336
rect 215251 9333 215263 9367
rect 215205 9327 215263 9333
rect 216493 9367 216551 9373
rect 216493 9333 216505 9367
rect 216539 9364 216551 9367
rect 217502 9364 217508 9376
rect 216539 9336 217508 9364
rect 216539 9333 216551 9336
rect 216493 9327 216551 9333
rect 217502 9324 217508 9336
rect 217560 9324 217566 9376
rect 217778 9324 217784 9376
rect 217836 9324 217842 9376
rect 218422 9324 218428 9376
rect 218480 9324 218486 9376
rect 219069 9367 219127 9373
rect 219069 9333 219081 9367
rect 219115 9364 219127 9367
rect 219342 9364 219348 9376
rect 219115 9336 219348 9364
rect 219115 9333 219127 9336
rect 219069 9327 219127 9333
rect 219342 9324 219348 9336
rect 219400 9324 219406 9376
rect 220354 9324 220360 9376
rect 220412 9324 220418 9376
rect 220998 9324 221004 9376
rect 221056 9324 221062 9376
rect 221642 9324 221648 9376
rect 221700 9324 221706 9376
rect 222930 9324 222936 9376
rect 222988 9324 222994 9376
rect 224034 9324 224040 9376
rect 224092 9324 224098 9376
rect 224589 9367 224647 9373
rect 224589 9333 224601 9367
rect 224635 9364 224647 9367
rect 225230 9364 225236 9376
rect 224635 9336 225236 9364
rect 224635 9333 224647 9336
rect 224589 9327 224647 9333
rect 225230 9324 225236 9336
rect 225288 9324 225294 9376
rect 226996 9364 227024 9404
rect 228266 9392 228272 9444
rect 228324 9392 228330 9444
rect 229002 9392 229008 9444
rect 229060 9392 229066 9444
rect 229830 9392 229836 9444
rect 229888 9392 229894 9444
rect 229940 9432 229968 9472
rect 230290 9460 230296 9512
rect 230348 9500 230354 9512
rect 234617 9503 234675 9509
rect 234617 9500 234629 9503
rect 230348 9472 234629 9500
rect 230348 9460 230354 9472
rect 234617 9469 234629 9472
rect 234663 9500 234675 9503
rect 235902 9500 235908 9512
rect 234663 9472 235908 9500
rect 234663 9469 234675 9472
rect 234617 9463 234675 9469
rect 235902 9460 235908 9472
rect 235960 9500 235966 9512
rect 235960 9472 237236 9500
rect 235960 9460 235966 9472
rect 229940 9404 231854 9432
rect 230290 9364 230296 9376
rect 226996 9336 230296 9364
rect 230290 9324 230296 9336
rect 230348 9324 230354 9376
rect 231029 9367 231087 9373
rect 231029 9333 231041 9367
rect 231075 9364 231087 9367
rect 231486 9364 231492 9376
rect 231075 9336 231492 9364
rect 231075 9333 231087 9336
rect 231029 9327 231087 9333
rect 231486 9324 231492 9336
rect 231544 9324 231550 9376
rect 231826 9364 231854 9404
rect 231946 9392 231952 9444
rect 232004 9392 232010 9444
rect 233418 9392 233424 9444
rect 233476 9392 233482 9444
rect 235994 9392 236000 9444
rect 236052 9392 236058 9444
rect 237208 9432 237236 9472
rect 237282 9460 237288 9512
rect 237340 9500 237346 9512
rect 241241 9503 241299 9509
rect 241241 9500 241253 9503
rect 237340 9472 241253 9500
rect 237340 9460 237346 9472
rect 241241 9469 241253 9472
rect 241287 9469 241299 9503
rect 241241 9463 241299 9469
rect 242526 9460 242532 9512
rect 242584 9460 242590 9512
rect 243446 9460 243452 9512
rect 243504 9500 243510 9512
rect 243924 9500 243952 9540
rect 244369 9537 244381 9540
rect 244415 9537 244427 9571
rect 244369 9531 244427 9537
rect 245105 9571 245163 9577
rect 245105 9537 245117 9571
rect 245151 9537 245163 9571
rect 245105 9531 245163 9537
rect 243504 9472 243952 9500
rect 243504 9460 243510 9472
rect 244182 9460 244188 9512
rect 244240 9500 244246 9512
rect 245120 9500 245148 9531
rect 246390 9528 246396 9580
rect 246448 9528 246454 9580
rect 247954 9528 247960 9580
rect 248012 9528 248018 9580
rect 249334 9528 249340 9580
rect 249392 9528 249398 9580
rect 251542 9528 251548 9580
rect 251600 9528 251606 9580
rect 253842 9528 253848 9580
rect 253900 9528 253906 9580
rect 244240 9472 245148 9500
rect 244240 9460 244246 9472
rect 246666 9460 246672 9512
rect 246724 9460 246730 9512
rect 249610 9460 249616 9512
rect 249668 9460 249674 9512
rect 249702 9460 249708 9512
rect 249760 9500 249766 9512
rect 251821 9503 251879 9509
rect 251821 9500 251833 9503
rect 249760 9472 251833 9500
rect 249760 9460 249766 9472
rect 251821 9469 251833 9472
rect 251867 9469 251879 9503
rect 251821 9463 251879 9469
rect 254118 9460 254124 9512
rect 254176 9460 254182 9512
rect 255148 9500 255176 9608
rect 255222 9596 255228 9648
rect 255280 9636 255286 9648
rect 260024 9636 260052 9667
rect 266262 9664 266268 9716
rect 266320 9664 266326 9716
rect 266998 9664 267004 9716
rect 267056 9704 267062 9716
rect 270402 9704 270408 9716
rect 267056 9676 270408 9704
rect 267056 9664 267062 9676
rect 270402 9664 270408 9676
rect 270460 9664 270466 9716
rect 255280 9608 260052 9636
rect 255280 9596 255286 9608
rect 264974 9596 264980 9648
rect 265032 9636 265038 9648
rect 265621 9639 265679 9645
rect 265621 9636 265633 9639
rect 265032 9608 265633 9636
rect 265032 9596 265038 9608
rect 265621 9605 265633 9608
rect 265667 9605 265679 9639
rect 268105 9639 268163 9645
rect 265621 9599 265679 9605
rect 266004 9608 267136 9636
rect 255314 9528 255320 9580
rect 255372 9568 255378 9580
rect 256421 9571 256479 9577
rect 256421 9568 256433 9571
rect 255372 9540 256433 9568
rect 255372 9528 255378 9540
rect 256421 9537 256433 9540
rect 256467 9537 256479 9571
rect 257890 9568 257896 9580
rect 256421 9531 256479 9537
rect 256620 9540 257896 9568
rect 256620 9500 256648 9540
rect 257890 9528 257896 9540
rect 257948 9528 257954 9580
rect 257982 9528 257988 9580
rect 258040 9528 258046 9580
rect 258077 9571 258135 9577
rect 258077 9537 258089 9571
rect 258123 9537 258135 9571
rect 258077 9531 258135 9537
rect 258997 9571 259055 9577
rect 258997 9537 259009 9571
rect 259043 9568 259055 9571
rect 259362 9568 259368 9580
rect 259043 9540 259368 9568
rect 259043 9537 259055 9540
rect 258997 9531 259055 9537
rect 255148 9472 256648 9500
rect 256697 9503 256755 9509
rect 256697 9469 256709 9503
rect 256743 9500 256755 9503
rect 256878 9500 256884 9512
rect 256743 9472 256884 9500
rect 256743 9469 256755 9472
rect 256697 9463 256755 9469
rect 256878 9460 256884 9472
rect 256936 9460 256942 9512
rect 258092 9500 258120 9531
rect 259362 9528 259368 9540
rect 259420 9528 259426 9580
rect 260190 9528 260196 9580
rect 260248 9528 260254 9580
rect 260837 9571 260895 9577
rect 260837 9568 260849 9571
rect 260576 9540 260849 9568
rect 259178 9500 259184 9512
rect 258092 9472 259184 9500
rect 259178 9460 259184 9472
rect 259236 9500 259242 9512
rect 260576 9500 260604 9540
rect 260837 9537 260849 9540
rect 260883 9568 260895 9571
rect 261757 9571 261815 9577
rect 261757 9568 261769 9571
rect 260883 9540 261769 9568
rect 260883 9537 260895 9540
rect 260837 9531 260895 9537
rect 261757 9537 261769 9540
rect 261803 9568 261815 9571
rect 262585 9571 262643 9577
rect 262585 9568 262597 9571
rect 261803 9540 262597 9568
rect 261803 9537 261815 9540
rect 261757 9531 261815 9537
rect 262585 9537 262597 9540
rect 262631 9568 262643 9571
rect 263413 9571 263471 9577
rect 263413 9568 263425 9571
rect 262631 9540 263425 9568
rect 262631 9537 262643 9540
rect 262585 9531 262643 9537
rect 263413 9537 263425 9540
rect 263459 9568 263471 9571
rect 263594 9568 263600 9580
rect 263459 9540 263600 9568
rect 263459 9537 263471 9540
rect 263413 9531 263471 9537
rect 263594 9528 263600 9540
rect 263652 9528 263658 9580
rect 264241 9571 264299 9577
rect 264241 9537 264253 9571
rect 264287 9568 264299 9571
rect 264422 9568 264428 9580
rect 264287 9540 264428 9568
rect 264287 9537 264299 9540
rect 264241 9531 264299 9537
rect 264422 9528 264428 9540
rect 264480 9568 264486 9580
rect 264885 9571 264943 9577
rect 264885 9568 264897 9571
rect 264480 9540 264897 9568
rect 264480 9528 264486 9540
rect 264885 9537 264897 9540
rect 264931 9537 264943 9571
rect 264885 9531 264943 9537
rect 265250 9528 265256 9580
rect 265308 9568 265314 9580
rect 266004 9568 266032 9608
rect 267108 9577 267136 9608
rect 268105 9605 268117 9639
rect 268151 9636 268163 9639
rect 269942 9636 269948 9648
rect 268151 9608 269948 9636
rect 268151 9605 268163 9608
rect 268105 9599 268163 9605
rect 269942 9596 269948 9608
rect 270000 9596 270006 9648
rect 265308 9540 266032 9568
rect 266081 9571 266139 9577
rect 265308 9528 265314 9540
rect 266081 9537 266093 9571
rect 266127 9537 266139 9571
rect 266081 9531 266139 9537
rect 267093 9571 267151 9577
rect 267093 9537 267105 9571
rect 267139 9568 267151 9571
rect 267642 9568 267648 9580
rect 267139 9540 267648 9568
rect 267139 9537 267151 9540
rect 267093 9531 267151 9537
rect 259236 9472 260604 9500
rect 260653 9503 260711 9509
rect 259236 9460 259242 9472
rect 260653 9469 260665 9503
rect 260699 9500 260711 9503
rect 261386 9500 261392 9512
rect 260699 9472 261392 9500
rect 260699 9469 260711 9472
rect 260653 9463 260711 9469
rect 237208 9404 238984 9432
rect 238846 9364 238852 9376
rect 231826 9336 238852 9364
rect 238846 9324 238852 9336
rect 238904 9324 238910 9376
rect 238956 9364 238984 9404
rect 240134 9392 240140 9444
rect 240192 9432 240198 9444
rect 243817 9435 243875 9441
rect 243817 9432 243829 9435
rect 240192 9404 243829 9432
rect 240192 9392 240198 9404
rect 243817 9401 243829 9404
rect 243863 9401 243875 9435
rect 258626 9432 258632 9444
rect 243817 9395 243875 9401
rect 243924 9404 258632 9432
rect 243924 9364 243952 9404
rect 258626 9392 258632 9404
rect 258684 9392 258690 9444
rect 258718 9392 258724 9444
rect 258776 9432 258782 9444
rect 260668 9432 260696 9463
rect 261386 9460 261392 9472
rect 261444 9460 261450 9512
rect 261570 9460 261576 9512
rect 261628 9460 261634 9512
rect 262122 9460 262128 9512
rect 262180 9500 262186 9512
rect 262401 9503 262459 9509
rect 262401 9500 262413 9503
rect 262180 9472 262413 9500
rect 262180 9460 262186 9472
rect 262401 9469 262413 9472
rect 262447 9469 262459 9503
rect 262401 9463 262459 9469
rect 263226 9460 263232 9512
rect 263284 9500 263290 9512
rect 263962 9500 263968 9512
rect 263284 9472 263968 9500
rect 263284 9460 263290 9472
rect 263962 9460 263968 9472
rect 264020 9460 264026 9512
rect 264698 9460 264704 9512
rect 264756 9500 264762 9512
rect 265069 9503 265127 9509
rect 265069 9500 265081 9503
rect 264756 9472 265081 9500
rect 264756 9460 264762 9472
rect 265069 9469 265081 9472
rect 265115 9469 265127 9503
rect 265069 9463 265127 9469
rect 265437 9503 265495 9509
rect 265437 9469 265449 9503
rect 265483 9500 265495 9503
rect 266096 9500 266124 9531
rect 267642 9528 267648 9540
rect 267700 9568 267706 9580
rect 267921 9571 267979 9577
rect 267921 9568 267933 9571
rect 267700 9540 267933 9568
rect 267700 9528 267706 9540
rect 267921 9537 267933 9540
rect 267967 9568 267979 9571
rect 268749 9571 268807 9577
rect 268749 9568 268761 9571
rect 267967 9540 268761 9568
rect 267967 9537 267979 9540
rect 267921 9531 267979 9537
rect 268749 9537 268761 9540
rect 268795 9537 268807 9571
rect 268749 9531 268807 9537
rect 268930 9528 268936 9580
rect 268988 9568 268994 9580
rect 269117 9571 269175 9577
rect 269117 9568 269129 9571
rect 268988 9540 269129 9568
rect 268988 9528 268994 9540
rect 269117 9537 269129 9540
rect 269163 9537 269175 9571
rect 269117 9531 269175 9537
rect 269577 9571 269635 9577
rect 269577 9537 269589 9571
rect 269623 9537 269635 9571
rect 269577 9531 269635 9537
rect 270129 9571 270187 9577
rect 270129 9537 270141 9571
rect 270175 9568 270187 9571
rect 270494 9568 270500 9580
rect 270175 9540 270500 9568
rect 270175 9537 270187 9540
rect 270129 9531 270187 9537
rect 265483 9472 266124 9500
rect 265483 9469 265495 9472
rect 265437 9463 265495 9469
rect 258776 9404 260696 9432
rect 258776 9392 258782 9404
rect 260834 9392 260840 9444
rect 260892 9432 260898 9444
rect 263686 9432 263692 9444
rect 260892 9404 263692 9432
rect 260892 9392 260898 9404
rect 263686 9392 263692 9404
rect 263744 9392 263750 9444
rect 263778 9392 263784 9444
rect 263836 9432 263842 9444
rect 264425 9435 264483 9441
rect 264425 9432 264437 9435
rect 263836 9404 264437 9432
rect 263836 9392 263842 9404
rect 264425 9401 264437 9404
rect 264471 9401 264483 9435
rect 265084 9432 265112 9463
rect 266906 9460 266912 9512
rect 266964 9500 266970 9512
rect 267458 9500 267464 9512
rect 266964 9472 267464 9500
rect 266964 9460 266970 9472
rect 267458 9460 267464 9472
rect 267516 9460 267522 9512
rect 267550 9460 267556 9512
rect 267608 9500 267614 9512
rect 267737 9503 267795 9509
rect 267737 9500 267749 9503
rect 267608 9472 267749 9500
rect 267608 9460 267614 9472
rect 267737 9469 267749 9472
rect 267783 9500 267795 9503
rect 268470 9500 268476 9512
rect 267783 9472 268476 9500
rect 267783 9469 267795 9472
rect 267737 9463 267795 9469
rect 268470 9460 268476 9472
rect 268528 9460 268534 9512
rect 268562 9460 268568 9512
rect 268620 9460 268626 9512
rect 268838 9460 268844 9512
rect 268896 9500 268902 9512
rect 269592 9500 269620 9531
rect 270494 9528 270500 9540
rect 270552 9528 270558 9580
rect 268896 9472 269620 9500
rect 268896 9460 268902 9472
rect 269850 9460 269856 9512
rect 269908 9500 269914 9512
rect 270405 9503 270463 9509
rect 270405 9500 270417 9503
rect 269908 9472 270417 9500
rect 269908 9460 269914 9472
rect 270405 9469 270417 9472
rect 270451 9469 270463 9503
rect 270405 9463 270463 9469
rect 265805 9435 265863 9441
rect 265805 9432 265817 9435
rect 265084 9404 265817 9432
rect 264425 9395 264483 9401
rect 265805 9401 265817 9404
rect 265851 9401 265863 9435
rect 268746 9432 268752 9444
rect 265805 9395 265863 9401
rect 266280 9404 268752 9432
rect 238956 9336 243952 9364
rect 243998 9324 244004 9376
rect 244056 9364 244062 9376
rect 244461 9367 244519 9373
rect 244461 9364 244473 9367
rect 244056 9336 244473 9364
rect 244056 9324 244062 9336
rect 244461 9333 244473 9336
rect 244507 9333 244519 9367
rect 244461 9327 244519 9333
rect 245194 9324 245200 9376
rect 245252 9324 245258 9376
rect 245562 9324 245568 9376
rect 245620 9364 245626 9376
rect 248049 9367 248107 9373
rect 248049 9364 248061 9367
rect 245620 9336 248061 9364
rect 245620 9324 245626 9336
rect 248049 9333 248061 9336
rect 248095 9333 248107 9367
rect 248049 9327 248107 9333
rect 258074 9324 258080 9376
rect 258132 9364 258138 9376
rect 258261 9367 258319 9373
rect 258261 9364 258273 9367
rect 258132 9336 258273 9364
rect 258132 9324 258138 9336
rect 258261 9333 258273 9336
rect 258307 9333 258319 9367
rect 258261 9327 258319 9333
rect 261021 9367 261079 9373
rect 261021 9333 261033 9367
rect 261067 9364 261079 9367
rect 261478 9364 261484 9376
rect 261067 9336 261484 9364
rect 261067 9333 261079 9336
rect 261021 9327 261079 9333
rect 261478 9324 261484 9336
rect 261536 9324 261542 9376
rect 261570 9324 261576 9376
rect 261628 9364 261634 9376
rect 261941 9367 261999 9373
rect 261941 9364 261953 9367
rect 261628 9336 261953 9364
rect 261628 9324 261634 9336
rect 261941 9333 261953 9336
rect 261987 9333 261999 9367
rect 261941 9327 261999 9333
rect 262306 9324 262312 9376
rect 262364 9364 262370 9376
rect 262769 9367 262827 9373
rect 262769 9364 262781 9367
rect 262364 9336 262781 9364
rect 262364 9324 262370 9336
rect 262769 9333 262781 9336
rect 262815 9333 262827 9367
rect 262769 9327 262827 9333
rect 263597 9367 263655 9373
rect 263597 9333 263609 9367
rect 263643 9364 263655 9367
rect 264146 9364 264152 9376
rect 263643 9336 264152 9364
rect 263643 9333 263655 9336
rect 263597 9327 263655 9333
rect 264146 9324 264152 9336
rect 264204 9324 264210 9376
rect 265526 9324 265532 9376
rect 265584 9364 265590 9376
rect 266280 9364 266308 9404
rect 268746 9392 268752 9404
rect 268804 9392 268810 9444
rect 268933 9435 268991 9441
rect 268933 9401 268945 9435
rect 268979 9432 268991 9435
rect 270586 9432 270592 9444
rect 268979 9404 270592 9432
rect 268979 9401 268991 9404
rect 268933 9395 268991 9401
rect 270586 9392 270592 9404
rect 270644 9392 270650 9444
rect 265584 9336 266308 9364
rect 265584 9324 265590 9336
rect 266354 9324 266360 9376
rect 266412 9364 266418 9376
rect 267277 9367 267335 9373
rect 267277 9364 267289 9367
rect 266412 9336 267289 9364
rect 266412 9324 266418 9336
rect 267277 9333 267289 9336
rect 267323 9333 267335 9367
rect 267277 9327 267335 9333
rect 269206 9324 269212 9376
rect 269264 9324 269270 9376
rect 269666 9324 269672 9376
rect 269724 9324 269730 9376
rect 1104 9274 271492 9296
rect 1104 9222 34748 9274
rect 34800 9222 34812 9274
rect 34864 9222 34876 9274
rect 34928 9222 34940 9274
rect 34992 9222 35004 9274
rect 35056 9222 102345 9274
rect 102397 9222 102409 9274
rect 102461 9222 102473 9274
rect 102525 9222 102537 9274
rect 102589 9222 102601 9274
rect 102653 9222 169942 9274
rect 169994 9222 170006 9274
rect 170058 9222 170070 9274
rect 170122 9222 170134 9274
rect 170186 9222 170198 9274
rect 170250 9222 237539 9274
rect 237591 9222 237603 9274
rect 237655 9222 237667 9274
rect 237719 9222 237731 9274
rect 237783 9222 237795 9274
rect 237847 9222 271492 9274
rect 1104 9200 271492 9222
rect 1394 9120 1400 9172
rect 1452 9160 1458 9172
rect 1765 9163 1823 9169
rect 1765 9160 1777 9163
rect 1452 9132 1777 9160
rect 1452 9120 1458 9132
rect 1765 9129 1777 9132
rect 1811 9129 1823 9163
rect 1765 9123 1823 9129
rect 3234 9120 3240 9172
rect 3292 9160 3298 9172
rect 3292 9132 23796 9160
rect 3292 9120 3298 9132
rect 7650 9052 7656 9104
rect 7708 9092 7714 9104
rect 7708 9064 23704 9092
rect 7708 9052 7714 9064
rect 5166 8984 5172 9036
rect 5224 9024 5230 9036
rect 17218 9024 17224 9036
rect 5224 8996 17224 9024
rect 5224 8984 5230 8996
rect 17218 8984 17224 8996
rect 17276 8984 17282 9036
rect 21726 9024 21732 9036
rect 20456 8996 21732 9024
rect 3142 8916 3148 8968
rect 3200 8916 3206 8968
rect 8202 8916 8208 8968
rect 8260 8956 8266 8968
rect 8297 8959 8355 8965
rect 8297 8956 8309 8959
rect 8260 8928 8309 8956
rect 8260 8916 8266 8928
rect 8297 8925 8309 8928
rect 8343 8925 8355 8959
rect 8297 8919 8355 8925
rect 13446 8916 13452 8968
rect 13504 8916 13510 8968
rect 14734 8916 14740 8968
rect 14792 8956 14798 8968
rect 18414 8956 18420 8968
rect 14792 8928 18420 8956
rect 14792 8916 14798 8928
rect 18414 8916 18420 8928
rect 18472 8916 18478 8968
rect 20254 8916 20260 8968
rect 20312 8916 20318 8968
rect 3326 8848 3332 8900
rect 3384 8848 3390 8900
rect 8478 8848 8484 8900
rect 8536 8848 8542 8900
rect 13630 8848 13636 8900
rect 13688 8848 13694 8900
rect 7558 8780 7564 8832
rect 7616 8820 7622 8832
rect 19334 8820 19340 8832
rect 7616 8792 19340 8820
rect 7616 8780 7622 8792
rect 19334 8780 19340 8792
rect 19392 8780 19398 8832
rect 20456 8829 20484 8996
rect 21726 8984 21732 8996
rect 21784 8984 21790 9036
rect 23198 8984 23204 9036
rect 23256 8984 23262 9036
rect 20901 8959 20959 8965
rect 20901 8925 20913 8959
rect 20947 8956 20959 8959
rect 21082 8956 21088 8968
rect 20947 8928 21088 8956
rect 20947 8925 20959 8928
rect 20901 8919 20959 8925
rect 21082 8916 21088 8928
rect 21140 8916 21146 8968
rect 21177 8959 21235 8965
rect 21177 8925 21189 8959
rect 21223 8956 21235 8959
rect 21450 8956 21456 8968
rect 21223 8928 21456 8956
rect 21223 8925 21235 8928
rect 21177 8919 21235 8925
rect 21450 8916 21456 8928
rect 21508 8916 21514 8968
rect 21634 8916 21640 8968
rect 21692 8956 21698 8968
rect 22097 8959 22155 8965
rect 22097 8958 22109 8959
rect 21928 8956 22109 8958
rect 21692 8930 22109 8956
rect 21692 8928 21956 8930
rect 21692 8916 21698 8928
rect 20441 8823 20499 8829
rect 20441 8789 20453 8823
rect 20487 8789 20499 8823
rect 20441 8783 20499 8789
rect 21361 8823 21419 8829
rect 21361 8789 21373 8823
rect 21407 8820 21419 8823
rect 21634 8820 21640 8832
rect 21407 8792 21640 8820
rect 21407 8789 21419 8792
rect 21361 8783 21419 8789
rect 21634 8780 21640 8792
rect 21692 8780 21698 8832
rect 21928 8820 21956 8928
rect 22097 8925 22109 8930
rect 22143 8925 22155 8959
rect 22097 8919 22155 8925
rect 22186 8916 22192 8968
rect 22244 8916 22250 8968
rect 22922 8916 22928 8968
rect 22980 8916 22986 8968
rect 23676 8888 23704 9064
rect 23768 9024 23796 9132
rect 23934 9120 23940 9172
rect 23992 9120 23998 9172
rect 30374 9120 30380 9172
rect 30432 9120 30438 9172
rect 32122 9120 32128 9172
rect 32180 9120 32186 9172
rect 33042 9120 33048 9172
rect 33100 9120 33106 9172
rect 35158 9120 35164 9172
rect 35216 9120 35222 9172
rect 53282 9120 53288 9172
rect 53340 9120 53346 9172
rect 53834 9120 53840 9172
rect 53892 9120 53898 9172
rect 54938 9120 54944 9172
rect 54996 9120 55002 9172
rect 55674 9120 55680 9172
rect 55732 9120 55738 9172
rect 56594 9120 56600 9172
rect 56652 9120 56658 9172
rect 57241 9163 57299 9169
rect 57241 9129 57253 9163
rect 57287 9160 57299 9163
rect 58066 9160 58072 9172
rect 57287 9132 58072 9160
rect 57287 9129 57299 9132
rect 57241 9123 57299 9129
rect 58066 9120 58072 9132
rect 58124 9120 58130 9172
rect 58526 9120 58532 9172
rect 58584 9120 58590 9172
rect 62206 9120 62212 9172
rect 62264 9120 62270 9172
rect 62758 9120 62764 9172
rect 62816 9120 62822 9172
rect 64046 9120 64052 9172
rect 64104 9160 64110 9172
rect 64104 9132 73660 9160
rect 64104 9120 64110 9132
rect 24026 9052 24032 9104
rect 24084 9092 24090 9104
rect 41506 9092 41512 9104
rect 24084 9064 41512 9092
rect 24084 9052 24090 9064
rect 41506 9052 41512 9064
rect 41564 9052 41570 9104
rect 46198 9052 46204 9104
rect 46256 9092 46262 9104
rect 57974 9092 57980 9104
rect 46256 9064 57980 9092
rect 46256 9052 46262 9064
rect 57974 9052 57980 9064
rect 58032 9052 58038 9104
rect 62298 9052 62304 9104
rect 62356 9092 62362 9104
rect 73632 9092 73660 9132
rect 73706 9120 73712 9172
rect 73764 9160 73770 9172
rect 84838 9160 84844 9172
rect 73764 9132 84844 9160
rect 73764 9120 73770 9132
rect 84838 9120 84844 9132
rect 84896 9120 84902 9172
rect 88242 9120 88248 9172
rect 88300 9160 88306 9172
rect 88429 9163 88487 9169
rect 88429 9160 88441 9163
rect 88300 9132 88441 9160
rect 88300 9120 88306 9132
rect 88429 9129 88441 9132
rect 88475 9129 88487 9163
rect 88429 9123 88487 9129
rect 90082 9120 90088 9172
rect 90140 9160 90146 9172
rect 90177 9163 90235 9169
rect 90177 9160 90189 9163
rect 90140 9132 90189 9160
rect 90140 9120 90146 9132
rect 90177 9129 90189 9132
rect 90223 9129 90235 9163
rect 90177 9123 90235 9129
rect 90542 9120 90548 9172
rect 90600 9160 90606 9172
rect 91646 9160 91652 9172
rect 90600 9132 91652 9160
rect 90600 9120 90606 9132
rect 91646 9120 91652 9132
rect 91704 9120 91710 9172
rect 91738 9120 91744 9172
rect 91796 9120 91802 9172
rect 93670 9120 93676 9172
rect 93728 9120 93734 9172
rect 94222 9160 94228 9172
rect 93964 9132 94228 9160
rect 81066 9092 81072 9104
rect 62356 9064 73568 9092
rect 73632 9064 81072 9092
rect 62356 9052 62362 9064
rect 25501 9027 25559 9033
rect 23768 8996 24164 9024
rect 23753 8959 23811 8965
rect 23753 8925 23765 8959
rect 23799 8956 23811 8959
rect 24026 8956 24032 8968
rect 23799 8928 24032 8956
rect 23799 8925 23811 8928
rect 23753 8919 23811 8925
rect 24026 8916 24032 8928
rect 24084 8916 24090 8968
rect 23934 8888 23940 8900
rect 23676 8860 23940 8888
rect 23934 8848 23940 8860
rect 23992 8848 23998 8900
rect 24136 8888 24164 8996
rect 25501 8993 25513 9027
rect 25547 9024 25559 9027
rect 31481 9027 31539 9033
rect 25547 8996 30972 9024
rect 25547 8993 25559 8996
rect 25501 8987 25559 8993
rect 27172 8968 27200 8996
rect 24670 8916 24676 8968
rect 24728 8916 24734 8968
rect 25682 8916 25688 8968
rect 25740 8956 25746 8968
rect 25777 8959 25835 8965
rect 25777 8956 25789 8959
rect 25740 8928 25789 8956
rect 25740 8916 25746 8928
rect 25777 8925 25789 8928
rect 25823 8925 25835 8959
rect 25777 8919 25835 8925
rect 26697 8959 26755 8965
rect 26697 8925 26709 8959
rect 26743 8956 26755 8959
rect 27062 8956 27068 8968
rect 26743 8928 27068 8956
rect 26743 8925 26755 8928
rect 26697 8919 26755 8925
rect 27062 8916 27068 8928
rect 27120 8916 27126 8968
rect 27154 8916 27160 8968
rect 27212 8916 27218 8968
rect 27706 8916 27712 8968
rect 27764 8956 27770 8968
rect 28000 8965 28028 8996
rect 27801 8959 27859 8965
rect 27801 8956 27813 8959
rect 27764 8928 27813 8956
rect 27764 8916 27770 8928
rect 27801 8925 27813 8928
rect 27847 8925 27859 8959
rect 27801 8919 27859 8925
rect 27985 8959 28043 8965
rect 27985 8925 27997 8959
rect 28031 8925 28043 8959
rect 27985 8919 28043 8925
rect 28534 8916 28540 8968
rect 28592 8956 28598 8968
rect 28828 8965 28856 8996
rect 28629 8959 28687 8965
rect 28629 8956 28641 8959
rect 28592 8928 28641 8956
rect 28592 8916 28598 8928
rect 28629 8925 28641 8928
rect 28675 8925 28687 8959
rect 28629 8919 28687 8925
rect 28813 8959 28871 8965
rect 28813 8925 28825 8959
rect 28859 8925 28871 8959
rect 28813 8919 28871 8925
rect 30098 8916 30104 8968
rect 30156 8916 30162 8968
rect 30208 8965 30236 8996
rect 30193 8959 30251 8965
rect 30193 8925 30205 8959
rect 30239 8925 30251 8959
rect 30193 8919 30251 8925
rect 30742 8916 30748 8968
rect 30800 8916 30806 8968
rect 30944 8965 30972 8996
rect 31481 8993 31493 9027
rect 31527 9024 31539 9027
rect 31757 9027 31815 9033
rect 31757 9024 31769 9027
rect 31527 8996 31769 9024
rect 31527 8993 31539 8996
rect 31481 8987 31539 8993
rect 31757 8993 31769 8996
rect 31803 9024 31815 9027
rect 31846 9024 31852 9036
rect 31803 8996 31852 9024
rect 31803 8993 31815 8996
rect 31757 8987 31815 8993
rect 31846 8984 31852 8996
rect 31904 9024 31910 9036
rect 32766 9024 32772 9036
rect 31904 8996 32772 9024
rect 31904 8984 31910 8996
rect 32766 8984 32772 8996
rect 32824 8984 32830 9036
rect 32950 8984 32956 9036
rect 33008 9024 33014 9036
rect 55674 9024 55680 9036
rect 33008 8996 41414 9024
rect 33008 8984 33014 8996
rect 30929 8959 30987 8965
rect 30929 8925 30941 8959
rect 30975 8956 30987 8959
rect 31938 8956 31944 8968
rect 30975 8928 31944 8956
rect 30975 8925 30987 8928
rect 30929 8919 30987 8925
rect 31938 8916 31944 8928
rect 31996 8916 32002 8968
rect 32861 8959 32919 8965
rect 32861 8925 32873 8959
rect 32907 8956 32919 8959
rect 33134 8956 33140 8968
rect 32907 8928 33140 8956
rect 32907 8925 32919 8928
rect 32861 8919 32919 8925
rect 33134 8916 33140 8928
rect 33192 8916 33198 8968
rect 40310 8916 40316 8968
rect 40368 8916 40374 8968
rect 36446 8888 36452 8900
rect 24136 8860 36452 8888
rect 36446 8848 36452 8860
rect 36504 8848 36510 8900
rect 39666 8888 39672 8900
rect 36556 8860 39672 8888
rect 22094 8820 22100 8832
rect 21928 8792 22100 8820
rect 22094 8780 22100 8792
rect 22152 8780 22158 8832
rect 22373 8823 22431 8829
rect 22373 8789 22385 8823
rect 22419 8820 22431 8823
rect 22738 8820 22744 8832
rect 22419 8792 22744 8820
rect 22419 8789 22431 8792
rect 22373 8783 22431 8789
rect 22738 8780 22744 8792
rect 22796 8780 22802 8832
rect 24762 8780 24768 8832
rect 24820 8780 24826 8832
rect 27246 8780 27252 8832
rect 27304 8820 27310 8832
rect 27341 8823 27399 8829
rect 27341 8820 27353 8823
rect 27304 8792 27353 8820
rect 27304 8780 27310 8792
rect 27341 8789 27353 8792
rect 27387 8789 27399 8823
rect 27341 8783 27399 8789
rect 27982 8780 27988 8832
rect 28040 8820 28046 8832
rect 28169 8823 28227 8829
rect 28169 8820 28181 8823
rect 28040 8792 28181 8820
rect 28040 8780 28046 8792
rect 28169 8789 28181 8792
rect 28215 8789 28227 8823
rect 28169 8783 28227 8789
rect 28718 8780 28724 8832
rect 28776 8820 28782 8832
rect 28997 8823 29055 8829
rect 28997 8820 29009 8823
rect 28776 8792 29009 8820
rect 28776 8780 28782 8792
rect 28997 8789 29009 8792
rect 29043 8789 29055 8823
rect 28997 8783 29055 8789
rect 30834 8780 30840 8832
rect 30892 8820 30898 8832
rect 31113 8823 31171 8829
rect 31113 8820 31125 8823
rect 30892 8792 31125 8820
rect 30892 8780 30898 8792
rect 31113 8789 31125 8792
rect 31159 8789 31171 8823
rect 31113 8783 31171 8789
rect 32766 8780 32772 8832
rect 32824 8820 32830 8832
rect 36556 8820 36584 8860
rect 39666 8848 39672 8860
rect 39724 8848 39730 8900
rect 41386 8888 41414 8996
rect 54772 8996 55680 9024
rect 45462 8916 45468 8968
rect 45520 8916 45526 8968
rect 53098 8916 53104 8968
rect 53156 8916 53162 8968
rect 53650 8916 53656 8968
rect 53708 8916 53714 8968
rect 54110 8916 54116 8968
rect 54168 8956 54174 8968
rect 54573 8959 54631 8965
rect 54573 8956 54585 8959
rect 54168 8928 54585 8956
rect 54168 8916 54174 8928
rect 54573 8925 54585 8928
rect 54619 8925 54631 8959
rect 54573 8919 54631 8925
rect 54662 8916 54668 8968
rect 54720 8956 54726 8968
rect 54772 8965 54800 8996
rect 55674 8984 55680 8996
rect 55732 9024 55738 9036
rect 57146 9024 57152 9036
rect 55732 8996 57152 9024
rect 55732 8984 55738 8996
rect 54757 8959 54815 8965
rect 54757 8956 54769 8959
rect 54720 8928 54769 8956
rect 54720 8916 54726 8928
rect 54757 8925 54769 8928
rect 54803 8925 54815 8959
rect 54757 8919 54815 8925
rect 55493 8959 55551 8965
rect 55493 8925 55505 8959
rect 55539 8956 55551 8959
rect 55858 8956 55864 8968
rect 55539 8928 55864 8956
rect 55539 8925 55551 8928
rect 55493 8919 55551 8925
rect 55858 8916 55864 8928
rect 55916 8916 55922 8968
rect 56318 8916 56324 8968
rect 56376 8916 56382 8968
rect 56428 8965 56456 8996
rect 56413 8959 56471 8965
rect 56413 8925 56425 8959
rect 56459 8925 56471 8959
rect 56413 8919 56471 8925
rect 56870 8916 56876 8968
rect 56928 8916 56934 8968
rect 57072 8965 57100 8996
rect 57146 8984 57152 8996
rect 57204 9024 57210 9036
rect 57204 8996 59952 9024
rect 57204 8984 57210 8996
rect 57057 8959 57115 8965
rect 57057 8925 57069 8959
rect 57103 8925 57115 8959
rect 57057 8919 57115 8925
rect 57609 8959 57667 8965
rect 57609 8925 57621 8959
rect 57655 8956 57667 8959
rect 57885 8959 57943 8965
rect 57885 8956 57897 8959
rect 57655 8928 57897 8956
rect 57655 8925 57667 8928
rect 57609 8919 57667 8925
rect 57885 8925 57897 8928
rect 57931 8956 57943 8959
rect 57974 8956 57980 8968
rect 57931 8928 57980 8956
rect 57931 8925 57943 8928
rect 57885 8919 57943 8925
rect 57974 8916 57980 8928
rect 58032 8916 58038 8968
rect 58084 8965 58112 8996
rect 58069 8959 58127 8965
rect 58069 8925 58081 8959
rect 58115 8925 58127 8959
rect 58069 8919 58127 8925
rect 58526 8916 58532 8968
rect 58584 8956 58590 8968
rect 59096 8965 59124 8996
rect 59924 8968 59952 8996
rect 60642 8984 60648 9036
rect 60700 8984 60706 9036
rect 65978 9024 65984 9036
rect 60844 8996 65984 9024
rect 58897 8959 58955 8965
rect 58897 8956 58909 8959
rect 58584 8928 58909 8956
rect 58584 8916 58590 8928
rect 58897 8925 58909 8928
rect 58943 8925 58955 8959
rect 58897 8919 58955 8925
rect 59081 8959 59139 8965
rect 59081 8925 59093 8959
rect 59127 8925 59139 8959
rect 59081 8919 59139 8925
rect 59722 8916 59728 8968
rect 59780 8916 59786 8968
rect 59906 8916 59912 8968
rect 59964 8916 59970 8968
rect 60844 8965 60872 8996
rect 60829 8959 60887 8965
rect 60829 8925 60841 8959
rect 60875 8925 60887 8959
rect 60829 8919 60887 8925
rect 61470 8916 61476 8968
rect 61528 8956 61534 8968
rect 62040 8965 62068 8996
rect 61841 8959 61899 8965
rect 61841 8956 61853 8959
rect 61528 8928 61853 8956
rect 61528 8916 61534 8928
rect 61841 8925 61853 8928
rect 61887 8925 61899 8959
rect 61841 8919 61899 8925
rect 62025 8959 62083 8965
rect 62025 8925 62037 8959
rect 62071 8925 62083 8959
rect 62025 8919 62083 8925
rect 62393 8959 62451 8965
rect 62393 8925 62405 8959
rect 62439 8925 62451 8959
rect 62393 8919 62451 8925
rect 62298 8888 62304 8900
rect 41386 8860 62304 8888
rect 62298 8848 62304 8860
rect 62356 8888 62362 8900
rect 62408 8888 62436 8919
rect 62482 8916 62488 8968
rect 62540 8956 62546 8968
rect 62592 8965 62620 8996
rect 62577 8959 62635 8965
rect 62577 8956 62589 8959
rect 62540 8928 62589 8956
rect 62540 8916 62546 8928
rect 62577 8925 62589 8928
rect 62623 8925 62635 8959
rect 62577 8919 62635 8925
rect 63218 8916 63224 8968
rect 63276 8916 63282 8968
rect 63420 8965 63448 8996
rect 63405 8959 63463 8965
rect 63405 8925 63417 8959
rect 63451 8925 63463 8959
rect 63405 8919 63463 8925
rect 64046 8916 64052 8968
rect 64104 8916 64110 8968
rect 64248 8965 64276 8996
rect 64233 8959 64291 8965
rect 64233 8925 64245 8959
rect 64279 8925 64291 8959
rect 64233 8919 64291 8925
rect 64966 8916 64972 8968
rect 65024 8916 65030 8968
rect 65076 8965 65104 8996
rect 65978 8984 65984 8996
rect 66036 9024 66042 9036
rect 66809 9027 66867 9033
rect 66036 8996 66208 9024
rect 66036 8984 66042 8996
rect 65061 8959 65119 8965
rect 65061 8925 65073 8959
rect 65107 8925 65119 8959
rect 65061 8919 65119 8925
rect 66070 8916 66076 8968
rect 66128 8916 66134 8968
rect 66180 8966 66208 8996
rect 66809 8993 66821 9027
rect 66855 9024 66867 9027
rect 70394 9024 70400 9036
rect 66855 8996 70400 9024
rect 66855 8993 66867 8996
rect 66809 8987 66867 8993
rect 66243 8969 66301 8975
rect 66243 8966 66255 8969
rect 66180 8938 66255 8966
rect 66243 8935 66255 8938
rect 66289 8935 66301 8969
rect 66243 8929 66301 8935
rect 66346 8916 66352 8968
rect 66404 8952 66410 8968
rect 66824 8956 66852 8987
rect 70394 8984 70400 8996
rect 70452 8984 70458 9036
rect 72050 8984 72056 9036
rect 72108 8984 72114 9036
rect 73430 8984 73436 9036
rect 73488 8984 73494 9036
rect 73540 9024 73568 9064
rect 81066 9052 81072 9064
rect 81124 9052 81130 9104
rect 93964 9092 93992 9132
rect 94222 9120 94228 9132
rect 94280 9160 94286 9172
rect 96062 9160 96068 9172
rect 94280 9132 96068 9160
rect 94280 9120 94286 9132
rect 96062 9120 96068 9132
rect 96120 9120 96126 9172
rect 96246 9120 96252 9172
rect 96304 9160 96310 9172
rect 96522 9160 96528 9172
rect 96304 9132 96528 9160
rect 96304 9120 96310 9132
rect 96522 9120 96528 9132
rect 96580 9160 96586 9172
rect 97718 9160 97724 9172
rect 96580 9132 97724 9160
rect 96580 9120 96586 9132
rect 97718 9120 97724 9132
rect 97776 9120 97782 9172
rect 98914 9120 98920 9172
rect 98972 9120 98978 9172
rect 100570 9120 100576 9172
rect 100628 9120 100634 9172
rect 101214 9120 101220 9172
rect 101272 9120 101278 9172
rect 107010 9120 107016 9172
rect 107068 9120 107074 9172
rect 111886 9120 111892 9172
rect 111944 9160 111950 9172
rect 115014 9160 115020 9172
rect 111944 9132 115020 9160
rect 111944 9120 111950 9132
rect 115014 9120 115020 9132
rect 115072 9120 115078 9172
rect 120994 9120 121000 9172
rect 121052 9160 121058 9172
rect 121052 9132 121960 9160
rect 121052 9120 121058 9132
rect 81176 9064 93992 9092
rect 81176 9024 81204 9064
rect 94038 9052 94044 9104
rect 94096 9092 94102 9104
rect 103698 9092 103704 9104
rect 94096 9064 103704 9092
rect 94096 9052 94102 9064
rect 103698 9052 103704 9064
rect 103756 9052 103762 9104
rect 104986 9052 104992 9104
rect 105044 9092 105050 9104
rect 108942 9092 108948 9104
rect 105044 9064 108948 9092
rect 105044 9052 105050 9064
rect 108942 9052 108948 9064
rect 109000 9052 109006 9104
rect 111150 9052 111156 9104
rect 111208 9092 111214 9104
rect 115750 9092 115756 9104
rect 111208 9064 115756 9092
rect 111208 9052 111214 9064
rect 115750 9052 115756 9064
rect 115808 9052 115814 9104
rect 121089 9095 121147 9101
rect 121089 9061 121101 9095
rect 121135 9092 121147 9095
rect 121822 9092 121828 9104
rect 121135 9064 121828 9092
rect 121135 9061 121147 9064
rect 121089 9055 121147 9061
rect 121822 9052 121828 9064
rect 121880 9052 121886 9104
rect 121932 9092 121960 9132
rect 124398 9120 124404 9172
rect 124456 9120 124462 9172
rect 124674 9120 124680 9172
rect 124732 9120 124738 9172
rect 126238 9120 126244 9172
rect 126296 9120 126302 9172
rect 127618 9120 127624 9172
rect 127676 9160 127682 9172
rect 128722 9160 128728 9172
rect 127676 9132 128728 9160
rect 127676 9120 127682 9132
rect 128722 9120 128728 9132
rect 128780 9120 128786 9172
rect 130562 9120 130568 9172
rect 130620 9120 130626 9172
rect 131390 9120 131396 9172
rect 131448 9120 131454 9172
rect 133046 9120 133052 9172
rect 133104 9120 133110 9172
rect 134058 9120 134064 9172
rect 134116 9120 134122 9172
rect 134702 9120 134708 9172
rect 134760 9120 134766 9172
rect 142798 9120 142804 9172
rect 142856 9160 142862 9172
rect 148594 9160 148600 9172
rect 142856 9132 148600 9160
rect 142856 9120 142862 9132
rect 148594 9120 148600 9132
rect 148652 9120 148658 9172
rect 152458 9120 152464 9172
rect 152516 9160 152522 9172
rect 175550 9160 175556 9172
rect 152516 9132 175556 9160
rect 152516 9120 152522 9132
rect 175550 9120 175556 9132
rect 175608 9120 175614 9172
rect 176838 9120 176844 9172
rect 176896 9120 176902 9172
rect 177574 9120 177580 9172
rect 177632 9120 177638 9172
rect 184566 9160 184572 9172
rect 180766 9132 184572 9160
rect 133874 9092 133880 9104
rect 121932 9064 128584 9092
rect 73540 8996 81204 9024
rect 81250 8984 81256 9036
rect 81308 8984 81314 9036
rect 81526 8984 81532 9036
rect 81584 8984 81590 9036
rect 81820 8996 82768 9024
rect 66456 8952 66852 8956
rect 66404 8928 66852 8952
rect 66404 8924 66484 8928
rect 66404 8916 66410 8924
rect 66990 8916 66996 8968
rect 67048 8916 67054 8968
rect 70026 8916 70032 8968
rect 70084 8916 70090 8968
rect 72326 8916 72332 8968
rect 72384 8916 72390 8968
rect 73706 8916 73712 8968
rect 73764 8916 73770 8968
rect 74718 8916 74724 8968
rect 74776 8916 74782 8968
rect 74994 8916 75000 8968
rect 75052 8916 75058 8968
rect 77202 8916 77208 8968
rect 77260 8916 77266 8968
rect 77478 8916 77484 8968
rect 77536 8916 77542 8968
rect 78674 8916 78680 8968
rect 78732 8916 78738 8968
rect 78950 8916 78956 8968
rect 79008 8916 79014 8968
rect 62356 8860 62436 8888
rect 62356 8848 62362 8860
rect 62666 8848 62672 8900
rect 62724 8888 62730 8900
rect 81820 8888 81848 8996
rect 82630 8916 82636 8968
rect 82688 8916 82694 8968
rect 82740 8956 82768 8996
rect 82814 8984 82820 9036
rect 82872 8984 82878 9036
rect 86402 8984 86408 9036
rect 86460 8984 86466 9036
rect 89530 9024 89536 9036
rect 86512 8996 89536 9024
rect 86512 8956 86540 8996
rect 89530 8984 89536 8996
rect 89588 8984 89594 9036
rect 89640 8996 94360 9024
rect 82740 8928 86540 8956
rect 86678 8916 86684 8968
rect 86736 8916 86742 8968
rect 88245 8959 88303 8965
rect 88245 8925 88257 8959
rect 88291 8925 88303 8959
rect 88245 8919 88303 8925
rect 88260 8888 88288 8919
rect 89070 8916 89076 8968
rect 89128 8916 89134 8968
rect 89165 8959 89223 8965
rect 89165 8925 89177 8959
rect 89211 8956 89223 8959
rect 89438 8956 89444 8968
rect 89211 8928 89444 8956
rect 89211 8925 89223 8928
rect 89165 8919 89223 8925
rect 89438 8916 89444 8928
rect 89496 8956 89502 8968
rect 89640 8956 89668 8996
rect 90008 8968 90036 8996
rect 89496 8928 89668 8956
rect 89496 8916 89502 8928
rect 89898 8916 89904 8968
rect 89956 8916 89962 8968
rect 89990 8916 89996 8968
rect 90048 8916 90054 8968
rect 90726 8916 90732 8968
rect 90784 8916 90790 8968
rect 90836 8965 90864 8996
rect 90821 8959 90879 8965
rect 90821 8925 90833 8959
rect 90867 8925 90879 8959
rect 90821 8919 90879 8925
rect 91557 8959 91615 8965
rect 91557 8925 91569 8959
rect 91603 8925 91615 8959
rect 91557 8919 91615 8925
rect 89349 8891 89407 8897
rect 89349 8888 89361 8891
rect 62724 8860 81848 8888
rect 81912 8860 82860 8888
rect 88260 8860 89361 8888
rect 62724 8848 62730 8860
rect 32824 8792 36584 8820
rect 32824 8780 32830 8792
rect 39390 8780 39396 8832
rect 39448 8820 39454 8832
rect 40129 8823 40187 8829
rect 40129 8820 40141 8823
rect 39448 8792 40141 8820
rect 39448 8780 39454 8792
rect 40129 8789 40141 8792
rect 40175 8789 40187 8823
rect 40129 8783 40187 8789
rect 44726 8780 44732 8832
rect 44784 8820 44790 8832
rect 45281 8823 45339 8829
rect 45281 8820 45293 8823
rect 44784 8792 45293 8820
rect 44784 8780 44790 8792
rect 45281 8789 45293 8792
rect 45327 8789 45339 8823
rect 45281 8783 45339 8789
rect 54110 8780 54116 8832
rect 54168 8820 54174 8832
rect 54205 8823 54263 8829
rect 54205 8820 54217 8823
rect 54168 8792 54217 8820
rect 54168 8780 54174 8792
rect 54205 8789 54217 8792
rect 54251 8789 54263 8823
rect 54205 8783 54263 8789
rect 56870 8780 56876 8832
rect 56928 8820 56934 8832
rect 57422 8820 57428 8832
rect 56928 8792 57428 8820
rect 56928 8780 56934 8792
rect 57422 8780 57428 8792
rect 57480 8780 57486 8832
rect 58250 8780 58256 8832
rect 58308 8780 58314 8832
rect 59265 8823 59323 8829
rect 59265 8789 59277 8823
rect 59311 8820 59323 8823
rect 59354 8820 59360 8832
rect 59311 8792 59360 8820
rect 59311 8789 59323 8792
rect 59265 8783 59323 8789
rect 59354 8780 59360 8792
rect 59412 8780 59418 8832
rect 60090 8780 60096 8832
rect 60148 8780 60154 8832
rect 60826 8780 60832 8832
rect 60884 8820 60890 8832
rect 61013 8823 61071 8829
rect 61013 8820 61025 8823
rect 60884 8792 61025 8820
rect 60884 8780 60890 8792
rect 61013 8789 61025 8792
rect 61059 8789 61071 8823
rect 61013 8783 61071 8789
rect 61470 8780 61476 8832
rect 61528 8780 61534 8832
rect 63589 8823 63647 8829
rect 63589 8789 63601 8823
rect 63635 8820 63647 8823
rect 63770 8820 63776 8832
rect 63635 8792 63776 8820
rect 63635 8789 63647 8792
rect 63589 8783 63647 8789
rect 63770 8780 63776 8792
rect 63828 8780 63834 8832
rect 64417 8823 64475 8829
rect 64417 8789 64429 8823
rect 64463 8820 64475 8823
rect 64506 8820 64512 8832
rect 64463 8792 64512 8820
rect 64463 8789 64475 8792
rect 64417 8783 64475 8789
rect 64506 8780 64512 8792
rect 64564 8780 64570 8832
rect 65245 8823 65303 8829
rect 65245 8789 65257 8823
rect 65291 8820 65303 8823
rect 65334 8820 65340 8832
rect 65291 8792 65340 8820
rect 65291 8789 65303 8792
rect 65245 8783 65303 8789
rect 65334 8780 65340 8792
rect 65392 8780 65398 8832
rect 66070 8780 66076 8832
rect 66128 8820 66134 8832
rect 66441 8823 66499 8829
rect 66441 8820 66453 8823
rect 66128 8792 66453 8820
rect 66128 8780 66134 8792
rect 66441 8789 66453 8792
rect 66487 8789 66499 8823
rect 66441 8783 66499 8789
rect 67174 8780 67180 8832
rect 67232 8780 67238 8832
rect 69845 8823 69903 8829
rect 69845 8789 69857 8823
rect 69891 8820 69903 8823
rect 81912 8820 81940 8860
rect 69891 8792 81940 8820
rect 82832 8820 82860 8860
rect 89349 8857 89361 8860
rect 89395 8857 89407 8891
rect 91094 8888 91100 8900
rect 89349 8851 89407 8857
rect 89456 8860 91100 8888
rect 89456 8820 89484 8860
rect 91094 8848 91100 8860
rect 91152 8848 91158 8900
rect 91572 8888 91600 8919
rect 91646 8916 91652 8968
rect 91704 8956 91710 8968
rect 92382 8956 92388 8968
rect 91704 8928 92388 8956
rect 91704 8916 91710 8928
rect 92382 8916 92388 8928
rect 92440 8916 92446 8968
rect 92492 8965 92520 8996
rect 93504 8968 93532 8996
rect 92477 8959 92535 8965
rect 92477 8925 92489 8959
rect 92523 8925 92535 8959
rect 92477 8919 92535 8925
rect 92842 8916 92848 8968
rect 92900 8956 92906 8968
rect 93029 8959 93087 8965
rect 93029 8956 93041 8959
rect 92900 8928 93041 8956
rect 92900 8916 92906 8928
rect 93029 8925 93041 8928
rect 93075 8956 93087 8959
rect 93394 8956 93400 8968
rect 93075 8928 93400 8956
rect 93075 8925 93087 8928
rect 93029 8919 93087 8925
rect 93394 8916 93400 8928
rect 93452 8916 93458 8968
rect 93486 8916 93492 8968
rect 93544 8916 93550 8968
rect 94332 8965 94360 8996
rect 94590 8984 94596 9036
rect 94648 9024 94654 9036
rect 94961 9027 95019 9033
rect 94961 9024 94973 9027
rect 94648 8996 94973 9024
rect 94648 8984 94654 8996
rect 94961 8993 94973 8996
rect 95007 8993 95019 9027
rect 95234 9024 95240 9036
rect 94961 8987 95019 8993
rect 95160 8996 95240 9024
rect 94133 8959 94191 8965
rect 94133 8925 94145 8959
rect 94179 8925 94191 8959
rect 94133 8919 94191 8925
rect 94317 8959 94375 8965
rect 94317 8925 94329 8959
rect 94363 8956 94375 8959
rect 94866 8956 94872 8968
rect 94363 8928 94872 8956
rect 94363 8925 94375 8928
rect 94317 8919 94375 8925
rect 92661 8891 92719 8897
rect 92661 8888 92673 8891
rect 91572 8860 92673 8888
rect 92661 8857 92673 8860
rect 92707 8857 92719 8891
rect 92661 8851 92719 8857
rect 92934 8848 92940 8900
rect 92992 8888 92998 8900
rect 93118 8888 93124 8900
rect 92992 8860 93124 8888
rect 92992 8848 92998 8860
rect 93118 8848 93124 8860
rect 93176 8888 93182 8900
rect 94148 8888 94176 8919
rect 94866 8916 94872 8928
rect 94924 8916 94930 8968
rect 95160 8965 95188 8996
rect 95234 8984 95240 8996
rect 95292 8984 95298 9036
rect 95970 8984 95976 9036
rect 96028 8984 96034 9036
rect 96522 8984 96528 9036
rect 96580 9024 96586 9036
rect 99190 9024 99196 9036
rect 96580 8996 99196 9024
rect 96580 8984 96586 8996
rect 99190 8984 99196 8996
rect 99248 8984 99254 9036
rect 99282 8984 99288 9036
rect 99340 9024 99346 9036
rect 123294 9024 123300 9036
rect 99340 8996 123300 9024
rect 99340 8984 99346 8996
rect 123294 8984 123300 8996
rect 123352 8984 123358 9036
rect 123389 9027 123447 9033
rect 123389 8993 123401 9027
rect 123435 9024 123447 9027
rect 123478 9024 123484 9036
rect 123435 8996 123484 9024
rect 123435 8993 123447 8996
rect 123389 8987 123447 8993
rect 123478 8984 123484 8996
rect 123536 8984 123542 9036
rect 128556 9033 128584 9064
rect 128648 9064 133880 9092
rect 128541 9027 128599 9033
rect 123588 8996 127848 9024
rect 95145 8959 95203 8965
rect 95145 8925 95157 8959
rect 95191 8925 95203 8959
rect 96614 8956 96620 8968
rect 95145 8919 95203 8925
rect 95620 8928 96620 8956
rect 95620 8897 95648 8928
rect 96614 8916 96620 8928
rect 96672 8916 96678 8968
rect 96982 8916 96988 8968
rect 97040 8916 97046 8968
rect 97077 8959 97135 8965
rect 97077 8925 97089 8959
rect 97123 8925 97135 8959
rect 97077 8919 97135 8925
rect 95605 8891 95663 8897
rect 95605 8888 95617 8891
rect 93176 8860 95617 8888
rect 93176 8848 93182 8860
rect 95605 8857 95617 8860
rect 95651 8857 95663 8891
rect 95605 8851 95663 8857
rect 82832 8792 89484 8820
rect 69891 8789 69903 8792
rect 69845 8783 69903 8789
rect 89530 8780 89536 8832
rect 89588 8820 89594 8832
rect 90542 8820 90548 8832
rect 89588 8792 90548 8820
rect 89588 8780 89594 8792
rect 90542 8780 90548 8792
rect 90600 8780 90606 8832
rect 90634 8780 90640 8832
rect 90692 8820 90698 8832
rect 91005 8823 91063 8829
rect 91005 8820 91017 8823
rect 90692 8792 91017 8820
rect 90692 8780 90698 8792
rect 91005 8789 91017 8792
rect 91051 8789 91063 8823
rect 91005 8783 91063 8789
rect 94406 8780 94412 8832
rect 94464 8820 94470 8832
rect 94501 8823 94559 8829
rect 94501 8820 94513 8823
rect 94464 8792 94513 8820
rect 94464 8780 94470 8792
rect 94501 8789 94513 8792
rect 94547 8789 94559 8823
rect 94501 8783 94559 8789
rect 94866 8780 94872 8832
rect 94924 8820 94930 8832
rect 95329 8823 95387 8829
rect 95329 8820 95341 8823
rect 94924 8792 95341 8820
rect 94924 8780 94930 8792
rect 95329 8789 95341 8792
rect 95375 8789 95387 8823
rect 95329 8783 95387 8789
rect 96062 8780 96068 8832
rect 96120 8820 96126 8832
rect 97000 8820 97028 8916
rect 97092 8888 97120 8919
rect 97718 8916 97724 8968
rect 97776 8916 97782 8968
rect 97905 8959 97963 8965
rect 97905 8925 97917 8959
rect 97951 8925 97963 8959
rect 97905 8919 97963 8925
rect 97350 8888 97356 8900
rect 97092 8860 97356 8888
rect 97350 8848 97356 8860
rect 97408 8848 97414 8900
rect 97534 8848 97540 8900
rect 97592 8888 97598 8900
rect 97920 8888 97948 8919
rect 98086 8916 98092 8968
rect 98144 8916 98150 8968
rect 98546 8916 98552 8968
rect 98604 8916 98610 8968
rect 98733 8959 98791 8965
rect 98733 8925 98745 8959
rect 98779 8925 98791 8959
rect 98733 8919 98791 8925
rect 99377 8959 99435 8965
rect 99377 8925 99389 8959
rect 99423 8956 99435 8959
rect 99929 8959 99987 8965
rect 99423 8928 99512 8956
rect 99423 8925 99435 8928
rect 99377 8919 99435 8925
rect 98748 8888 98776 8919
rect 99484 8888 99512 8928
rect 99929 8925 99941 8959
rect 99975 8956 99987 8959
rect 100294 8956 100300 8968
rect 99975 8928 100300 8956
rect 99975 8925 99987 8928
rect 99929 8919 99987 8925
rect 100294 8916 100300 8928
rect 100352 8916 100358 8968
rect 100389 8959 100447 8965
rect 100389 8925 100401 8959
rect 100435 8956 100447 8959
rect 100938 8956 100944 8968
rect 100435 8928 100944 8956
rect 100435 8925 100447 8928
rect 100389 8919 100447 8925
rect 100404 8888 100432 8919
rect 100938 8916 100944 8928
rect 100996 8916 101002 8968
rect 101030 8916 101036 8968
rect 101088 8916 101094 8968
rect 101490 8916 101496 8968
rect 101548 8956 101554 8968
rect 106366 8956 106372 8968
rect 101548 8928 106372 8956
rect 101548 8916 101554 8928
rect 106366 8916 106372 8928
rect 106424 8916 106430 8968
rect 107194 8916 107200 8968
rect 107252 8916 107258 8968
rect 112346 8916 112352 8968
rect 112404 8916 112410 8968
rect 117222 8916 117228 8968
rect 117280 8956 117286 8968
rect 117501 8959 117559 8965
rect 117501 8956 117513 8959
rect 117280 8928 117513 8956
rect 117280 8916 117286 8928
rect 117501 8925 117513 8928
rect 117547 8925 117559 8959
rect 117501 8919 117559 8925
rect 120905 8959 120963 8965
rect 120905 8925 120917 8959
rect 120951 8956 120963 8959
rect 120994 8956 121000 8968
rect 120951 8928 121000 8956
rect 120951 8925 120963 8928
rect 120905 8919 120963 8925
rect 120994 8916 121000 8928
rect 121052 8916 121058 8968
rect 121641 8959 121699 8965
rect 121641 8925 121653 8959
rect 121687 8925 121699 8959
rect 121641 8919 121699 8925
rect 121733 8959 121791 8965
rect 121733 8925 121745 8959
rect 121779 8925 121791 8959
rect 121733 8919 121791 8925
rect 97592 8860 100432 8888
rect 97592 8848 97598 8860
rect 105078 8848 105084 8900
rect 105136 8888 105142 8900
rect 110598 8888 110604 8900
rect 105136 8860 110604 8888
rect 105136 8848 105142 8860
rect 110598 8848 110604 8860
rect 110656 8848 110662 8900
rect 96120 8792 97028 8820
rect 96120 8780 96126 8792
rect 97258 8780 97264 8832
rect 97316 8780 97322 8832
rect 99561 8823 99619 8829
rect 99561 8789 99573 8823
rect 99607 8820 99619 8823
rect 99650 8820 99656 8832
rect 99607 8792 99656 8820
rect 99607 8789 99619 8792
rect 99561 8783 99619 8789
rect 99650 8780 99656 8792
rect 99708 8780 99714 8832
rect 100202 8780 100208 8832
rect 100260 8820 100266 8832
rect 111334 8820 111340 8832
rect 100260 8792 111340 8820
rect 100260 8780 100266 8792
rect 111334 8780 111340 8792
rect 111392 8780 111398 8832
rect 112162 8780 112168 8832
rect 112220 8780 112226 8832
rect 116486 8780 116492 8832
rect 116544 8820 116550 8832
rect 117317 8823 117375 8829
rect 117317 8820 117329 8823
rect 116544 8792 117329 8820
rect 116544 8780 116550 8792
rect 117317 8789 117329 8792
rect 117363 8789 117375 8823
rect 121656 8820 121684 8919
rect 121748 8888 121776 8919
rect 122650 8916 122656 8968
rect 122708 8916 122714 8968
rect 123588 8965 123616 8996
rect 122745 8959 122803 8965
rect 122745 8925 122757 8959
rect 122791 8956 122803 8959
rect 123573 8959 123631 8965
rect 123573 8956 123585 8959
rect 122791 8928 123585 8956
rect 122791 8925 122803 8928
rect 122745 8919 122803 8925
rect 123573 8925 123585 8928
rect 123619 8925 123631 8959
rect 123573 8919 123631 8925
rect 121822 8888 121828 8900
rect 121748 8860 121828 8888
rect 121822 8848 121828 8860
rect 121880 8888 121886 8900
rect 122760 8888 122788 8919
rect 124122 8916 124128 8968
rect 124180 8916 124186 8968
rect 124232 8965 124260 8996
rect 124217 8959 124275 8965
rect 124217 8925 124229 8959
rect 124263 8925 124275 8959
rect 124217 8919 124275 8925
rect 124674 8916 124680 8968
rect 124732 8956 124738 8968
rect 125042 8956 125048 8968
rect 124732 8928 125048 8956
rect 124732 8916 124738 8928
rect 125042 8916 125048 8928
rect 125100 8916 125106 8968
rect 125244 8965 125272 8996
rect 125229 8959 125287 8965
rect 125229 8925 125241 8959
rect 125275 8925 125287 8959
rect 125229 8919 125287 8925
rect 125870 8916 125876 8968
rect 125928 8916 125934 8968
rect 126072 8965 126100 8996
rect 126057 8959 126115 8965
rect 126057 8925 126069 8959
rect 126103 8925 126115 8959
rect 126057 8919 126115 8925
rect 126330 8916 126336 8968
rect 126388 8956 126394 8968
rect 126698 8956 126704 8968
rect 126388 8928 126704 8956
rect 126388 8916 126394 8928
rect 126698 8916 126704 8928
rect 126756 8916 126762 8968
rect 126900 8965 126928 8996
rect 127820 8968 127848 8996
rect 128541 8993 128553 9027
rect 128587 8993 128599 9027
rect 128541 8987 128599 8993
rect 126885 8959 126943 8965
rect 126885 8925 126897 8959
rect 126931 8925 126943 8959
rect 126885 8919 126943 8925
rect 127618 8916 127624 8968
rect 127676 8916 127682 8968
rect 127802 8916 127808 8968
rect 127860 8916 127866 8968
rect 121880 8860 122788 8888
rect 121880 8848 121886 8860
rect 122834 8848 122840 8900
rect 122892 8888 122898 8900
rect 123205 8891 123263 8897
rect 123205 8888 123217 8891
rect 122892 8860 123217 8888
rect 122892 8848 122898 8860
rect 123205 8857 123217 8860
rect 123251 8857 123263 8891
rect 123205 8851 123263 8857
rect 123386 8848 123392 8900
rect 123444 8888 123450 8900
rect 128648 8888 128676 9064
rect 133874 9052 133880 9064
rect 133932 9052 133938 9104
rect 141418 9052 141424 9104
rect 141476 9092 141482 9104
rect 169662 9092 169668 9104
rect 141476 9064 169668 9092
rect 141476 9052 141482 9064
rect 169662 9052 169668 9064
rect 169720 9052 169726 9104
rect 169754 9052 169760 9104
rect 169812 9092 169818 9104
rect 170217 9095 170275 9101
rect 170217 9092 170229 9095
rect 169812 9064 170229 9092
rect 169812 9052 169818 9064
rect 170217 9061 170229 9064
rect 170263 9061 170275 9095
rect 170217 9055 170275 9061
rect 174262 9052 174268 9104
rect 174320 9052 174326 9104
rect 175274 9052 175280 9104
rect 175332 9092 175338 9104
rect 180766 9092 180794 9132
rect 184566 9120 184572 9132
rect 184624 9120 184630 9172
rect 192018 9120 192024 9172
rect 192076 9160 192082 9172
rect 192757 9163 192815 9169
rect 192757 9160 192769 9163
rect 192076 9132 192769 9160
rect 192076 9120 192082 9132
rect 192757 9129 192769 9132
rect 192803 9129 192815 9163
rect 192757 9123 192815 9129
rect 194594 9120 194600 9172
rect 194652 9160 194658 9172
rect 195793 9163 195851 9169
rect 195793 9160 195805 9163
rect 194652 9132 195805 9160
rect 194652 9120 194658 9132
rect 195793 9129 195805 9132
rect 195839 9129 195851 9163
rect 195793 9123 195851 9129
rect 197998 9120 198004 9172
rect 198056 9160 198062 9172
rect 199105 9163 199163 9169
rect 199105 9160 199117 9163
rect 198056 9132 199117 9160
rect 198056 9120 198062 9132
rect 199105 9129 199117 9132
rect 199151 9129 199163 9163
rect 199105 9123 199163 9129
rect 199746 9120 199752 9172
rect 199804 9160 199810 9172
rect 200114 9160 200120 9172
rect 199804 9132 200120 9160
rect 199804 9120 199810 9132
rect 200114 9120 200120 9132
rect 200172 9120 200178 9172
rect 200666 9120 200672 9172
rect 200724 9160 200730 9172
rect 203334 9160 203340 9172
rect 200724 9132 203340 9160
rect 200724 9120 200730 9132
rect 203334 9120 203340 9132
rect 203392 9120 203398 9172
rect 203426 9120 203432 9172
rect 203484 9120 203490 9172
rect 204070 9120 204076 9172
rect 204128 9120 204134 9172
rect 204180 9132 228312 9160
rect 175332 9064 180794 9092
rect 175332 9052 175338 9064
rect 182082 9052 182088 9104
rect 182140 9052 182146 9104
rect 194502 9092 194508 9104
rect 182376 9064 194508 9092
rect 128814 8984 128820 9036
rect 128872 9024 128878 9036
rect 145006 9024 145012 9036
rect 128872 8996 133920 9024
rect 128872 8984 128878 8996
rect 130102 8916 130108 8968
rect 130160 8956 130166 8968
rect 130396 8965 130424 8996
rect 130197 8959 130255 8965
rect 130197 8956 130209 8959
rect 130160 8928 130209 8956
rect 130160 8916 130166 8928
rect 130197 8925 130209 8928
rect 130243 8925 130255 8959
rect 130197 8919 130255 8925
rect 130381 8959 130439 8965
rect 130381 8925 130393 8959
rect 130427 8925 130439 8959
rect 130381 8919 130439 8925
rect 131025 8959 131083 8965
rect 131025 8925 131037 8959
rect 131071 8956 131083 8959
rect 131114 8956 131120 8968
rect 131071 8928 131120 8956
rect 131071 8925 131083 8928
rect 131025 8919 131083 8925
rect 131114 8916 131120 8928
rect 131172 8916 131178 8968
rect 131224 8965 131252 8996
rect 131209 8959 131267 8965
rect 131209 8925 131221 8959
rect 131255 8925 131267 8959
rect 131209 8919 131267 8925
rect 131850 8916 131856 8968
rect 131908 8916 131914 8968
rect 132052 8965 132080 8996
rect 132880 8968 132908 8996
rect 132037 8959 132095 8965
rect 132037 8925 132049 8959
rect 132083 8925 132095 8959
rect 132037 8919 132095 8925
rect 132586 8916 132592 8968
rect 132644 8956 132650 8968
rect 132770 8956 132776 8968
rect 132644 8928 132776 8956
rect 132644 8916 132650 8928
rect 132770 8916 132776 8928
rect 132828 8916 132834 8968
rect 132862 8916 132868 8968
rect 132920 8916 132926 8968
rect 133782 8916 133788 8968
rect 133840 8916 133846 8968
rect 133892 8965 133920 8996
rect 137986 8996 145012 9024
rect 133877 8959 133935 8965
rect 133877 8925 133889 8959
rect 133923 8925 133935 8959
rect 133877 8919 133935 8925
rect 134518 8916 134524 8968
rect 134576 8916 134582 8968
rect 123444 8860 128676 8888
rect 123444 8848 123450 8860
rect 130838 8848 130844 8900
rect 130896 8888 130902 8900
rect 137986 8888 138014 8996
rect 145006 8984 145012 8996
rect 145064 8984 145070 9036
rect 149606 8984 149612 9036
rect 149664 9024 149670 9036
rect 149664 8996 150204 9024
rect 149664 8984 149670 8996
rect 139762 8916 139768 8968
rect 139820 8916 139826 8968
rect 144914 8916 144920 8968
rect 144972 8916 144978 8968
rect 150066 8916 150072 8968
rect 150124 8916 150130 8968
rect 150176 8956 150204 8996
rect 150802 8984 150808 9036
rect 150860 9024 150866 9036
rect 153470 9024 153476 9036
rect 150860 8996 153476 9024
rect 150860 8984 150866 8996
rect 153470 8984 153476 8996
rect 153528 8984 153534 9036
rect 156046 9024 156052 9036
rect 153580 8996 156052 9024
rect 153580 8956 153608 8996
rect 156046 8984 156052 8996
rect 156104 8984 156110 9036
rect 156141 9027 156199 9033
rect 156141 8993 156153 9027
rect 156187 9024 156199 9027
rect 156690 9024 156696 9036
rect 156187 8996 156696 9024
rect 156187 8993 156199 8996
rect 156141 8987 156199 8993
rect 156690 8984 156696 8996
rect 156748 8984 156754 9036
rect 157334 8984 157340 9036
rect 157392 8984 157398 9036
rect 157426 8984 157432 9036
rect 157484 9024 157490 9036
rect 157484 8996 171824 9024
rect 157484 8984 157490 8996
rect 150176 8928 153608 8956
rect 155218 8916 155224 8968
rect 155276 8916 155282 8968
rect 156325 8959 156383 8965
rect 156325 8925 156337 8959
rect 156371 8958 156383 8959
rect 156371 8930 156460 8958
rect 156371 8925 156383 8930
rect 156325 8919 156383 8925
rect 130896 8860 138014 8888
rect 130896 8848 130902 8860
rect 142798 8848 142804 8900
rect 142856 8888 142862 8900
rect 156230 8888 156236 8900
rect 142856 8860 156236 8888
rect 142856 8848 142862 8860
rect 156230 8848 156236 8860
rect 156288 8848 156294 8900
rect 156432 8888 156460 8930
rect 157058 8916 157064 8968
rect 157116 8916 157122 8968
rect 157153 8959 157211 8965
rect 157153 8925 157165 8959
rect 157199 8956 157211 8959
rect 157518 8956 157524 8968
rect 157199 8928 157524 8956
rect 157199 8925 157211 8928
rect 157153 8919 157211 8925
rect 157168 8888 157196 8919
rect 157518 8916 157524 8928
rect 157576 8916 157582 8968
rect 158625 8959 158683 8965
rect 158625 8925 158637 8959
rect 158671 8956 158683 8959
rect 159634 8956 159640 8968
rect 158671 8928 159640 8956
rect 158671 8925 158683 8928
rect 158625 8919 158683 8925
rect 159634 8916 159640 8928
rect 159692 8916 159698 8968
rect 160373 8959 160431 8965
rect 160373 8925 160385 8959
rect 160419 8956 160431 8959
rect 161569 8959 161627 8965
rect 160419 8928 161520 8956
rect 160419 8925 160431 8928
rect 160373 8919 160431 8925
rect 156432 8860 157196 8888
rect 157794 8848 157800 8900
rect 157852 8888 157858 8900
rect 159174 8888 159180 8900
rect 157852 8860 159180 8888
rect 157852 8848 157858 8860
rect 159174 8848 159180 8860
rect 159232 8848 159238 8900
rect 161017 8891 161075 8897
rect 161017 8857 161029 8891
rect 161063 8888 161075 8891
rect 161106 8888 161112 8900
rect 161063 8860 161112 8888
rect 161063 8857 161075 8860
rect 161017 8851 161075 8857
rect 161106 8848 161112 8860
rect 161164 8848 161170 8900
rect 161492 8888 161520 8928
rect 161569 8925 161581 8959
rect 161615 8956 161627 8959
rect 161934 8956 161940 8968
rect 161615 8928 161940 8956
rect 161615 8925 161627 8928
rect 161569 8919 161627 8925
rect 161934 8916 161940 8928
rect 161992 8916 161998 8968
rect 162854 8956 162860 8968
rect 162044 8928 162860 8956
rect 162044 8888 162072 8928
rect 162854 8916 162860 8928
rect 162912 8916 162918 8968
rect 163133 8959 163191 8965
rect 163133 8925 163145 8959
rect 163179 8956 163191 8959
rect 163774 8956 163780 8968
rect 163179 8928 163780 8956
rect 163179 8925 163191 8928
rect 163133 8919 163191 8925
rect 163774 8916 163780 8928
rect 163832 8916 163838 8968
rect 164973 8959 165031 8965
rect 164973 8925 164985 8959
rect 165019 8956 165031 8959
rect 165019 8928 166028 8956
rect 165019 8925 165031 8928
rect 164973 8919 165031 8925
rect 161492 8860 162072 8888
rect 162302 8848 162308 8900
rect 162360 8848 162366 8900
rect 162578 8848 162584 8900
rect 162636 8888 162642 8900
rect 162762 8888 162768 8900
rect 162636 8860 162768 8888
rect 162636 8848 162642 8860
rect 162762 8848 162768 8860
rect 162820 8888 162826 8900
rect 164145 8891 164203 8897
rect 164145 8888 164157 8891
rect 162820 8860 164157 8888
rect 162820 8848 162826 8860
rect 164145 8857 164157 8860
rect 164191 8857 164203 8891
rect 164145 8851 164203 8857
rect 164510 8848 164516 8900
rect 164568 8888 164574 8900
rect 165341 8891 165399 8897
rect 165341 8888 165353 8891
rect 164568 8860 165353 8888
rect 164568 8848 164574 8860
rect 165341 8857 165353 8860
rect 165387 8857 165399 8891
rect 165341 8851 165399 8857
rect 121730 8820 121736 8832
rect 121656 8792 121736 8820
rect 117317 8783 117375 8789
rect 121730 8780 121736 8792
rect 121788 8780 121794 8832
rect 121917 8823 121975 8829
rect 121917 8789 121929 8823
rect 121963 8820 121975 8823
rect 122190 8820 122196 8832
rect 121963 8792 122196 8820
rect 121963 8789 121975 8792
rect 121917 8783 121975 8789
rect 122190 8780 122196 8792
rect 122248 8780 122254 8832
rect 122929 8823 122987 8829
rect 122929 8789 122941 8823
rect 122975 8820 122987 8823
rect 123018 8820 123024 8832
rect 122975 8792 123024 8820
rect 122975 8789 122987 8792
rect 122929 8783 122987 8789
rect 123018 8780 123024 8792
rect 123076 8780 123082 8832
rect 123757 8823 123815 8829
rect 123757 8789 123769 8823
rect 123803 8820 123815 8823
rect 123846 8820 123852 8832
rect 123803 8792 123852 8820
rect 123803 8789 123815 8792
rect 123757 8783 123815 8789
rect 123846 8780 123852 8792
rect 123904 8780 123910 8832
rect 125410 8780 125416 8832
rect 125468 8780 125474 8832
rect 126790 8780 126796 8832
rect 126848 8820 126854 8832
rect 127069 8823 127127 8829
rect 127069 8820 127081 8823
rect 126848 8792 127081 8820
rect 126848 8780 126854 8792
rect 127069 8789 127081 8792
rect 127115 8789 127127 8823
rect 127069 8783 127127 8789
rect 127526 8780 127532 8832
rect 127584 8820 127590 8832
rect 127989 8823 128047 8829
rect 127989 8820 128001 8823
rect 127584 8792 128001 8820
rect 127584 8780 127590 8792
rect 127989 8789 128001 8792
rect 128035 8789 128047 8823
rect 127989 8783 128047 8789
rect 131942 8780 131948 8832
rect 132000 8820 132006 8832
rect 132221 8823 132279 8829
rect 132221 8820 132233 8823
rect 132000 8792 132233 8820
rect 132000 8780 132006 8792
rect 132221 8789 132233 8792
rect 132267 8789 132279 8823
rect 132221 8783 132279 8789
rect 133417 8823 133475 8829
rect 133417 8789 133429 8823
rect 133463 8820 133475 8823
rect 133874 8820 133880 8832
rect 133463 8792 133880 8820
rect 133463 8789 133475 8792
rect 133417 8783 133475 8789
rect 133874 8780 133880 8792
rect 133932 8820 133938 8832
rect 134150 8820 134156 8832
rect 133932 8792 134156 8820
rect 133932 8780 133938 8792
rect 134150 8780 134156 8792
rect 134208 8780 134214 8832
rect 139302 8780 139308 8832
rect 139360 8820 139366 8832
rect 139581 8823 139639 8829
rect 139581 8820 139593 8823
rect 139360 8792 139593 8820
rect 139360 8780 139366 8792
rect 139581 8789 139593 8792
rect 139627 8789 139639 8823
rect 139581 8783 139639 8789
rect 144730 8780 144736 8832
rect 144788 8780 144794 8832
rect 149885 8823 149943 8829
rect 149885 8789 149897 8823
rect 149931 8820 149943 8823
rect 150342 8820 150348 8832
rect 149931 8792 150348 8820
rect 149931 8789 149943 8792
rect 149885 8783 149943 8789
rect 150342 8780 150348 8792
rect 150400 8780 150406 8832
rect 155034 8780 155040 8832
rect 155092 8780 155098 8832
rect 155954 8780 155960 8832
rect 156012 8820 156018 8832
rect 156509 8823 156567 8829
rect 156509 8820 156521 8823
rect 156012 8792 156521 8820
rect 156012 8780 156018 8792
rect 156509 8789 156521 8792
rect 156555 8789 156567 8823
rect 156509 8783 156567 8789
rect 161842 8780 161848 8832
rect 161900 8820 161906 8832
rect 165798 8820 165804 8832
rect 161900 8792 165804 8820
rect 161900 8780 161906 8792
rect 165798 8780 165804 8792
rect 165856 8780 165862 8832
rect 166000 8829 166028 8928
rect 166166 8916 166172 8968
rect 166224 8916 166230 8968
rect 166442 8916 166448 8968
rect 166500 8956 166506 8968
rect 166537 8959 166595 8965
rect 166537 8956 166549 8959
rect 166500 8928 166549 8956
rect 166500 8916 166506 8928
rect 166537 8925 166549 8928
rect 166583 8925 166595 8959
rect 166537 8919 166595 8925
rect 167365 8959 167423 8965
rect 167365 8925 167377 8959
rect 167411 8956 167423 8959
rect 168742 8956 168748 8968
rect 167411 8928 168748 8956
rect 167411 8925 167423 8928
rect 167365 8919 167423 8925
rect 168742 8916 168748 8928
rect 168800 8916 168806 8968
rect 168926 8916 168932 8968
rect 168984 8916 168990 8968
rect 169018 8916 169024 8968
rect 169076 8956 169082 8968
rect 170033 8959 170091 8965
rect 170033 8956 170045 8959
rect 169076 8928 170045 8956
rect 169076 8916 169082 8928
rect 170033 8925 170045 8928
rect 170079 8925 170091 8959
rect 170033 8919 170091 8925
rect 167086 8848 167092 8900
rect 167144 8888 167150 8900
rect 167733 8891 167791 8897
rect 167733 8888 167745 8891
rect 167144 8860 167745 8888
rect 167144 8848 167150 8860
rect 167733 8857 167745 8860
rect 167779 8857 167791 8891
rect 167733 8851 167791 8857
rect 167822 8848 167828 8900
rect 167880 8888 167886 8900
rect 169297 8891 169355 8897
rect 169297 8888 169309 8891
rect 167880 8860 169309 8888
rect 167880 8848 167886 8860
rect 169297 8857 169309 8860
rect 169343 8857 169355 8891
rect 171796 8888 171824 8996
rect 171870 8984 171876 9036
rect 171928 9024 171934 9036
rect 182376 9024 182404 9064
rect 194502 9052 194508 9064
rect 194560 9052 194566 9104
rect 194686 9052 194692 9104
rect 194744 9092 194750 9104
rect 195330 9092 195336 9104
rect 194744 9064 195336 9092
rect 194744 9052 194750 9064
rect 195330 9052 195336 9064
rect 195388 9052 195394 9104
rect 195514 9052 195520 9104
rect 195572 9092 195578 9104
rect 195572 9064 199976 9092
rect 195572 9052 195578 9064
rect 171928 8996 182404 9024
rect 171928 8984 171934 8996
rect 184290 8984 184296 9036
rect 184348 8984 184354 9036
rect 184750 8984 184756 9036
rect 184808 9024 184814 9036
rect 185581 9027 185639 9033
rect 185581 9024 185593 9027
rect 184808 8996 185593 9024
rect 184808 8984 184814 8996
rect 185581 8993 185593 8996
rect 185627 8993 185639 9027
rect 185581 8987 185639 8993
rect 186222 8984 186228 9036
rect 186280 9024 186286 9036
rect 186869 9027 186927 9033
rect 186869 9024 186881 9027
rect 186280 8996 186881 9024
rect 186280 8984 186286 8996
rect 186869 8993 186881 8996
rect 186915 8993 186927 9027
rect 186869 8987 186927 8993
rect 189442 8984 189448 9036
rect 189500 8984 189506 9036
rect 190822 8984 190828 9036
rect 190880 9024 190886 9036
rect 197633 9027 197691 9033
rect 197633 9024 197645 9027
rect 190880 8996 197645 9024
rect 190880 8984 190886 8996
rect 197633 8993 197645 8996
rect 197679 8993 197691 9027
rect 197633 8987 197691 8993
rect 197722 8984 197728 9036
rect 197780 9024 197786 9036
rect 197909 9027 197967 9033
rect 197909 9024 197921 9027
rect 197780 8996 197921 9024
rect 197780 8984 197786 8996
rect 197909 8993 197921 8996
rect 197955 9024 197967 9027
rect 199948 9024 199976 9064
rect 201310 9052 201316 9104
rect 201368 9092 201374 9104
rect 204180 9092 204208 9132
rect 201368 9064 204208 9092
rect 201368 9052 201374 9064
rect 204254 9052 204260 9104
rect 204312 9092 204318 9104
rect 220262 9092 220268 9104
rect 204312 9064 220268 9092
rect 204312 9052 204318 9064
rect 220262 9052 220268 9064
rect 220320 9052 220326 9104
rect 223666 9092 223672 9104
rect 221568 9064 223672 9092
rect 220078 9024 220084 9036
rect 197955 8996 199884 9024
rect 199948 8996 220084 9024
rect 197955 8993 197967 8996
rect 197909 8987 197967 8993
rect 173894 8916 173900 8968
rect 173952 8956 173958 8968
rect 174081 8959 174139 8965
rect 174081 8956 174093 8959
rect 173952 8928 174093 8956
rect 173952 8916 173958 8928
rect 174081 8925 174093 8928
rect 174127 8925 174139 8959
rect 174081 8919 174139 8925
rect 175182 8916 175188 8968
rect 175240 8956 175246 8968
rect 175277 8959 175335 8965
rect 175277 8956 175289 8959
rect 175240 8928 175289 8956
rect 175240 8916 175246 8928
rect 175277 8925 175289 8928
rect 175323 8925 175335 8959
rect 175277 8919 175335 8925
rect 176746 8916 176752 8968
rect 176804 8916 176810 8968
rect 177482 8916 177488 8968
rect 177540 8916 177546 8968
rect 180426 8916 180432 8968
rect 180484 8916 180490 8968
rect 181898 8916 181904 8968
rect 181956 8916 181962 8968
rect 184569 8959 184627 8965
rect 184569 8925 184581 8959
rect 184615 8925 184627 8959
rect 184569 8919 184627 8925
rect 180613 8891 180671 8897
rect 180613 8888 180625 8891
rect 171796 8860 180625 8888
rect 169297 8851 169355 8857
rect 180613 8857 180625 8860
rect 180659 8857 180671 8891
rect 184584 8888 184612 8919
rect 185854 8916 185860 8968
rect 185912 8916 185918 8968
rect 187145 8959 187203 8965
rect 187145 8925 187157 8959
rect 187191 8925 187203 8959
rect 187145 8919 187203 8925
rect 180613 8851 180671 8857
rect 180766 8860 184612 8888
rect 165985 8823 166043 8829
rect 165985 8789 165997 8823
rect 166031 8820 166043 8823
rect 168834 8820 168840 8832
rect 166031 8792 168840 8820
rect 166031 8789 166043 8792
rect 165985 8783 166043 8789
rect 168834 8780 168840 8792
rect 168892 8780 168898 8832
rect 168926 8780 168932 8832
rect 168984 8820 168990 8832
rect 171042 8820 171048 8832
rect 168984 8792 171048 8820
rect 168984 8780 168990 8792
rect 171042 8780 171048 8792
rect 171100 8780 171106 8832
rect 172698 8780 172704 8832
rect 172756 8820 172762 8832
rect 175369 8823 175427 8829
rect 175369 8820 175381 8823
rect 172756 8792 175381 8820
rect 172756 8780 172762 8792
rect 175369 8789 175381 8792
rect 175415 8789 175427 8823
rect 175369 8783 175427 8789
rect 177666 8780 177672 8832
rect 177724 8820 177730 8832
rect 180766 8820 180794 8860
rect 177724 8792 180794 8820
rect 177724 8780 177730 8792
rect 182082 8780 182088 8832
rect 182140 8820 182146 8832
rect 187160 8820 187188 8919
rect 189718 8916 189724 8968
rect 189776 8916 189782 8968
rect 190638 8916 190644 8968
rect 190696 8956 190702 8968
rect 190733 8959 190791 8965
rect 190733 8956 190745 8959
rect 190696 8928 190745 8956
rect 190696 8916 190702 8928
rect 190733 8925 190745 8928
rect 190779 8925 190791 8959
rect 190733 8919 190791 8925
rect 190914 8916 190920 8968
rect 190972 8916 190978 8968
rect 191006 8916 191012 8968
rect 191064 8956 191070 8968
rect 191561 8959 191619 8965
rect 191561 8956 191573 8959
rect 191064 8928 191573 8956
rect 191064 8916 191070 8928
rect 191561 8925 191573 8928
rect 191607 8925 191619 8959
rect 191561 8919 191619 8925
rect 191745 8959 191803 8965
rect 191745 8925 191757 8959
rect 191791 8925 191803 8959
rect 191745 8919 191803 8925
rect 190932 8888 190960 8916
rect 191760 8888 191788 8919
rect 192110 8916 192116 8968
rect 192168 8956 192174 8968
rect 192389 8959 192447 8965
rect 192389 8956 192401 8959
rect 192168 8928 192401 8956
rect 192168 8916 192174 8928
rect 192389 8925 192401 8928
rect 192435 8925 192447 8959
rect 192389 8919 192447 8925
rect 192573 8959 192631 8965
rect 192573 8925 192585 8959
rect 192619 8925 192631 8959
rect 192573 8919 192631 8925
rect 192478 8888 192484 8900
rect 190932 8860 192484 8888
rect 192478 8848 192484 8860
rect 192536 8888 192542 8900
rect 192588 8888 192616 8919
rect 193306 8916 193312 8968
rect 193364 8916 193370 8968
rect 193401 8959 193459 8965
rect 193401 8925 193413 8959
rect 193447 8925 193459 8959
rect 193401 8919 193459 8925
rect 193416 8888 193444 8919
rect 194686 8916 194692 8968
rect 194744 8916 194750 8968
rect 194781 8959 194839 8965
rect 194781 8925 194793 8959
rect 194827 8925 194839 8959
rect 194781 8919 194839 8925
rect 194796 8888 194824 8919
rect 195514 8916 195520 8968
rect 195572 8916 195578 8968
rect 195609 8959 195667 8965
rect 195609 8925 195621 8959
rect 195655 8925 195667 8959
rect 195609 8919 195667 8925
rect 195624 8888 195652 8919
rect 196342 8916 196348 8968
rect 196400 8916 196406 8968
rect 196437 8959 196495 8965
rect 196437 8925 196449 8959
rect 196483 8925 196495 8959
rect 196437 8919 196495 8925
rect 195974 8888 195980 8900
rect 192536 8860 195980 8888
rect 192536 8848 192542 8860
rect 195974 8848 195980 8860
rect 196032 8888 196038 8900
rect 196452 8888 196480 8919
rect 198550 8916 198556 8968
rect 198608 8956 198614 8968
rect 198921 8959 198979 8965
rect 198921 8956 198933 8959
rect 198608 8928 198933 8956
rect 198608 8916 198614 8928
rect 198921 8925 198933 8928
rect 198967 8925 198979 8959
rect 198921 8919 198979 8925
rect 199746 8916 199752 8968
rect 199804 8916 199810 8968
rect 199856 8956 199884 8996
rect 220078 8984 220084 8996
rect 220136 8984 220142 9036
rect 220170 8984 220176 9036
rect 220228 9024 220234 9036
rect 221568 9024 221596 9064
rect 223666 9052 223672 9064
rect 223724 9052 223730 9104
rect 223758 9052 223764 9104
rect 223816 9052 223822 9104
rect 225414 9092 225420 9104
rect 223868 9064 225420 9092
rect 220228 8996 221596 9024
rect 220228 8984 220234 8996
rect 221642 8984 221648 9036
rect 221700 9024 221706 9036
rect 223868 9024 223896 9064
rect 225414 9052 225420 9064
rect 225472 9052 225478 9104
rect 228284 9092 228312 9132
rect 228358 9120 228364 9172
rect 228416 9120 228422 9172
rect 228542 9120 228548 9172
rect 228600 9160 228606 9172
rect 228600 9132 230704 9160
rect 228600 9120 228606 9132
rect 230566 9092 230572 9104
rect 228284 9064 230572 9092
rect 230566 9052 230572 9064
rect 230624 9052 230630 9104
rect 230676 9092 230704 9132
rect 230934 9120 230940 9172
rect 230992 9160 230998 9172
rect 230992 9132 233556 9160
rect 230992 9120 230998 9132
rect 233528 9092 233556 9132
rect 233970 9120 233976 9172
rect 234028 9120 234034 9172
rect 234706 9120 234712 9172
rect 234764 9160 234770 9172
rect 235626 9160 235632 9172
rect 234764 9132 235632 9160
rect 234764 9120 234770 9132
rect 235626 9120 235632 9132
rect 235684 9160 235690 9172
rect 236454 9160 236460 9172
rect 235684 9132 236460 9160
rect 235684 9120 235690 9132
rect 236454 9120 236460 9132
rect 236512 9120 236518 9172
rect 236822 9120 236828 9172
rect 236880 9120 236886 9172
rect 244918 9120 244924 9172
rect 244976 9160 244982 9172
rect 249702 9160 249708 9172
rect 244976 9132 249708 9160
rect 244976 9120 244982 9132
rect 249702 9120 249708 9132
rect 249760 9120 249766 9172
rect 249794 9120 249800 9172
rect 249852 9160 249858 9172
rect 252511 9163 252569 9169
rect 252511 9160 252523 9163
rect 249852 9132 252523 9160
rect 249852 9120 249858 9132
rect 252511 9129 252523 9132
rect 252557 9129 252569 9163
rect 252511 9123 252569 9129
rect 254670 9120 254676 9172
rect 254728 9160 254734 9172
rect 258718 9160 258724 9172
rect 254728 9132 258724 9160
rect 254728 9120 254734 9132
rect 258718 9120 258724 9132
rect 258776 9120 258782 9172
rect 259362 9120 259368 9172
rect 259420 9120 259426 9172
rect 261662 9120 261668 9172
rect 261720 9160 261726 9172
rect 261757 9163 261815 9169
rect 261757 9160 261769 9163
rect 261720 9132 261769 9160
rect 261720 9120 261726 9132
rect 261757 9129 261769 9132
rect 261803 9129 261815 9163
rect 261757 9123 261815 9129
rect 262122 9120 262128 9172
rect 262180 9160 262186 9172
rect 262677 9163 262735 9169
rect 262677 9160 262689 9163
rect 262180 9132 262689 9160
rect 262180 9120 262186 9132
rect 262677 9129 262689 9132
rect 262723 9129 262735 9163
rect 262677 9123 262735 9129
rect 265066 9120 265072 9172
rect 265124 9160 265130 9172
rect 268654 9160 268660 9172
rect 265124 9132 268660 9160
rect 265124 9120 265130 9132
rect 268654 9120 268660 9132
rect 268712 9120 268718 9172
rect 270402 9120 270408 9172
rect 270460 9160 270466 9172
rect 270589 9163 270647 9169
rect 270589 9160 270601 9163
rect 270460 9132 270601 9160
rect 270460 9120 270466 9132
rect 270589 9129 270601 9132
rect 270635 9129 270647 9163
rect 270589 9123 270647 9129
rect 254762 9092 254768 9104
rect 230676 9064 233004 9092
rect 233528 9064 254768 9092
rect 221700 8996 223896 9024
rect 224236 8996 224448 9024
rect 221700 8984 221706 8996
rect 199933 8959 199991 8965
rect 199933 8956 199945 8959
rect 199856 8928 199945 8956
rect 199933 8925 199945 8928
rect 199979 8925 199991 8959
rect 199933 8919 199991 8925
rect 196032 8860 196480 8888
rect 199948 8888 199976 8919
rect 200666 8916 200672 8968
rect 200724 8916 200730 8968
rect 200761 8959 200819 8965
rect 200761 8925 200773 8959
rect 200807 8925 200819 8959
rect 200761 8919 200819 8925
rect 200776 8888 200804 8919
rect 201310 8916 201316 8968
rect 201368 8956 201374 8968
rect 201405 8959 201463 8965
rect 201405 8956 201417 8959
rect 201368 8928 201417 8956
rect 201368 8916 201374 8928
rect 201405 8925 201417 8928
rect 201451 8925 201463 8959
rect 201405 8919 201463 8925
rect 201589 8959 201647 8965
rect 201589 8925 201601 8959
rect 201635 8925 201647 8959
rect 201589 8919 201647 8925
rect 201604 8888 201632 8919
rect 202322 8916 202328 8968
rect 202380 8916 202386 8968
rect 202417 8959 202475 8965
rect 202417 8925 202429 8959
rect 202463 8925 202475 8959
rect 202417 8919 202475 8925
rect 202432 8888 202460 8919
rect 203058 8916 203064 8968
rect 203116 8916 203122 8968
rect 203245 8959 203303 8965
rect 203245 8925 203257 8959
rect 203291 8925 203303 8959
rect 203245 8919 203303 8925
rect 202506 8888 202512 8900
rect 199948 8860 202512 8888
rect 196032 8848 196038 8860
rect 202506 8848 202512 8860
rect 202564 8888 202570 8900
rect 203260 8888 203288 8919
rect 203518 8916 203524 8968
rect 203576 8956 203582 8968
rect 203889 8959 203947 8965
rect 203889 8956 203901 8959
rect 203576 8928 203901 8956
rect 203576 8916 203582 8928
rect 203889 8925 203901 8928
rect 203935 8925 203947 8959
rect 203889 8919 203947 8925
rect 211706 8916 211712 8968
rect 211764 8916 211770 8968
rect 211798 8916 211804 8968
rect 211856 8956 211862 8968
rect 215110 8956 215116 8968
rect 211856 8928 215116 8956
rect 211856 8916 211862 8928
rect 215110 8916 215116 8928
rect 215168 8916 215174 8968
rect 216858 8916 216864 8968
rect 216916 8916 216922 8968
rect 222010 8916 222016 8968
rect 222068 8916 222074 8968
rect 223022 8916 223028 8968
rect 223080 8956 223086 8968
rect 223393 8959 223451 8965
rect 223393 8956 223405 8959
rect 223080 8928 223405 8956
rect 223080 8916 223086 8928
rect 223393 8925 223405 8928
rect 223439 8925 223451 8959
rect 223393 8919 223451 8925
rect 223577 8959 223635 8965
rect 223577 8925 223589 8959
rect 223623 8956 223635 8959
rect 224236 8956 224264 8996
rect 224420 8968 224448 8996
rect 224586 8984 224592 9036
rect 224644 9024 224650 9036
rect 230661 9027 230719 9033
rect 230661 9024 230673 9027
rect 224644 8996 230673 9024
rect 224644 8984 224650 8996
rect 230661 8993 230673 8996
rect 230707 8993 230719 9027
rect 230661 8987 230719 8993
rect 232774 8984 232780 9036
rect 232832 8984 232838 9036
rect 232976 9024 233004 9064
rect 254762 9052 254768 9064
rect 254820 9052 254826 9104
rect 254946 9052 254952 9104
rect 255004 9092 255010 9104
rect 263226 9092 263232 9104
rect 255004 9064 263232 9092
rect 255004 9052 255010 9064
rect 263226 9052 263232 9064
rect 263284 9052 263290 9104
rect 263686 9052 263692 9104
rect 263744 9092 263750 9104
rect 267918 9092 267924 9104
rect 263744 9064 267924 9092
rect 263744 9052 263750 9064
rect 267918 9052 267924 9064
rect 267976 9052 267982 9104
rect 268470 9052 268476 9104
rect 268528 9092 268534 9104
rect 268841 9095 268899 9101
rect 268841 9092 268853 9095
rect 268528 9064 268853 9092
rect 268528 9052 268534 9064
rect 268841 9061 268853 9064
rect 268887 9061 268899 9095
rect 268841 9055 268899 9061
rect 254670 9024 254676 9036
rect 232976 8996 254676 9024
rect 254670 8984 254676 8996
rect 254728 8984 254734 9036
rect 255038 8984 255044 9036
rect 255096 8984 255102 9036
rect 256418 8984 256424 9036
rect 256476 8984 256482 9036
rect 257706 8984 257712 9036
rect 257764 8984 257770 9036
rect 257890 8984 257896 9036
rect 257948 9024 257954 9036
rect 260742 9024 260748 9036
rect 257948 8996 260748 9024
rect 257948 8984 257954 8996
rect 260742 8984 260748 8996
rect 260800 9024 260806 9036
rect 260800 8996 261708 9024
rect 260800 8984 260806 8996
rect 223623 8928 224264 8956
rect 223623 8925 223635 8928
rect 223577 8919 223635 8925
rect 224310 8916 224316 8968
rect 224368 8916 224374 8968
rect 224402 8916 224408 8968
rect 224460 8956 224466 8968
rect 224460 8928 225552 8956
rect 224460 8916 224466 8928
rect 202564 8860 203288 8888
rect 202564 8848 202570 8860
rect 203334 8848 203340 8900
rect 203392 8888 203398 8900
rect 225138 8888 225144 8900
rect 203392 8860 225144 8888
rect 203392 8848 203398 8860
rect 225138 8848 225144 8860
rect 225196 8848 225202 8900
rect 225524 8888 225552 8928
rect 225598 8916 225604 8968
rect 225656 8916 225662 8968
rect 225693 8959 225751 8965
rect 225693 8925 225705 8959
rect 225739 8925 225751 8959
rect 225693 8919 225751 8925
rect 225708 8888 225736 8919
rect 226426 8916 226432 8968
rect 226484 8916 226490 8968
rect 226521 8959 226579 8965
rect 226521 8925 226533 8959
rect 226567 8925 226579 8959
rect 226521 8919 226579 8925
rect 226536 8888 226564 8919
rect 227162 8916 227168 8968
rect 227220 8916 227226 8968
rect 227349 8959 227407 8965
rect 227349 8925 227361 8959
rect 227395 8925 227407 8959
rect 227349 8919 227407 8925
rect 227364 8888 227392 8919
rect 228082 8916 228088 8968
rect 228140 8916 228146 8968
rect 228177 8959 228235 8965
rect 228177 8925 228189 8959
rect 228223 8925 228235 8959
rect 228177 8919 228235 8925
rect 228192 8888 228220 8919
rect 228818 8916 228824 8968
rect 228876 8916 228882 8968
rect 229005 8959 229063 8965
rect 229005 8956 229017 8959
rect 228928 8928 229017 8956
rect 228266 8888 228272 8900
rect 225524 8860 228272 8888
rect 228266 8848 228272 8860
rect 228324 8888 228330 8900
rect 228928 8888 228956 8928
rect 229005 8925 229017 8928
rect 229051 8956 229063 8959
rect 229051 8928 229140 8956
rect 229051 8925 229063 8928
rect 229005 8919 229063 8925
rect 228324 8860 228956 8888
rect 229112 8888 229140 8928
rect 229646 8916 229652 8968
rect 229704 8916 229710 8968
rect 229833 8959 229891 8965
rect 229833 8925 229845 8959
rect 229879 8925 229891 8959
rect 229833 8919 229891 8925
rect 229848 8888 229876 8919
rect 230014 8916 230020 8968
rect 230072 8916 230078 8968
rect 230106 8916 230112 8968
rect 230164 8956 230170 8968
rect 230842 8956 230848 8968
rect 230164 8928 230848 8956
rect 230164 8916 230170 8928
rect 230842 8916 230848 8928
rect 230900 8956 230906 8968
rect 230937 8959 230995 8965
rect 230937 8956 230949 8959
rect 230900 8928 230949 8956
rect 230900 8916 230906 8928
rect 230937 8925 230949 8928
rect 230983 8925 230995 8959
rect 230937 8919 230995 8925
rect 230198 8888 230204 8900
rect 229112 8860 230204 8888
rect 228324 8848 228330 8860
rect 230198 8848 230204 8860
rect 230256 8848 230262 8900
rect 230658 8848 230664 8900
rect 230716 8848 230722 8900
rect 230952 8888 230980 8919
rect 231854 8916 231860 8968
rect 231912 8956 231918 8968
rect 231949 8959 232007 8965
rect 231949 8956 231961 8959
rect 231912 8928 231961 8956
rect 231912 8916 231918 8928
rect 231949 8925 231961 8928
rect 231995 8956 232007 8959
rect 232038 8956 232044 8968
rect 231995 8928 232044 8956
rect 231995 8925 232007 8928
rect 231949 8919 232007 8925
rect 232038 8916 232044 8928
rect 232096 8916 232102 8968
rect 232133 8959 232191 8965
rect 232133 8925 232145 8959
rect 232179 8925 232191 8959
rect 232133 8919 232191 8925
rect 232148 8888 232176 8919
rect 232314 8916 232320 8968
rect 232372 8916 232378 8968
rect 232961 8959 233019 8965
rect 232961 8958 232973 8959
rect 232884 8930 232973 8958
rect 232884 8888 232912 8930
rect 232961 8925 232973 8930
rect 233007 8925 233019 8959
rect 232961 8919 233019 8925
rect 233602 8916 233608 8968
rect 233660 8916 233666 8968
rect 233789 8959 233847 8965
rect 233789 8925 233801 8959
rect 233835 8925 233847 8959
rect 233789 8919 233847 8925
rect 233694 8888 233700 8900
rect 230952 8860 233700 8888
rect 233694 8848 233700 8860
rect 233752 8888 233758 8900
rect 233804 8888 233832 8919
rect 234522 8916 234528 8968
rect 234580 8916 234586 8968
rect 234617 8959 234675 8965
rect 234617 8925 234629 8959
rect 234663 8956 234675 8959
rect 234798 8956 234804 8968
rect 234663 8928 234804 8956
rect 234663 8925 234675 8928
rect 234617 8919 234675 8925
rect 234632 8888 234660 8919
rect 234798 8916 234804 8928
rect 234856 8916 234862 8968
rect 235810 8916 235816 8968
rect 235868 8916 235874 8968
rect 235997 8959 236055 8965
rect 235997 8925 236009 8959
rect 236043 8925 236055 8959
rect 235997 8919 236055 8925
rect 236181 8959 236239 8965
rect 236181 8925 236193 8959
rect 236227 8956 236239 8959
rect 236641 8959 236699 8965
rect 236641 8956 236653 8959
rect 236227 8928 236653 8956
rect 236227 8925 236239 8928
rect 236181 8919 236239 8925
rect 236641 8925 236653 8928
rect 236687 8925 236699 8959
rect 236641 8919 236699 8925
rect 236012 8888 236040 8919
rect 241238 8916 241244 8968
rect 241296 8916 241302 8968
rect 241517 8959 241575 8965
rect 241517 8925 241529 8959
rect 241563 8956 241575 8959
rect 241606 8956 241612 8968
rect 241563 8928 241612 8956
rect 241563 8925 241575 8928
rect 241517 8919 241575 8925
rect 241606 8916 241612 8928
rect 241664 8916 241670 8968
rect 245010 8916 245016 8968
rect 245068 8916 245074 8968
rect 246206 8916 246212 8968
rect 246264 8916 246270 8968
rect 247126 8916 247132 8968
rect 247184 8916 247190 8968
rect 247402 8916 247408 8968
rect 247460 8916 247466 8968
rect 248690 8916 248696 8968
rect 248748 8916 248754 8968
rect 250162 8916 250168 8968
rect 250220 8916 250226 8968
rect 251174 8916 251180 8968
rect 251232 8956 251238 8968
rect 251361 8959 251419 8965
rect 251361 8956 251373 8959
rect 251232 8928 251373 8956
rect 251232 8916 251238 8928
rect 251361 8925 251373 8928
rect 251407 8925 251419 8959
rect 251361 8919 251419 8925
rect 252278 8916 252284 8968
rect 252336 8916 252342 8968
rect 253750 8916 253756 8968
rect 253808 8916 253814 8968
rect 254029 8959 254087 8965
rect 254029 8956 254041 8959
rect 253906 8928 254041 8956
rect 233752 8860 236040 8888
rect 233752 8848 233758 8860
rect 238846 8848 238852 8900
rect 238904 8888 238910 8900
rect 246942 8888 246948 8900
rect 238904 8860 246948 8888
rect 238904 8848 238910 8860
rect 246942 8848 246948 8860
rect 247000 8848 247006 8900
rect 249058 8848 249064 8900
rect 249116 8888 249122 8900
rect 253906 8888 253934 8928
rect 254029 8925 254041 8928
rect 254075 8925 254087 8959
rect 254029 8919 254087 8925
rect 255314 8916 255320 8968
rect 255372 8916 255378 8968
rect 256697 8959 256755 8965
rect 256697 8925 256709 8959
rect 256743 8956 256755 8959
rect 256786 8956 256792 8968
rect 256743 8928 256792 8956
rect 256743 8925 256755 8928
rect 256697 8919 256755 8925
rect 256786 8916 256792 8928
rect 256844 8916 256850 8968
rect 257985 8959 258043 8965
rect 257985 8925 257997 8959
rect 258031 8925 258043 8959
rect 257985 8919 258043 8925
rect 249116 8860 253934 8888
rect 249116 8848 249122 8860
rect 182140 8792 187188 8820
rect 182140 8780 182146 8792
rect 190362 8780 190368 8832
rect 190420 8820 190426 8832
rect 191101 8823 191159 8829
rect 191101 8820 191113 8823
rect 190420 8792 191113 8820
rect 190420 8780 190426 8792
rect 191101 8789 191113 8792
rect 191147 8789 191159 8823
rect 191101 8783 191159 8789
rect 191926 8780 191932 8832
rect 191984 8780 191990 8832
rect 193122 8780 193128 8832
rect 193180 8820 193186 8832
rect 193585 8823 193643 8829
rect 193585 8820 193597 8823
rect 193180 8792 193597 8820
rect 193180 8780 193186 8792
rect 193585 8789 193597 8792
rect 193631 8789 193643 8823
rect 193585 8783 193643 8789
rect 193858 8780 193864 8832
rect 193916 8820 193922 8832
rect 194965 8823 195023 8829
rect 194965 8820 194977 8823
rect 193916 8792 194977 8820
rect 193916 8780 193922 8792
rect 194965 8789 194977 8792
rect 195011 8789 195023 8823
rect 194965 8783 195023 8789
rect 195330 8780 195336 8832
rect 195388 8780 195394 8832
rect 196066 8780 196072 8832
rect 196124 8820 196130 8832
rect 196621 8823 196679 8829
rect 196621 8820 196633 8823
rect 196124 8792 196633 8820
rect 196124 8780 196130 8792
rect 196621 8789 196633 8792
rect 196667 8789 196679 8823
rect 196621 8783 196679 8789
rect 199194 8780 199200 8832
rect 199252 8820 199258 8832
rect 200117 8823 200175 8829
rect 200117 8820 200129 8823
rect 199252 8792 200129 8820
rect 199252 8780 199258 8792
rect 200117 8789 200129 8792
rect 200163 8789 200175 8823
rect 200117 8783 200175 8789
rect 200206 8780 200212 8832
rect 200264 8820 200270 8832
rect 200945 8823 201003 8829
rect 200945 8820 200957 8823
rect 200264 8792 200957 8820
rect 200264 8780 200270 8792
rect 200945 8789 200957 8792
rect 200991 8789 201003 8823
rect 200945 8783 201003 8789
rect 201034 8780 201040 8832
rect 201092 8820 201098 8832
rect 201773 8823 201831 8829
rect 201773 8820 201785 8823
rect 201092 8792 201785 8820
rect 201092 8780 201098 8792
rect 201773 8789 201785 8792
rect 201819 8789 201831 8823
rect 201773 8783 201831 8789
rect 201862 8780 201868 8832
rect 201920 8820 201926 8832
rect 202601 8823 202659 8829
rect 202601 8820 202613 8823
rect 201920 8792 202613 8820
rect 201920 8780 201926 8792
rect 202601 8789 202613 8792
rect 202647 8789 202659 8823
rect 202601 8783 202659 8789
rect 211525 8823 211583 8829
rect 211525 8789 211537 8823
rect 211571 8820 211583 8823
rect 214558 8820 214564 8832
rect 211571 8792 214564 8820
rect 211571 8789 211583 8792
rect 211525 8783 211583 8789
rect 214558 8780 214564 8792
rect 214616 8780 214622 8832
rect 216677 8823 216735 8829
rect 216677 8789 216689 8823
rect 216723 8820 216735 8823
rect 217686 8820 217692 8832
rect 216723 8792 217692 8820
rect 216723 8789 216735 8792
rect 216677 8783 216735 8789
rect 217686 8780 217692 8792
rect 217744 8780 217750 8832
rect 217962 8780 217968 8832
rect 218020 8820 218026 8832
rect 221274 8820 221280 8832
rect 218020 8792 221280 8820
rect 218020 8780 218026 8792
rect 221274 8780 221280 8792
rect 221332 8780 221338 8832
rect 221829 8823 221887 8829
rect 221829 8789 221841 8823
rect 221875 8820 221887 8823
rect 223390 8820 223396 8832
rect 221875 8792 223396 8820
rect 221875 8789 221887 8792
rect 221829 8783 221887 8789
rect 223390 8780 223396 8792
rect 223448 8780 223454 8832
rect 224494 8780 224500 8832
rect 224552 8820 224558 8832
rect 224589 8823 224647 8829
rect 224589 8820 224601 8823
rect 224552 8792 224601 8820
rect 224552 8780 224558 8792
rect 224589 8789 224601 8792
rect 224635 8789 224647 8823
rect 224589 8783 224647 8789
rect 225322 8780 225328 8832
rect 225380 8820 225386 8832
rect 225877 8823 225935 8829
rect 225877 8820 225889 8823
rect 225380 8792 225889 8820
rect 225380 8780 225386 8792
rect 225877 8789 225889 8792
rect 225923 8789 225935 8823
rect 225877 8783 225935 8789
rect 226058 8780 226064 8832
rect 226116 8820 226122 8832
rect 226705 8823 226763 8829
rect 226705 8820 226717 8823
rect 226116 8792 226717 8820
rect 226116 8780 226122 8792
rect 226705 8789 226717 8792
rect 226751 8789 226763 8823
rect 226705 8783 226763 8789
rect 226794 8780 226800 8832
rect 226852 8820 226858 8832
rect 227533 8823 227591 8829
rect 227533 8820 227545 8823
rect 226852 8792 227545 8820
rect 226852 8780 226858 8792
rect 227533 8789 227545 8792
rect 227579 8789 227591 8823
rect 227533 8783 227591 8789
rect 228082 8780 228088 8832
rect 228140 8820 228146 8832
rect 228542 8820 228548 8832
rect 228140 8792 228548 8820
rect 228140 8780 228146 8792
rect 228542 8780 228548 8792
rect 228600 8780 228606 8832
rect 229002 8780 229008 8832
rect 229060 8820 229066 8832
rect 229189 8823 229247 8829
rect 229189 8820 229201 8823
rect 229060 8792 229201 8820
rect 229060 8780 229066 8792
rect 229189 8789 229201 8792
rect 229235 8789 229247 8823
rect 230676 8820 230704 8848
rect 231302 8820 231308 8832
rect 230676 8792 231308 8820
rect 229189 8783 229247 8789
rect 231302 8780 231308 8792
rect 231360 8780 231366 8832
rect 232406 8780 232412 8832
rect 232464 8820 232470 8832
rect 233145 8823 233203 8829
rect 233145 8820 233157 8823
rect 232464 8792 233157 8820
rect 232464 8780 232470 8792
rect 233145 8789 233157 8792
rect 233191 8789 233203 8823
rect 233145 8783 233203 8789
rect 234706 8780 234712 8832
rect 234764 8820 234770 8832
rect 234801 8823 234859 8829
rect 234801 8820 234813 8823
rect 234764 8792 234813 8820
rect 234764 8780 234770 8792
rect 234801 8789 234813 8792
rect 234847 8789 234859 8823
rect 234801 8783 234859 8789
rect 245102 8780 245108 8832
rect 245160 8780 245166 8832
rect 246298 8780 246304 8832
rect 246356 8780 246362 8832
rect 247034 8780 247040 8832
rect 247092 8820 247098 8832
rect 248785 8823 248843 8829
rect 248785 8820 248797 8823
rect 247092 8792 248797 8820
rect 247092 8780 247098 8792
rect 248785 8789 248797 8792
rect 248831 8789 248843 8823
rect 248785 8783 248843 8789
rect 250254 8780 250260 8832
rect 250312 8780 250318 8832
rect 250346 8780 250352 8832
rect 250404 8820 250410 8832
rect 251453 8823 251511 8829
rect 251453 8820 251465 8823
rect 250404 8792 251465 8820
rect 250404 8780 250410 8792
rect 251453 8789 251465 8792
rect 251499 8789 251511 8823
rect 251453 8783 251511 8789
rect 251542 8780 251548 8832
rect 251600 8820 251606 8832
rect 258000 8820 258028 8919
rect 259086 8916 259092 8968
rect 259144 8916 259150 8968
rect 259178 8916 259184 8968
rect 259236 8916 259242 8968
rect 259822 8916 259828 8968
rect 259880 8916 259886 8968
rect 260009 8959 260067 8965
rect 260009 8925 260021 8959
rect 260055 8925 260067 8959
rect 260009 8919 260067 8925
rect 259196 8888 259224 8916
rect 260024 8888 260052 8919
rect 260558 8916 260564 8968
rect 260616 8956 260622 8968
rect 261680 8965 261708 8996
rect 264054 8984 264060 9036
rect 264112 9024 264118 9036
rect 265805 9027 265863 9033
rect 265805 9024 265817 9027
rect 264112 8996 265817 9024
rect 264112 8984 264118 8996
rect 265805 8993 265817 8996
rect 265851 9024 265863 9027
rect 267182 9024 267188 9036
rect 265851 8996 267188 9024
rect 265851 8993 265863 8996
rect 265805 8987 265863 8993
rect 267182 8984 267188 8996
rect 267240 8984 267246 9036
rect 267274 8984 267280 9036
rect 267332 9024 267338 9036
rect 269666 9024 269672 9036
rect 267332 8996 269672 9024
rect 267332 8984 267338 8996
rect 269666 8984 269672 8996
rect 269724 8984 269730 9036
rect 260653 8959 260711 8965
rect 260653 8956 260665 8959
rect 260616 8928 260665 8956
rect 260616 8916 260622 8928
rect 260653 8925 260665 8928
rect 260699 8925 260711 8959
rect 260653 8919 260711 8925
rect 260837 8959 260895 8965
rect 260837 8925 260849 8959
rect 260883 8925 260895 8959
rect 260837 8919 260895 8925
rect 261665 8959 261723 8965
rect 261665 8925 261677 8959
rect 261711 8956 261723 8959
rect 262309 8959 262367 8965
rect 262309 8956 262321 8959
rect 261711 8928 262321 8956
rect 261711 8925 261723 8928
rect 261665 8919 261723 8925
rect 262309 8925 262321 8928
rect 262355 8925 262367 8959
rect 262309 8919 262367 8925
rect 260852 8888 260880 8919
rect 262950 8916 262956 8968
rect 263008 8956 263014 8968
rect 263413 8959 263471 8965
rect 263413 8956 263425 8959
rect 263008 8928 263425 8956
rect 263008 8916 263014 8928
rect 263413 8925 263425 8928
rect 263459 8925 263471 8959
rect 263413 8919 263471 8925
rect 263594 8916 263600 8968
rect 263652 8916 263658 8968
rect 263870 8916 263876 8968
rect 263928 8956 263934 8968
rect 264241 8959 264299 8965
rect 264241 8956 264253 8959
rect 263928 8928 264253 8956
rect 263928 8916 263934 8928
rect 264241 8925 264253 8928
rect 264287 8925 264299 8959
rect 264241 8919 264299 8925
rect 264517 8959 264575 8965
rect 264517 8925 264529 8959
rect 264563 8956 264575 8959
rect 265250 8956 265256 8968
rect 264563 8928 265256 8956
rect 264563 8925 264575 8928
rect 264517 8919 264575 8925
rect 265250 8916 265256 8928
rect 265308 8916 265314 8968
rect 266446 8916 266452 8968
rect 266504 8956 266510 8968
rect 267737 8959 267795 8965
rect 267737 8956 267749 8959
rect 266504 8928 267749 8956
rect 266504 8916 266510 8928
rect 267737 8925 267749 8928
rect 267783 8925 267795 8959
rect 267737 8919 267795 8925
rect 267918 8916 267924 8968
rect 267976 8956 267982 8968
rect 268657 8959 268715 8965
rect 268657 8956 268669 8959
rect 267976 8928 268669 8956
rect 267976 8916 267982 8928
rect 268657 8925 268669 8928
rect 268703 8956 268715 8959
rect 269301 8959 269359 8965
rect 269301 8956 269313 8959
rect 268703 8928 269313 8956
rect 268703 8925 268715 8928
rect 268657 8919 268715 8925
rect 259196 8860 260880 8888
rect 262030 8848 262036 8900
rect 262088 8888 262094 8900
rect 262585 8891 262643 8897
rect 262585 8888 262597 8891
rect 262088 8860 262597 8888
rect 262088 8848 262094 8860
rect 262585 8857 262597 8860
rect 262631 8857 262643 8891
rect 263612 8888 263640 8916
rect 266722 8888 266728 8900
rect 263612 8860 266728 8888
rect 262585 8851 262643 8857
rect 266722 8848 266728 8860
rect 266780 8848 266786 8900
rect 266817 8891 266875 8897
rect 266817 8857 266829 8891
rect 266863 8888 266875 8891
rect 267182 8888 267188 8900
rect 266863 8860 267188 8888
rect 266863 8857 266875 8860
rect 266817 8851 266875 8857
rect 267182 8848 267188 8860
rect 267240 8848 267246 8900
rect 267366 8848 267372 8900
rect 267424 8888 267430 8900
rect 268010 8888 268016 8900
rect 267424 8860 268016 8888
rect 267424 8848 267430 8860
rect 268010 8848 268016 8860
rect 268068 8848 268074 8900
rect 269040 8832 269068 8928
rect 269301 8925 269313 8928
rect 269347 8925 269359 8959
rect 269301 8919 269359 8925
rect 270129 8891 270187 8897
rect 270129 8857 270141 8891
rect 270175 8888 270187 8891
rect 270497 8891 270555 8897
rect 270497 8888 270509 8891
rect 270175 8860 270509 8888
rect 270175 8857 270187 8860
rect 270129 8851 270187 8857
rect 270497 8857 270509 8860
rect 270543 8888 270555 8891
rect 270862 8888 270868 8900
rect 270543 8860 270868 8888
rect 270543 8857 270555 8860
rect 270497 8851 270555 8857
rect 270862 8848 270868 8860
rect 270920 8848 270926 8900
rect 251600 8792 258028 8820
rect 251600 8780 251606 8792
rect 259730 8780 259736 8832
rect 259788 8820 259794 8832
rect 260193 8823 260251 8829
rect 260193 8820 260205 8823
rect 259788 8792 260205 8820
rect 259788 8780 259794 8792
rect 260193 8789 260205 8792
rect 260239 8789 260251 8823
rect 260193 8783 260251 8789
rect 260282 8780 260288 8832
rect 260340 8820 260346 8832
rect 261021 8823 261079 8829
rect 261021 8820 261033 8823
rect 260340 8792 261033 8820
rect 260340 8780 260346 8792
rect 261021 8789 261033 8792
rect 261067 8789 261079 8823
rect 261021 8783 261079 8789
rect 263134 8780 263140 8832
rect 263192 8820 263198 8832
rect 263781 8823 263839 8829
rect 263781 8820 263793 8823
rect 263192 8792 263793 8820
rect 263192 8780 263198 8792
rect 263781 8789 263793 8792
rect 263827 8789 263839 8823
rect 263781 8783 263839 8789
rect 266173 8823 266231 8829
rect 266173 8789 266185 8823
rect 266219 8820 266231 8823
rect 266446 8820 266452 8832
rect 266219 8792 266452 8820
rect 266219 8789 266231 8792
rect 266173 8783 266231 8789
rect 266446 8780 266452 8792
rect 266504 8780 266510 8832
rect 266538 8780 266544 8832
rect 266596 8820 266602 8832
rect 266909 8823 266967 8829
rect 266909 8820 266921 8823
rect 266596 8792 266921 8820
rect 266596 8780 266602 8792
rect 266909 8789 266921 8792
rect 266955 8789 266967 8823
rect 266909 8783 266967 8789
rect 267458 8780 267464 8832
rect 267516 8820 267522 8832
rect 267829 8823 267887 8829
rect 267829 8820 267841 8823
rect 267516 8792 267841 8820
rect 267516 8780 267522 8792
rect 267829 8789 267841 8792
rect 267875 8789 267887 8823
rect 267829 8783 267887 8789
rect 269022 8780 269028 8832
rect 269080 8780 269086 8832
rect 269206 8780 269212 8832
rect 269264 8820 269270 8832
rect 270402 8820 270408 8832
rect 269264 8792 270408 8820
rect 269264 8780 269270 8792
rect 270402 8780 270408 8792
rect 270460 8780 270466 8832
rect 1104 8730 271651 8752
rect 1104 8678 68546 8730
rect 68598 8678 68610 8730
rect 68662 8678 68674 8730
rect 68726 8678 68738 8730
rect 68790 8678 68802 8730
rect 68854 8678 136143 8730
rect 136195 8678 136207 8730
rect 136259 8678 136271 8730
rect 136323 8678 136335 8730
rect 136387 8678 136399 8730
rect 136451 8678 203740 8730
rect 203792 8678 203804 8730
rect 203856 8678 203868 8730
rect 203920 8678 203932 8730
rect 203984 8678 203996 8730
rect 204048 8678 271337 8730
rect 271389 8678 271401 8730
rect 271453 8678 271465 8730
rect 271517 8678 271529 8730
rect 271581 8678 271593 8730
rect 271645 8678 271651 8730
rect 1104 8656 271651 8678
rect 10318 8576 10324 8628
rect 10376 8616 10382 8628
rect 20806 8616 20812 8628
rect 10376 8588 20812 8616
rect 10376 8576 10382 8588
rect 20806 8576 20812 8588
rect 20864 8576 20870 8628
rect 21358 8576 21364 8628
rect 21416 8576 21422 8628
rect 21450 8576 21456 8628
rect 21508 8616 21514 8628
rect 22186 8616 22192 8628
rect 21508 8588 22192 8616
rect 21508 8576 21514 8588
rect 22186 8576 22192 8588
rect 22244 8576 22250 8628
rect 24026 8576 24032 8628
rect 24084 8576 24090 8628
rect 26510 8576 26516 8628
rect 26568 8576 26574 8628
rect 27430 8576 27436 8628
rect 27488 8576 27494 8628
rect 28166 8576 28172 8628
rect 28224 8576 28230 8628
rect 28902 8576 28908 8628
rect 28960 8576 28966 8628
rect 29822 8576 29828 8628
rect 29880 8576 29886 8628
rect 31018 8576 31024 8628
rect 31076 8576 31082 8628
rect 33134 8576 33140 8628
rect 33192 8576 33198 8628
rect 53650 8576 53656 8628
rect 53708 8616 53714 8628
rect 54849 8619 54907 8625
rect 54849 8616 54861 8619
rect 53708 8588 54861 8616
rect 53708 8576 53714 8588
rect 54849 8585 54861 8588
rect 54895 8585 54907 8619
rect 54849 8579 54907 8585
rect 55858 8576 55864 8628
rect 55916 8576 55922 8628
rect 56410 8576 56416 8628
rect 56468 8616 56474 8628
rect 56597 8619 56655 8625
rect 56597 8616 56609 8619
rect 56468 8588 56609 8616
rect 56468 8576 56474 8588
rect 56597 8585 56609 8588
rect 56643 8585 56655 8619
rect 56597 8579 56655 8585
rect 57330 8576 57336 8628
rect 57388 8576 57394 8628
rect 58802 8576 58808 8628
rect 58860 8576 58866 8628
rect 59262 8576 59268 8628
rect 59320 8616 59326 8628
rect 59541 8619 59599 8625
rect 59541 8616 59553 8619
rect 59320 8588 59553 8616
rect 59320 8576 59326 8588
rect 59541 8585 59553 8588
rect 59587 8585 59599 8619
rect 59541 8579 59599 8585
rect 60274 8576 60280 8628
rect 60332 8576 60338 8628
rect 60642 8576 60648 8628
rect 60700 8616 60706 8628
rect 61657 8619 61715 8625
rect 61657 8616 61669 8619
rect 60700 8588 61669 8616
rect 60700 8576 60706 8588
rect 61657 8585 61669 8588
rect 61703 8585 61715 8619
rect 61657 8579 61715 8585
rect 62574 8576 62580 8628
rect 62632 8576 62638 8628
rect 63954 8576 63960 8628
rect 64012 8576 64018 8628
rect 64690 8576 64696 8628
rect 64748 8576 64754 8628
rect 64846 8588 80054 8616
rect 11054 8508 11060 8560
rect 11112 8548 11118 8560
rect 20714 8548 20720 8560
rect 11112 8520 20720 8548
rect 11112 8508 11118 8520
rect 20714 8508 20720 8520
rect 20772 8508 20778 8560
rect 22373 8551 22431 8557
rect 22373 8548 22385 8551
rect 22066 8520 22385 8548
rect 21177 8483 21235 8489
rect 21177 8449 21189 8483
rect 21223 8480 21235 8483
rect 22066 8480 22094 8520
rect 22373 8517 22385 8520
rect 22419 8517 22431 8551
rect 22373 8511 22431 8517
rect 23382 8508 23388 8560
rect 23440 8548 23446 8560
rect 25222 8548 25228 8560
rect 23440 8520 25228 8548
rect 23440 8508 23446 8520
rect 21223 8452 22094 8480
rect 21223 8449 21235 8452
rect 21177 8443 21235 8449
rect 22186 8440 22192 8492
rect 22244 8480 22250 8492
rect 23768 8489 23796 8520
rect 25222 8508 25228 8520
rect 25280 8508 25286 8560
rect 25682 8508 25688 8560
rect 25740 8508 25746 8560
rect 27062 8508 27068 8560
rect 27120 8548 27126 8560
rect 64846 8548 64874 8588
rect 27120 8520 57284 8548
rect 27120 8508 27126 8520
rect 22833 8483 22891 8489
rect 22833 8480 22845 8483
rect 22244 8452 22845 8480
rect 22244 8440 22250 8452
rect 22833 8449 22845 8452
rect 22879 8480 22891 8483
rect 23753 8483 23811 8489
rect 22879 8452 23612 8480
rect 22879 8449 22891 8452
rect 22833 8443 22891 8449
rect 22005 8415 22063 8421
rect 22005 8381 22017 8415
rect 22051 8412 22063 8415
rect 22278 8412 22284 8424
rect 22051 8384 22284 8412
rect 22051 8381 22063 8384
rect 22005 8375 22063 8381
rect 22278 8372 22284 8384
rect 22336 8372 22342 8424
rect 22646 8372 22652 8424
rect 22704 8372 22710 8424
rect 23106 8412 23112 8424
rect 22756 8384 23112 8412
rect 18598 8304 18604 8356
rect 18656 8344 18662 8356
rect 18656 8316 20760 8344
rect 18656 8304 18662 8316
rect 20732 8276 20760 8316
rect 21082 8304 21088 8356
rect 21140 8344 21146 8356
rect 22756 8344 22784 8384
rect 23106 8372 23112 8384
rect 23164 8372 23170 8424
rect 23584 8412 23612 8452
rect 23753 8449 23765 8483
rect 23799 8449 23811 8483
rect 23753 8443 23811 8449
rect 23845 8483 23903 8489
rect 23845 8449 23857 8483
rect 23891 8480 23903 8483
rect 24857 8483 24915 8489
rect 24857 8480 24869 8483
rect 23891 8452 24869 8480
rect 23891 8449 23903 8452
rect 23845 8443 23903 8449
rect 24857 8449 24869 8452
rect 24903 8480 24915 8483
rect 25700 8480 25728 8508
rect 24903 8452 25728 8480
rect 25869 8483 25927 8489
rect 24903 8449 24915 8452
rect 24857 8443 24915 8449
rect 25869 8449 25881 8483
rect 25915 8480 25927 8483
rect 26142 8480 26148 8492
rect 25915 8452 26148 8480
rect 25915 8449 25927 8452
rect 25869 8443 25927 8449
rect 23860 8412 23888 8443
rect 23584 8384 23888 8412
rect 24397 8415 24455 8421
rect 24397 8381 24409 8415
rect 24443 8412 24455 8415
rect 24486 8412 24492 8424
rect 24443 8384 24492 8412
rect 24443 8381 24455 8384
rect 24397 8375 24455 8381
rect 24486 8372 24492 8384
rect 24544 8412 24550 8424
rect 24673 8415 24731 8421
rect 24673 8412 24685 8415
rect 24544 8384 24685 8412
rect 24544 8372 24550 8384
rect 24673 8381 24685 8384
rect 24719 8381 24731 8415
rect 24673 8375 24731 8381
rect 25682 8372 25688 8424
rect 25740 8412 25746 8424
rect 25884 8412 25912 8443
rect 26142 8440 26148 8452
rect 26200 8440 26206 8492
rect 26329 8483 26387 8489
rect 26329 8449 26341 8483
rect 26375 8480 26387 8483
rect 27154 8480 27160 8492
rect 26375 8452 27160 8480
rect 26375 8449 26387 8452
rect 26329 8443 26387 8449
rect 27154 8440 27160 8452
rect 27212 8440 27218 8492
rect 27246 8440 27252 8492
rect 27304 8440 27310 8492
rect 27982 8440 27988 8492
rect 28040 8440 28046 8492
rect 28718 8440 28724 8492
rect 28776 8440 28782 8492
rect 29546 8440 29552 8492
rect 29604 8440 29610 8492
rect 29641 8483 29699 8489
rect 29641 8449 29653 8483
rect 29687 8449 29699 8483
rect 29641 8443 29699 8449
rect 25740 8384 25912 8412
rect 29656 8412 29684 8443
rect 30834 8440 30840 8492
rect 30892 8440 30898 8492
rect 32858 8440 32864 8492
rect 32916 8440 32922 8492
rect 32953 8483 33011 8489
rect 32953 8449 32965 8483
rect 32999 8449 33011 8483
rect 32953 8443 33011 8449
rect 31938 8412 31944 8424
rect 29656 8384 31944 8412
rect 25740 8372 25746 8384
rect 31938 8372 31944 8384
rect 31996 8412 32002 8424
rect 32968 8412 32996 8443
rect 33686 8440 33692 8492
rect 33744 8440 33750 8492
rect 54662 8440 54668 8492
rect 54720 8440 54726 8492
rect 55582 8440 55588 8492
rect 55640 8440 55646 8492
rect 55674 8440 55680 8492
rect 55732 8440 55738 8492
rect 57146 8440 57152 8492
rect 57204 8440 57210 8492
rect 33873 8415 33931 8421
rect 33873 8412 33885 8415
rect 31996 8384 33885 8412
rect 31996 8372 32002 8384
rect 33873 8381 33885 8384
rect 33919 8381 33931 8415
rect 33873 8375 33931 8381
rect 54386 8372 54392 8424
rect 54444 8412 54450 8424
rect 54481 8415 54539 8421
rect 54481 8412 54493 8415
rect 54444 8384 54493 8412
rect 54444 8372 54450 8384
rect 54481 8381 54493 8384
rect 54527 8381 54539 8415
rect 54481 8375 54539 8381
rect 56410 8372 56416 8424
rect 56468 8412 56474 8424
rect 56965 8415 57023 8421
rect 56965 8412 56977 8415
rect 56468 8384 56977 8412
rect 56468 8372 56474 8384
rect 56965 8381 56977 8384
rect 57011 8381 57023 8415
rect 57256 8412 57284 8520
rect 57440 8520 64874 8548
rect 57330 8440 57336 8492
rect 57388 8480 57394 8492
rect 57440 8480 57468 8520
rect 65978 8508 65984 8560
rect 66036 8548 66042 8560
rect 67082 8548 67088 8560
rect 66036 8520 67088 8548
rect 66036 8508 66042 8520
rect 67082 8508 67088 8520
rect 67140 8548 67146 8560
rect 80026 8548 80054 8588
rect 87506 8576 87512 8628
rect 87564 8616 87570 8628
rect 88981 8619 89039 8625
rect 88981 8616 88993 8619
rect 87564 8588 88993 8616
rect 87564 8576 87570 8588
rect 88981 8585 88993 8588
rect 89027 8585 89039 8619
rect 88981 8579 89039 8585
rect 90818 8576 90824 8628
rect 90876 8576 90882 8628
rect 91554 8576 91560 8628
rect 91612 8616 91618 8628
rect 91925 8619 91983 8625
rect 91925 8616 91937 8619
rect 91612 8588 91937 8616
rect 91612 8576 91618 8588
rect 91925 8585 91937 8588
rect 91971 8585 91983 8619
rect 91925 8579 91983 8585
rect 92566 8576 92572 8628
rect 92624 8616 92630 8628
rect 93397 8619 93455 8625
rect 93397 8616 93409 8619
rect 92624 8588 93409 8616
rect 92624 8576 92630 8588
rect 93397 8585 93409 8588
rect 93443 8585 93455 8619
rect 93397 8579 93455 8585
rect 94590 8576 94596 8628
rect 94648 8576 94654 8628
rect 95050 8576 95056 8628
rect 95108 8576 95114 8628
rect 95418 8576 95424 8628
rect 95476 8576 95482 8628
rect 96154 8576 96160 8628
rect 96212 8576 96218 8628
rect 96890 8576 96896 8628
rect 96948 8576 96954 8628
rect 97258 8576 97264 8628
rect 97316 8616 97322 8628
rect 97316 8588 97396 8616
rect 97316 8576 97322 8588
rect 89349 8551 89407 8557
rect 89349 8548 89361 8551
rect 67140 8520 67312 8548
rect 80026 8520 89361 8548
rect 67140 8508 67146 8520
rect 57388 8452 57468 8480
rect 57388 8440 57394 8452
rect 58250 8440 58256 8492
rect 58308 8480 58314 8492
rect 58621 8483 58679 8489
rect 58621 8480 58633 8483
rect 58308 8452 58633 8480
rect 58308 8440 58314 8452
rect 58621 8449 58633 8452
rect 58667 8449 58679 8483
rect 58621 8443 58679 8449
rect 59354 8440 59360 8492
rect 59412 8440 59418 8492
rect 60090 8440 60096 8492
rect 60148 8440 60154 8492
rect 60826 8440 60832 8492
rect 60884 8440 60890 8492
rect 62022 8440 62028 8492
rect 62080 8480 62086 8492
rect 62209 8483 62267 8489
rect 62209 8480 62221 8483
rect 62080 8452 62221 8480
rect 62080 8440 62086 8452
rect 62209 8449 62221 8452
rect 62255 8449 62267 8483
rect 62209 8443 62267 8449
rect 62393 8483 62451 8489
rect 62393 8449 62405 8483
rect 62439 8480 62451 8483
rect 62482 8480 62488 8492
rect 62439 8452 62488 8480
rect 62439 8449 62451 8452
rect 62393 8443 62451 8449
rect 62482 8440 62488 8452
rect 62540 8440 62546 8492
rect 63770 8440 63776 8492
rect 63828 8440 63834 8492
rect 64506 8440 64512 8492
rect 64564 8440 64570 8492
rect 65334 8440 65340 8492
rect 65392 8440 65398 8492
rect 66070 8440 66076 8492
rect 66128 8440 66134 8492
rect 67284 8489 67312 8520
rect 89349 8517 89361 8520
rect 89395 8548 89407 8551
rect 89622 8548 89628 8560
rect 89395 8520 89628 8548
rect 89395 8517 89407 8520
rect 89349 8511 89407 8517
rect 89622 8508 89628 8520
rect 89680 8548 89686 8560
rect 97166 8548 97172 8560
rect 89680 8520 89760 8548
rect 89680 8508 89686 8520
rect 67269 8483 67327 8489
rect 67269 8449 67281 8483
rect 67315 8449 67327 8483
rect 67269 8443 67327 8449
rect 74258 8440 74264 8492
rect 74316 8440 74322 8492
rect 74534 8440 74540 8492
rect 74592 8440 74598 8492
rect 76466 8440 76472 8492
rect 76524 8440 76530 8492
rect 88794 8440 88800 8492
rect 88852 8440 88858 8492
rect 89732 8489 89760 8520
rect 93596 8520 97172 8548
rect 89717 8483 89775 8489
rect 89717 8449 89729 8483
rect 89763 8449 89775 8483
rect 89717 8443 89775 8449
rect 89901 8483 89959 8489
rect 89901 8449 89913 8483
rect 89947 8480 89959 8483
rect 89990 8480 89996 8492
rect 89947 8452 89996 8480
rect 89947 8449 89959 8452
rect 89901 8443 89959 8449
rect 89990 8440 89996 8452
rect 90048 8440 90054 8492
rect 90634 8440 90640 8492
rect 90692 8440 90698 8492
rect 91002 8440 91008 8492
rect 91060 8480 91066 8492
rect 91281 8483 91339 8489
rect 91281 8480 91293 8483
rect 91060 8452 91293 8480
rect 91060 8440 91066 8452
rect 91281 8449 91293 8452
rect 91327 8480 91339 8483
rect 91557 8483 91615 8489
rect 91557 8480 91569 8483
rect 91327 8452 91569 8480
rect 91327 8449 91339 8452
rect 91281 8443 91339 8449
rect 91557 8449 91569 8452
rect 91603 8449 91615 8483
rect 91557 8443 91615 8449
rect 91741 8483 91799 8489
rect 91741 8449 91753 8483
rect 91787 8480 91799 8483
rect 93213 8483 93271 8489
rect 93213 8480 93225 8483
rect 91787 8452 93225 8480
rect 91787 8449 91799 8452
rect 91741 8443 91799 8449
rect 93213 8449 93225 8452
rect 93259 8480 93271 8483
rect 93486 8480 93492 8492
rect 93259 8452 93492 8480
rect 93259 8449 93271 8452
rect 93213 8443 93271 8449
rect 93486 8440 93492 8452
rect 93544 8440 93550 8492
rect 61286 8412 61292 8424
rect 57256 8384 61292 8412
rect 56965 8375 57023 8381
rect 61286 8372 61292 8384
rect 61344 8412 61350 8424
rect 61470 8412 61476 8424
rect 61344 8384 61476 8412
rect 61344 8372 61350 8384
rect 61470 8372 61476 8384
rect 61528 8372 61534 8424
rect 66993 8415 67051 8421
rect 66993 8381 67005 8415
rect 67039 8412 67051 8415
rect 67358 8412 67364 8424
rect 67039 8384 67364 8412
rect 67039 8381 67051 8384
rect 66993 8375 67051 8381
rect 67358 8372 67364 8384
rect 67416 8372 67422 8424
rect 76745 8415 76803 8421
rect 76745 8381 76757 8415
rect 76791 8412 76803 8415
rect 82722 8412 82728 8424
rect 76791 8384 82728 8412
rect 76791 8381 76803 8384
rect 76745 8375 76803 8381
rect 82722 8372 82728 8384
rect 82780 8372 82786 8424
rect 84838 8372 84844 8424
rect 84896 8412 84902 8424
rect 92934 8412 92940 8424
rect 84896 8384 92940 8412
rect 84896 8372 84902 8384
rect 92934 8372 92940 8384
rect 92992 8372 92998 8424
rect 93026 8372 93032 8424
rect 93084 8372 93090 8424
rect 21140 8316 22784 8344
rect 23017 8347 23075 8353
rect 21140 8304 21146 8316
rect 23017 8313 23029 8347
rect 23063 8344 23075 8347
rect 23474 8344 23480 8356
rect 23063 8316 23480 8344
rect 23063 8313 23075 8316
rect 23017 8307 23075 8313
rect 23474 8304 23480 8316
rect 23532 8304 23538 8356
rect 24228 8316 24440 8344
rect 24228 8276 24256 8316
rect 20732 8248 24256 8276
rect 24412 8276 24440 8316
rect 24964 8316 25176 8344
rect 24964 8276 24992 8316
rect 24412 8248 24992 8276
rect 25038 8236 25044 8288
rect 25096 8236 25102 8288
rect 25148 8276 25176 8316
rect 25700 8316 25912 8344
rect 25700 8276 25728 8316
rect 25148 8248 25728 8276
rect 25884 8276 25912 8316
rect 28534 8304 28540 8356
rect 28592 8344 28598 8356
rect 32950 8344 32956 8356
rect 28592 8316 32956 8344
rect 28592 8304 28598 8316
rect 32950 8304 32956 8316
rect 33008 8304 33014 8356
rect 33060 8316 33916 8344
rect 33060 8276 33088 8316
rect 25884 8248 33088 8276
rect 33888 8276 33916 8316
rect 54110 8304 54116 8356
rect 54168 8344 54174 8356
rect 57330 8344 57336 8356
rect 54168 8316 57336 8344
rect 54168 8304 54174 8316
rect 57330 8304 57336 8316
rect 57388 8304 57394 8356
rect 57422 8304 57428 8356
rect 57480 8344 57486 8356
rect 62666 8344 62672 8356
rect 57480 8316 62672 8344
rect 57480 8304 57486 8316
rect 62666 8304 62672 8316
rect 62724 8304 62730 8356
rect 65518 8304 65524 8356
rect 65576 8304 65582 8356
rect 65886 8304 65892 8356
rect 65944 8344 65950 8356
rect 66257 8347 66315 8353
rect 66257 8344 66269 8347
rect 65944 8316 66269 8344
rect 65944 8304 65950 8316
rect 66257 8313 66269 8316
rect 66303 8313 66315 8347
rect 93596 8344 93624 8520
rect 97166 8508 97172 8520
rect 97224 8508 97230 8560
rect 94406 8440 94412 8492
rect 94464 8440 94470 8492
rect 94866 8440 94872 8492
rect 94924 8440 94930 8492
rect 95050 8440 95056 8492
rect 95108 8480 95114 8492
rect 95418 8480 95424 8492
rect 95108 8452 95424 8480
rect 95108 8440 95114 8452
rect 95418 8440 95424 8452
rect 95476 8480 95482 8492
rect 95694 8480 95700 8492
rect 95476 8452 95700 8480
rect 95476 8440 95482 8452
rect 95694 8440 95700 8452
rect 95752 8478 95758 8492
rect 95789 8483 95847 8489
rect 95789 8478 95801 8483
rect 95752 8450 95801 8478
rect 95752 8440 95758 8450
rect 95789 8449 95801 8450
rect 95835 8449 95847 8483
rect 95789 8443 95847 8449
rect 95878 8440 95884 8492
rect 95936 8480 95942 8492
rect 95973 8483 96031 8489
rect 95973 8480 95985 8483
rect 95936 8452 95985 8480
rect 95936 8440 95942 8452
rect 95973 8449 95985 8452
rect 96019 8480 96031 8483
rect 96709 8483 96767 8489
rect 96709 8480 96721 8483
rect 96019 8452 96721 8480
rect 96019 8449 96031 8452
rect 95973 8443 96031 8449
rect 96709 8449 96721 8452
rect 96755 8480 96767 8483
rect 97258 8480 97264 8492
rect 96755 8452 97264 8480
rect 96755 8449 96767 8452
rect 96709 8443 96767 8449
rect 97258 8440 97264 8452
rect 97316 8440 97322 8492
rect 97368 8489 97396 8588
rect 97534 8576 97540 8628
rect 97592 8576 97598 8628
rect 97994 8576 98000 8628
rect 98052 8616 98058 8628
rect 98273 8619 98331 8625
rect 98273 8616 98285 8619
rect 98052 8588 98285 8616
rect 98052 8576 98058 8588
rect 98273 8585 98285 8588
rect 98319 8585 98331 8619
rect 98273 8579 98331 8585
rect 99374 8576 99380 8628
rect 99432 8616 99438 8628
rect 99837 8619 99895 8625
rect 99837 8616 99849 8619
rect 99432 8588 99849 8616
rect 99432 8576 99438 8588
rect 99837 8585 99849 8588
rect 99883 8585 99895 8619
rect 121546 8616 121552 8628
rect 99837 8579 99895 8585
rect 99944 8588 121552 8616
rect 99466 8508 99472 8560
rect 99524 8548 99530 8560
rect 99944 8548 99972 8588
rect 121546 8576 121552 8588
rect 121604 8576 121610 8628
rect 121638 8576 121644 8628
rect 121696 8576 121702 8628
rect 122374 8576 122380 8628
rect 122432 8576 122438 8628
rect 123202 8576 123208 8628
rect 123260 8576 123266 8628
rect 124030 8576 124036 8628
rect 124088 8576 124094 8628
rect 125594 8576 125600 8628
rect 125652 8576 125658 8628
rect 126974 8576 126980 8628
rect 127032 8576 127038 8628
rect 127710 8576 127716 8628
rect 127768 8576 127774 8628
rect 128262 8576 128268 8628
rect 128320 8576 128326 8628
rect 129366 8576 129372 8628
rect 129424 8616 129430 8628
rect 130565 8619 130623 8625
rect 130565 8616 130577 8619
rect 129424 8588 130577 8616
rect 129424 8576 129430 8588
rect 130565 8585 130577 8588
rect 130611 8585 130623 8619
rect 130565 8579 130623 8585
rect 132126 8576 132132 8628
rect 132184 8576 132190 8628
rect 134518 8576 134524 8628
rect 134576 8576 134582 8628
rect 137186 8576 137192 8628
rect 137244 8616 137250 8628
rect 153838 8616 153844 8628
rect 137244 8588 153844 8616
rect 137244 8576 137250 8588
rect 153838 8576 153844 8588
rect 153896 8576 153902 8628
rect 156046 8576 156052 8628
rect 156104 8616 156110 8628
rect 156141 8619 156199 8625
rect 156141 8616 156153 8619
rect 156104 8588 156153 8616
rect 156104 8576 156110 8588
rect 156141 8585 156153 8588
rect 156187 8585 156199 8619
rect 156141 8579 156199 8585
rect 156230 8576 156236 8628
rect 156288 8616 156294 8628
rect 161842 8616 161848 8628
rect 156288 8588 161848 8616
rect 156288 8576 156294 8588
rect 161842 8576 161848 8588
rect 161900 8576 161906 8628
rect 161934 8576 161940 8628
rect 161992 8616 161998 8628
rect 161992 8588 214052 8616
rect 161992 8576 161998 8588
rect 99524 8520 99972 8548
rect 99524 8508 99530 8520
rect 100294 8508 100300 8560
rect 100352 8548 100358 8560
rect 123386 8548 123392 8560
rect 100352 8520 123392 8548
rect 100352 8508 100358 8520
rect 123386 8508 123392 8520
rect 123444 8508 123450 8560
rect 127802 8508 127808 8560
rect 127860 8548 127866 8560
rect 127860 8520 134380 8548
rect 127860 8508 127866 8520
rect 97353 8483 97411 8489
rect 97353 8449 97365 8483
rect 97399 8449 97411 8483
rect 97353 8443 97411 8449
rect 98086 8440 98092 8492
rect 98144 8440 98150 8492
rect 99650 8440 99656 8492
rect 99708 8440 99714 8492
rect 102042 8440 102048 8492
rect 102100 8480 102106 8492
rect 121457 8483 121515 8489
rect 102100 8452 121408 8480
rect 102100 8440 102106 8452
rect 96430 8372 96436 8424
rect 96488 8412 96494 8424
rect 96525 8415 96583 8421
rect 96525 8412 96537 8415
rect 96488 8384 96537 8412
rect 96488 8372 96494 8384
rect 96525 8381 96537 8384
rect 96571 8381 96583 8415
rect 96525 8375 96583 8381
rect 96614 8372 96620 8424
rect 96672 8412 96678 8424
rect 97994 8412 98000 8424
rect 96672 8384 98000 8412
rect 96672 8372 96678 8384
rect 97994 8372 98000 8384
rect 98052 8372 98058 8424
rect 100665 8415 100723 8421
rect 98114 8384 100064 8412
rect 66257 8307 66315 8313
rect 86926 8316 93624 8344
rect 95344 8316 95556 8344
rect 51166 8276 51172 8288
rect 33888 8248 51172 8276
rect 51166 8236 51172 8248
rect 51224 8236 51230 8288
rect 61010 8236 61016 8288
rect 61068 8236 61074 8288
rect 70394 8236 70400 8288
rect 70452 8276 70458 8288
rect 86926 8276 86954 8316
rect 70452 8248 86954 8276
rect 70452 8236 70458 8248
rect 90082 8236 90088 8288
rect 90140 8236 90146 8288
rect 93210 8236 93216 8288
rect 93268 8276 93274 8288
rect 95344 8276 95372 8316
rect 93268 8248 95372 8276
rect 95528 8276 95556 8316
rect 95694 8304 95700 8356
rect 95752 8344 95758 8356
rect 98114 8344 98142 8384
rect 100036 8344 100064 8384
rect 100665 8381 100677 8415
rect 100711 8412 100723 8415
rect 100754 8412 100760 8424
rect 100711 8384 100760 8412
rect 100711 8381 100723 8384
rect 100665 8375 100723 8381
rect 100754 8372 100760 8384
rect 100812 8372 100818 8424
rect 100938 8372 100944 8424
rect 100996 8372 101002 8424
rect 101950 8372 101956 8424
rect 102008 8372 102014 8424
rect 120810 8372 120816 8424
rect 120868 8412 120874 8424
rect 121273 8415 121331 8421
rect 121273 8412 121285 8415
rect 120868 8384 121285 8412
rect 120868 8372 120874 8384
rect 121273 8381 121285 8384
rect 121319 8381 121331 8415
rect 121380 8412 121408 8452
rect 121457 8449 121469 8483
rect 121503 8480 121515 8483
rect 121822 8480 121828 8492
rect 121503 8452 121828 8480
rect 121503 8449 121515 8452
rect 121457 8443 121515 8449
rect 121822 8440 121828 8452
rect 121880 8440 121886 8492
rect 122190 8440 122196 8492
rect 122248 8440 122254 8492
rect 123018 8440 123024 8492
rect 123076 8440 123082 8492
rect 123846 8440 123852 8492
rect 123904 8440 123910 8492
rect 125410 8440 125416 8492
rect 125468 8440 125474 8492
rect 126790 8440 126796 8492
rect 126848 8440 126854 8492
rect 127526 8440 127532 8492
rect 127584 8440 127590 8492
rect 128078 8440 128084 8492
rect 128136 8440 128142 8492
rect 128814 8440 128820 8492
rect 128872 8480 128878 8492
rect 129185 8483 129243 8489
rect 129185 8480 129197 8483
rect 128872 8452 129197 8480
rect 128872 8440 128878 8452
rect 129185 8449 129197 8452
rect 129231 8480 129243 8483
rect 130381 8483 130439 8489
rect 130381 8480 130393 8483
rect 129231 8452 130393 8480
rect 129231 8449 129243 8452
rect 129185 8443 129243 8449
rect 130381 8449 130393 8452
rect 130427 8449 130439 8483
rect 130381 8443 130439 8449
rect 131942 8440 131948 8492
rect 132000 8440 132006 8492
rect 132862 8440 132868 8492
rect 132920 8440 132926 8492
rect 134242 8440 134248 8492
rect 134300 8440 134306 8492
rect 134352 8489 134380 8520
rect 135530 8508 135536 8560
rect 135588 8548 135594 8560
rect 135588 8520 138014 8548
rect 135588 8508 135594 8520
rect 134337 8483 134395 8489
rect 134337 8449 134349 8483
rect 134383 8449 134395 8483
rect 137986 8480 138014 8520
rect 143718 8508 143724 8560
rect 143776 8548 143782 8560
rect 152458 8548 152464 8560
rect 143776 8520 152464 8548
rect 143776 8508 143782 8520
rect 152458 8508 152464 8520
rect 152516 8508 152522 8560
rect 154022 8508 154028 8560
rect 154080 8548 154086 8560
rect 156506 8548 156512 8560
rect 154080 8520 156512 8548
rect 154080 8508 154086 8520
rect 156506 8508 156512 8520
rect 156564 8508 156570 8560
rect 171870 8548 171876 8560
rect 158916 8520 171876 8548
rect 153746 8480 153752 8492
rect 137986 8452 153752 8480
rect 134337 8443 134395 8449
rect 153746 8440 153752 8452
rect 153804 8440 153810 8492
rect 155954 8440 155960 8492
rect 156012 8440 156018 8492
rect 158916 8489 158944 8520
rect 171870 8508 171876 8520
rect 171928 8508 171934 8560
rect 213914 8548 213920 8560
rect 180766 8520 213920 8548
rect 156877 8483 156935 8489
rect 156877 8449 156889 8483
rect 156923 8480 156935 8483
rect 157981 8483 158039 8489
rect 157981 8480 157993 8483
rect 156923 8452 157993 8480
rect 156923 8449 156935 8452
rect 156877 8443 156935 8449
rect 157981 8449 157993 8452
rect 158027 8449 158039 8483
rect 157981 8443 158039 8449
rect 158533 8483 158591 8489
rect 158533 8449 158545 8483
rect 158579 8480 158591 8483
rect 158901 8483 158959 8489
rect 158901 8480 158913 8483
rect 158579 8452 158913 8480
rect 158579 8449 158591 8452
rect 158533 8443 158591 8449
rect 158901 8449 158913 8452
rect 158947 8449 158959 8483
rect 160189 8483 160247 8489
rect 160189 8480 160201 8483
rect 158901 8443 158959 8449
rect 159008 8452 160201 8480
rect 128633 8415 128691 8421
rect 128633 8412 128645 8415
rect 121380 8384 128645 8412
rect 121273 8375 121331 8381
rect 128633 8381 128645 8384
rect 128679 8412 128691 8415
rect 128906 8412 128912 8424
rect 128679 8384 128912 8412
rect 128679 8381 128691 8384
rect 128633 8375 128691 8381
rect 128906 8372 128912 8384
rect 128964 8412 128970 8424
rect 129001 8415 129059 8421
rect 129001 8412 129013 8415
rect 128964 8384 129013 8412
rect 128964 8372 128970 8384
rect 129001 8381 129013 8384
rect 129047 8381 129059 8415
rect 129001 8375 129059 8381
rect 113818 8344 113824 8356
rect 95752 8316 98142 8344
rect 99760 8316 99972 8344
rect 100036 8316 113824 8344
rect 95752 8304 95758 8316
rect 99760 8276 99788 8316
rect 95528 8248 99788 8276
rect 99944 8276 99972 8316
rect 113818 8304 113824 8316
rect 113876 8304 113882 8356
rect 129016 8344 129044 8375
rect 130194 8372 130200 8424
rect 130252 8412 130258 8424
rect 130838 8412 130844 8424
rect 130252 8384 130844 8412
rect 130252 8372 130258 8384
rect 130838 8372 130844 8384
rect 130896 8372 130902 8424
rect 132678 8372 132684 8424
rect 132736 8412 132742 8424
rect 142798 8412 142804 8424
rect 132736 8384 142804 8412
rect 132736 8372 132742 8384
rect 142798 8372 142804 8384
rect 142856 8372 142862 8424
rect 148778 8372 148784 8424
rect 148836 8412 148842 8424
rect 156138 8412 156144 8424
rect 148836 8384 156144 8412
rect 148836 8372 148842 8384
rect 156138 8372 156144 8384
rect 156196 8372 156202 8424
rect 156230 8372 156236 8424
rect 156288 8412 156294 8424
rect 156693 8415 156751 8421
rect 156693 8412 156705 8415
rect 156288 8384 156705 8412
rect 156288 8372 156294 8384
rect 156693 8381 156705 8384
rect 156739 8381 156751 8415
rect 156693 8375 156751 8381
rect 157794 8372 157800 8424
rect 157852 8372 157858 8424
rect 157996 8412 158024 8443
rect 159008 8412 159036 8452
rect 160189 8449 160201 8452
rect 160235 8480 160247 8483
rect 161201 8483 161259 8489
rect 161201 8480 161213 8483
rect 160235 8452 161213 8480
rect 160235 8449 160247 8452
rect 160189 8443 160247 8449
rect 161201 8449 161213 8452
rect 161247 8480 161259 8483
rect 161290 8480 161296 8492
rect 161247 8452 161296 8480
rect 161247 8449 161259 8452
rect 161201 8443 161259 8449
rect 161290 8440 161296 8452
rect 161348 8440 161354 8492
rect 161753 8483 161811 8489
rect 161753 8449 161765 8483
rect 161799 8480 161811 8483
rect 162118 8480 162124 8492
rect 161799 8452 162124 8480
rect 161799 8449 161811 8452
rect 161753 8443 161811 8449
rect 162118 8440 162124 8452
rect 162176 8440 162182 8492
rect 163317 8483 163375 8489
rect 163317 8449 163329 8483
rect 163363 8480 163375 8483
rect 163685 8483 163743 8489
rect 163685 8480 163697 8483
rect 163363 8452 163697 8480
rect 163363 8449 163375 8452
rect 163317 8443 163375 8449
rect 163685 8449 163697 8452
rect 163731 8480 163743 8483
rect 163866 8480 163872 8492
rect 163731 8452 163872 8480
rect 163731 8449 163743 8452
rect 163685 8443 163743 8449
rect 163866 8440 163872 8452
rect 163924 8440 163930 8492
rect 164697 8483 164755 8489
rect 164697 8449 164709 8483
rect 164743 8480 164755 8483
rect 165062 8480 165068 8492
rect 164743 8452 165068 8480
rect 164743 8449 164755 8452
rect 164697 8443 164755 8449
rect 165062 8440 165068 8452
rect 165120 8440 165126 8492
rect 166350 8440 166356 8492
rect 166408 8440 166414 8492
rect 166445 8483 166503 8489
rect 166445 8449 166457 8483
rect 166491 8480 166503 8483
rect 166534 8480 166540 8492
rect 166491 8452 166540 8480
rect 166491 8449 166503 8452
rect 166445 8443 166503 8449
rect 166534 8440 166540 8452
rect 166592 8480 166598 8492
rect 166810 8480 166816 8492
rect 166592 8452 166816 8480
rect 166592 8440 166598 8452
rect 166810 8440 166816 8452
rect 166868 8440 166874 8492
rect 166902 8440 166908 8492
rect 166960 8440 166966 8492
rect 166997 8483 167055 8489
rect 166997 8449 167009 8483
rect 167043 8480 167055 8483
rect 167365 8483 167423 8489
rect 167365 8480 167377 8483
rect 167043 8452 167377 8480
rect 167043 8449 167055 8452
rect 166997 8443 167055 8449
rect 167365 8449 167377 8452
rect 167411 8480 167423 8483
rect 180766 8480 180794 8520
rect 213914 8508 213920 8520
rect 213972 8508 213978 8560
rect 167411 8452 180794 8480
rect 167411 8449 167423 8452
rect 167365 8443 167423 8449
rect 186958 8440 186964 8492
rect 187016 8440 187022 8492
rect 190362 8440 190368 8492
rect 190420 8440 190426 8492
rect 191101 8483 191159 8489
rect 191101 8449 191113 8483
rect 191147 8480 191159 8483
rect 191926 8480 191932 8492
rect 191147 8452 191932 8480
rect 191147 8449 191159 8452
rect 191101 8443 191159 8449
rect 191926 8440 191932 8452
rect 191984 8440 191990 8492
rect 192386 8440 192392 8492
rect 192444 8440 192450 8492
rect 192478 8440 192484 8492
rect 192536 8440 192542 8492
rect 192662 8440 192668 8492
rect 192720 8440 192726 8492
rect 193122 8440 193128 8492
rect 193180 8440 193186 8492
rect 193858 8440 193864 8492
rect 193916 8440 193922 8492
rect 195425 8483 195483 8489
rect 195425 8449 195437 8483
rect 195471 8449 195483 8483
rect 195425 8443 195483 8449
rect 157996 8384 159036 8412
rect 159453 8415 159511 8421
rect 159453 8381 159465 8415
rect 159499 8412 159511 8415
rect 159542 8412 159548 8424
rect 159499 8384 159548 8412
rect 159499 8381 159511 8384
rect 159453 8375 159511 8381
rect 159542 8372 159548 8384
rect 159600 8372 159606 8424
rect 159910 8372 159916 8424
rect 159968 8412 159974 8424
rect 160005 8415 160063 8421
rect 160005 8412 160017 8415
rect 159968 8384 160017 8412
rect 159968 8372 159974 8384
rect 160005 8381 160017 8384
rect 160051 8381 160063 8415
rect 160005 8375 160063 8381
rect 161017 8415 161075 8421
rect 161017 8381 161029 8415
rect 161063 8412 161075 8415
rect 161106 8412 161112 8424
rect 161063 8384 161112 8412
rect 161063 8381 161075 8384
rect 161017 8375 161075 8381
rect 161106 8372 161112 8384
rect 161164 8372 161170 8424
rect 161658 8372 161664 8424
rect 161716 8412 161722 8424
rect 162302 8412 162308 8424
rect 161716 8384 162308 8412
rect 161716 8372 161722 8384
rect 162302 8372 162308 8384
rect 162360 8372 162366 8424
rect 162670 8372 162676 8424
rect 162728 8372 162734 8424
rect 163590 8372 163596 8424
rect 163648 8412 163654 8424
rect 163961 8415 164019 8421
rect 163961 8412 163973 8415
rect 163648 8384 163973 8412
rect 163648 8372 163654 8384
rect 163961 8381 163973 8384
rect 164007 8381 164019 8415
rect 165338 8412 165344 8424
rect 163961 8375 164019 8381
rect 165080 8384 165344 8412
rect 129016 8316 147674 8344
rect 111518 8276 111524 8288
rect 99944 8248 111524 8276
rect 93268 8236 93274 8248
rect 111518 8236 111524 8248
rect 111576 8236 111582 8288
rect 129090 8236 129096 8288
rect 129148 8276 129154 8288
rect 129369 8279 129427 8285
rect 129369 8276 129381 8279
rect 129148 8248 129381 8276
rect 129148 8236 129154 8248
rect 129369 8245 129381 8248
rect 129415 8245 129427 8279
rect 129369 8239 129427 8245
rect 132770 8236 132776 8288
rect 132828 8276 132834 8288
rect 133049 8279 133107 8285
rect 133049 8276 133061 8279
rect 132828 8248 133061 8276
rect 132828 8236 132834 8248
rect 133049 8245 133061 8248
rect 133095 8245 133107 8279
rect 147646 8276 147674 8316
rect 151446 8304 151452 8356
rect 151504 8344 151510 8356
rect 154022 8344 154028 8356
rect 151504 8316 154028 8344
rect 151504 8304 151510 8316
rect 154022 8304 154028 8316
rect 154080 8304 154086 8356
rect 154666 8304 154672 8356
rect 154724 8344 154730 8356
rect 157812 8344 157840 8372
rect 165080 8356 165108 8384
rect 165338 8372 165344 8384
rect 165396 8372 165402 8424
rect 166920 8412 166948 8440
rect 167641 8415 167699 8421
rect 167641 8412 167653 8415
rect 166920 8384 167653 8412
rect 167641 8381 167653 8384
rect 167687 8381 167699 8415
rect 167641 8375 167699 8381
rect 168650 8372 168656 8424
rect 168708 8372 168714 8424
rect 168926 8372 168932 8424
rect 168984 8372 168990 8424
rect 169754 8372 169760 8424
rect 169812 8412 169818 8424
rect 169941 8415 169999 8421
rect 169941 8412 169953 8415
rect 169812 8384 169953 8412
rect 169812 8372 169818 8384
rect 169941 8381 169953 8384
rect 169987 8381 169999 8415
rect 187237 8415 187295 8421
rect 187237 8412 187249 8415
rect 169941 8375 169999 8381
rect 180766 8384 187249 8412
rect 154724 8316 157840 8344
rect 158165 8347 158223 8353
rect 154724 8304 154730 8316
rect 158165 8313 158177 8347
rect 158211 8344 158223 8347
rect 159266 8344 159272 8356
rect 158211 8316 159272 8344
rect 158211 8313 158223 8316
rect 158165 8307 158223 8313
rect 159266 8304 159272 8316
rect 159324 8304 159330 8356
rect 161385 8347 161443 8353
rect 161385 8313 161397 8347
rect 161431 8344 161443 8347
rect 161474 8344 161480 8356
rect 161431 8316 161480 8344
rect 161431 8313 161443 8316
rect 161385 8307 161443 8313
rect 161474 8304 161480 8316
rect 161532 8304 161538 8356
rect 165062 8304 165068 8356
rect 165120 8304 165126 8356
rect 166552 8316 167132 8344
rect 151722 8276 151728 8288
rect 147646 8248 151728 8276
rect 133049 8239 133107 8245
rect 151722 8236 151728 8248
rect 151780 8236 151786 8288
rect 157058 8236 157064 8288
rect 157116 8236 157122 8288
rect 160373 8279 160431 8285
rect 160373 8245 160385 8279
rect 160419 8276 160431 8279
rect 160738 8276 160744 8288
rect 160419 8248 160744 8276
rect 160419 8245 160431 8248
rect 160373 8239 160431 8245
rect 160738 8236 160744 8248
rect 160796 8236 160802 8288
rect 161934 8236 161940 8288
rect 161992 8276 161998 8288
rect 164234 8276 164240 8288
rect 161992 8248 164240 8276
rect 161992 8236 161998 8248
rect 164234 8236 164240 8248
rect 164292 8236 164298 8288
rect 164694 8236 164700 8288
rect 164752 8276 164758 8288
rect 166552 8276 166580 8316
rect 164752 8248 166580 8276
rect 164752 8236 164758 8248
rect 166626 8236 166632 8288
rect 166684 8236 166690 8288
rect 167104 8276 167132 8316
rect 168834 8304 168840 8356
rect 168892 8344 168898 8356
rect 169662 8344 169668 8356
rect 168892 8316 169668 8344
rect 168892 8304 168898 8316
rect 169662 8304 169668 8316
rect 169720 8304 169726 8356
rect 180766 8276 180794 8384
rect 187237 8381 187249 8384
rect 187283 8381 187295 8415
rect 187237 8375 187295 8381
rect 195241 8415 195299 8421
rect 195241 8381 195253 8415
rect 195287 8381 195299 8415
rect 195440 8412 195468 8443
rect 195606 8440 195612 8492
rect 195664 8440 195670 8492
rect 196066 8440 196072 8492
rect 196124 8440 196130 8492
rect 197357 8483 197415 8489
rect 197357 8480 197369 8483
rect 196268 8452 197369 8480
rect 195974 8412 195980 8424
rect 195440 8384 195980 8412
rect 195241 8375 195299 8381
rect 189902 8304 189908 8356
rect 189960 8344 189966 8356
rect 190549 8347 190607 8353
rect 190549 8344 190561 8347
rect 189960 8316 190561 8344
rect 189960 8304 189966 8316
rect 190549 8313 190561 8316
rect 190595 8313 190607 8347
rect 190549 8307 190607 8313
rect 191282 8304 191288 8356
rect 191340 8304 191346 8356
rect 192846 8304 192852 8356
rect 192904 8344 192910 8356
rect 193309 8347 193367 8353
rect 193309 8344 193321 8347
rect 192904 8316 193321 8344
rect 192904 8304 192910 8316
rect 193309 8313 193321 8316
rect 193355 8313 193367 8347
rect 193309 8307 193367 8313
rect 194042 8304 194048 8356
rect 194100 8304 194106 8356
rect 195256 8344 195284 8375
rect 195974 8372 195980 8384
rect 196032 8412 196038 8424
rect 196268 8412 196296 8452
rect 197357 8449 197369 8452
rect 197403 8449 197415 8483
rect 197357 8443 197415 8449
rect 197538 8440 197544 8492
rect 197596 8440 197602 8492
rect 197722 8440 197728 8492
rect 197780 8480 197786 8492
rect 198369 8483 198427 8489
rect 198369 8480 198381 8483
rect 197780 8452 198381 8480
rect 197780 8440 197786 8452
rect 198369 8449 198381 8452
rect 198415 8449 198427 8483
rect 198369 8443 198427 8449
rect 198550 8440 198556 8492
rect 198608 8440 198614 8492
rect 199013 8483 199071 8489
rect 199013 8449 199025 8483
rect 199059 8480 199071 8483
rect 199194 8480 199200 8492
rect 199059 8452 199200 8480
rect 199059 8449 199071 8452
rect 199013 8443 199071 8449
rect 199194 8440 199200 8452
rect 199252 8440 199258 8492
rect 199749 8483 199807 8489
rect 199749 8449 199761 8483
rect 199795 8480 199807 8483
rect 200206 8480 200212 8492
rect 199795 8452 200212 8480
rect 199795 8449 199807 8452
rect 199749 8443 199807 8449
rect 200206 8440 200212 8452
rect 200264 8440 200270 8492
rect 200577 8483 200635 8489
rect 200577 8449 200589 8483
rect 200623 8480 200635 8483
rect 201034 8480 201040 8492
rect 200623 8452 201040 8480
rect 200623 8449 200635 8452
rect 200577 8443 200635 8449
rect 201034 8440 201040 8452
rect 201092 8440 201098 8492
rect 201313 8483 201371 8489
rect 201313 8449 201325 8483
rect 201359 8480 201371 8483
rect 201862 8480 201868 8492
rect 201359 8452 201868 8480
rect 201359 8449 201371 8452
rect 201313 8443 201371 8449
rect 201862 8440 201868 8452
rect 201920 8440 201926 8492
rect 202506 8440 202512 8492
rect 202564 8440 202570 8492
rect 202690 8440 202696 8492
rect 202748 8440 202754 8492
rect 203337 8483 203395 8489
rect 203337 8480 203349 8483
rect 202800 8452 203349 8480
rect 196032 8384 196296 8412
rect 196032 8372 196038 8384
rect 197078 8372 197084 8424
rect 197136 8412 197142 8424
rect 197173 8415 197231 8421
rect 197173 8412 197185 8415
rect 197136 8384 197185 8412
rect 197136 8372 197142 8384
rect 197173 8381 197185 8384
rect 197219 8381 197231 8415
rect 197173 8375 197231 8381
rect 198185 8415 198243 8421
rect 198185 8381 198197 8415
rect 198231 8412 198243 8415
rect 198734 8412 198740 8424
rect 198231 8384 198740 8412
rect 198231 8381 198243 8384
rect 198185 8375 198243 8381
rect 198734 8372 198740 8384
rect 198792 8372 198798 8424
rect 202325 8415 202383 8421
rect 202325 8381 202337 8415
rect 202371 8381 202383 8415
rect 202524 8412 202552 8440
rect 202800 8412 202828 8452
rect 203337 8449 203349 8452
rect 203383 8449 203395 8483
rect 203337 8443 203395 8449
rect 203518 8440 203524 8492
rect 203576 8440 203582 8492
rect 202524 8384 202828 8412
rect 202325 8375 202383 8381
rect 195256 8316 195744 8344
rect 167104 8248 180794 8276
rect 195716 8276 195744 8316
rect 195790 8304 195796 8356
rect 195848 8344 195854 8356
rect 196253 8347 196311 8353
rect 196253 8344 196265 8347
rect 195848 8316 196265 8344
rect 195848 8304 195854 8316
rect 196253 8313 196265 8316
rect 196299 8313 196311 8347
rect 196253 8307 196311 8313
rect 199102 8304 199108 8356
rect 199160 8344 199166 8356
rect 199197 8347 199255 8353
rect 199197 8344 199209 8347
rect 199160 8316 199209 8344
rect 199160 8304 199166 8316
rect 199197 8313 199209 8316
rect 199243 8313 199255 8347
rect 199197 8307 199255 8313
rect 199930 8304 199936 8356
rect 199988 8304 199994 8356
rect 200758 8304 200764 8356
rect 200816 8304 200822 8356
rect 200942 8304 200948 8356
rect 201000 8344 201006 8356
rect 201497 8347 201555 8353
rect 201497 8344 201509 8347
rect 201000 8316 201509 8344
rect 201000 8304 201006 8316
rect 201497 8313 201509 8316
rect 201543 8313 201555 8347
rect 202340 8344 202368 8375
rect 202966 8372 202972 8424
rect 203024 8412 203030 8424
rect 203153 8415 203211 8421
rect 203153 8412 203165 8415
rect 203024 8384 203165 8412
rect 203024 8372 203030 8384
rect 203153 8381 203165 8384
rect 203199 8381 203211 8415
rect 203153 8375 203211 8381
rect 203242 8344 203248 8356
rect 202340 8316 203248 8344
rect 201497 8307 201555 8313
rect 203242 8304 203248 8316
rect 203300 8344 203306 8356
rect 211798 8344 211804 8356
rect 203300 8316 211804 8344
rect 203300 8304 203306 8316
rect 211798 8304 211804 8316
rect 211856 8304 211862 8356
rect 214024 8344 214052 8588
rect 216398 8576 216404 8628
rect 216456 8616 216462 8628
rect 219434 8616 219440 8628
rect 216456 8588 219440 8616
rect 216456 8576 216462 8588
rect 219434 8576 219440 8588
rect 219492 8576 219498 8628
rect 220906 8576 220912 8628
rect 220964 8616 220970 8628
rect 223482 8616 223488 8628
rect 220964 8588 223488 8616
rect 220964 8576 220970 8588
rect 223482 8576 223488 8588
rect 223540 8576 223546 8628
rect 224678 8576 224684 8628
rect 224736 8576 224742 8628
rect 224954 8576 224960 8628
rect 225012 8616 225018 8628
rect 225012 8588 225460 8616
rect 225012 8576 225018 8588
rect 215478 8508 215484 8560
rect 215536 8548 215542 8560
rect 217962 8548 217968 8560
rect 215536 8520 217968 8548
rect 215536 8508 215542 8520
rect 217962 8508 217968 8520
rect 218020 8508 218026 8560
rect 219250 8508 219256 8560
rect 219308 8548 219314 8560
rect 223206 8548 223212 8560
rect 219308 8520 223212 8548
rect 219308 8508 219314 8520
rect 223206 8508 223212 8520
rect 223264 8508 223270 8560
rect 223853 8551 223911 8557
rect 223853 8517 223865 8551
rect 223899 8548 223911 8551
rect 224402 8548 224408 8560
rect 223899 8520 224408 8548
rect 223899 8517 223911 8520
rect 223853 8511 223911 8517
rect 224402 8508 224408 8520
rect 224460 8508 224466 8560
rect 225432 8548 225460 8588
rect 225506 8576 225512 8628
rect 225564 8576 225570 8628
rect 225984 8588 226196 8616
rect 225984 8548 226012 8588
rect 225432 8520 226012 8548
rect 226168 8548 226196 8588
rect 226242 8576 226248 8628
rect 226300 8576 226306 8628
rect 226978 8576 226984 8628
rect 227036 8576 227042 8628
rect 227824 8588 228404 8616
rect 227824 8548 227852 8588
rect 226168 8520 227852 8548
rect 228376 8548 228404 8588
rect 228450 8576 228456 8628
rect 228508 8576 228514 8628
rect 229186 8576 229192 8628
rect 229244 8576 229250 8628
rect 230842 8616 230848 8628
rect 230032 8588 230848 8616
rect 230032 8548 230060 8588
rect 230842 8576 230848 8588
rect 230900 8576 230906 8628
rect 230934 8576 230940 8628
rect 230992 8576 230998 8628
rect 231670 8576 231676 8628
rect 231728 8576 231734 8628
rect 231762 8576 231768 8628
rect 231820 8616 231826 8628
rect 232498 8616 232504 8628
rect 231820 8588 232504 8616
rect 231820 8576 231826 8588
rect 232498 8576 232504 8588
rect 232556 8576 232562 8628
rect 232590 8576 232596 8628
rect 232648 8576 232654 8628
rect 234430 8576 234436 8628
rect 234488 8576 234494 8628
rect 236270 8576 236276 8628
rect 236328 8576 236334 8628
rect 248874 8616 248880 8628
rect 236564 8588 248880 8616
rect 228376 8520 230060 8548
rect 215202 8440 215208 8492
rect 215260 8480 215266 8492
rect 220446 8480 220452 8492
rect 215260 8452 220452 8480
rect 215260 8440 215266 8452
rect 220446 8440 220452 8452
rect 220504 8440 220510 8492
rect 221458 8440 221464 8492
rect 221516 8480 221522 8492
rect 223669 8483 223727 8489
rect 223669 8480 223681 8483
rect 221516 8452 223681 8480
rect 221516 8440 221522 8452
rect 223669 8449 223681 8452
rect 223715 8480 223727 8483
rect 223715 8452 223896 8480
rect 223715 8449 223727 8452
rect 223669 8443 223727 8449
rect 219084 8384 220952 8412
rect 214024 8316 215294 8344
rect 195974 8276 195980 8288
rect 195716 8248 195980 8276
rect 195974 8236 195980 8248
rect 196032 8276 196038 8288
rect 196158 8276 196164 8288
rect 196032 8248 196164 8276
rect 196032 8236 196038 8248
rect 196158 8236 196164 8248
rect 196216 8236 196222 8288
rect 215266 8276 215294 8316
rect 219084 8276 219112 8384
rect 219158 8304 219164 8356
rect 219216 8344 219222 8356
rect 220924 8344 220952 8384
rect 221274 8372 221280 8424
rect 221332 8412 221338 8424
rect 223758 8412 223764 8424
rect 221332 8384 223764 8412
rect 221332 8372 221338 8384
rect 223758 8372 223764 8384
rect 223816 8372 223822 8424
rect 223868 8412 223896 8452
rect 224034 8440 224040 8492
rect 224092 8480 224098 8492
rect 224092 8452 224356 8480
rect 224092 8440 224098 8452
rect 224218 8412 224224 8424
rect 223868 8384 224224 8412
rect 224218 8372 224224 8384
rect 224276 8372 224282 8424
rect 224328 8412 224356 8452
rect 224494 8440 224500 8492
rect 224552 8440 224558 8492
rect 225322 8440 225328 8492
rect 225380 8440 225386 8492
rect 226058 8440 226064 8492
rect 226116 8440 226122 8492
rect 226794 8440 226800 8492
rect 226852 8440 226858 8492
rect 227806 8440 227812 8492
rect 227864 8480 227870 8492
rect 228085 8483 228143 8489
rect 228085 8480 228097 8483
rect 227864 8452 228097 8480
rect 227864 8440 227870 8452
rect 228085 8449 228097 8452
rect 228131 8449 228143 8483
rect 228085 8443 228143 8449
rect 226242 8412 226248 8424
rect 224328 8384 226248 8412
rect 226242 8372 226248 8384
rect 226300 8372 226306 8424
rect 228100 8412 228128 8443
rect 228266 8440 228272 8492
rect 228324 8440 228330 8492
rect 229002 8440 229008 8492
rect 229060 8440 229066 8492
rect 230032 8489 230060 8520
rect 230198 8508 230204 8560
rect 230256 8548 230262 8560
rect 232314 8548 232320 8560
rect 230256 8520 232320 8548
rect 230256 8508 230262 8520
rect 232314 8508 232320 8520
rect 232372 8508 232378 8560
rect 236564 8548 236592 8588
rect 248874 8576 248880 8588
rect 248932 8576 248938 8628
rect 248966 8576 248972 8628
rect 249024 8616 249030 8628
rect 251542 8616 251548 8628
rect 249024 8588 251548 8616
rect 249024 8576 249030 8588
rect 251542 8576 251548 8588
rect 251600 8576 251606 8628
rect 258258 8576 258264 8628
rect 258316 8576 258322 8628
rect 259178 8576 259184 8628
rect 259236 8576 259242 8628
rect 259914 8576 259920 8628
rect 259972 8576 259978 8628
rect 260466 8576 260472 8628
rect 260524 8576 260530 8628
rect 261846 8576 261852 8628
rect 261904 8616 261910 8628
rect 262309 8619 262367 8625
rect 262309 8616 262321 8619
rect 261904 8588 262321 8616
rect 261904 8576 261910 8588
rect 262309 8585 262321 8588
rect 262355 8585 262367 8619
rect 262309 8579 262367 8585
rect 262582 8576 262588 8628
rect 262640 8616 262646 8628
rect 262640 8588 265388 8616
rect 262640 8576 262646 8588
rect 232700 8520 236592 8548
rect 230017 8483 230075 8489
rect 230017 8449 230029 8483
rect 230063 8449 230075 8483
rect 230017 8443 230075 8449
rect 230106 8440 230112 8492
rect 230164 8440 230170 8492
rect 230293 8483 230351 8489
rect 230293 8449 230305 8483
rect 230339 8480 230351 8483
rect 230753 8483 230811 8489
rect 230753 8480 230765 8483
rect 230339 8452 230765 8480
rect 230339 8449 230351 8452
rect 230293 8443 230351 8449
rect 230753 8449 230765 8452
rect 230799 8449 230811 8483
rect 230753 8443 230811 8449
rect 231486 8440 231492 8492
rect 231544 8440 231550 8492
rect 232406 8440 232412 8492
rect 232464 8440 232470 8492
rect 232700 8486 232728 8520
rect 239306 8508 239312 8560
rect 239364 8548 239370 8560
rect 263870 8548 263876 8560
rect 239364 8520 257108 8548
rect 239364 8508 239370 8520
rect 232516 8458 232728 8486
rect 233605 8483 233663 8489
rect 228910 8412 228916 8424
rect 228100 8384 228916 8412
rect 228910 8372 228916 8384
rect 228968 8372 228974 8424
rect 229094 8372 229100 8424
rect 229152 8412 229158 8424
rect 229646 8412 229652 8424
rect 229152 8384 229652 8412
rect 229152 8372 229158 8384
rect 229646 8372 229652 8384
rect 229704 8372 229710 8424
rect 232516 8412 232544 8458
rect 233605 8449 233617 8483
rect 233651 8480 233663 8483
rect 233694 8480 233700 8492
rect 233651 8452 233700 8480
rect 233651 8449 233663 8452
rect 233605 8443 233663 8449
rect 233694 8440 233700 8452
rect 233752 8440 233758 8492
rect 233789 8483 233847 8489
rect 233789 8449 233801 8483
rect 233835 8480 233847 8483
rect 234249 8483 234307 8489
rect 234249 8480 234261 8483
rect 233835 8452 234261 8480
rect 233835 8449 233847 8452
rect 233789 8443 233847 8449
rect 234249 8449 234261 8452
rect 234295 8449 234307 8483
rect 234249 8443 234307 8449
rect 234430 8440 234436 8492
rect 234488 8480 234494 8492
rect 235261 8483 235319 8489
rect 235261 8480 235273 8483
rect 234488 8452 235273 8480
rect 234488 8440 234494 8452
rect 235261 8449 235273 8452
rect 235307 8449 235319 8483
rect 235261 8443 235319 8449
rect 235445 8483 235503 8489
rect 235445 8449 235457 8483
rect 235491 8480 235503 8483
rect 236089 8483 236147 8489
rect 236089 8480 236101 8483
rect 235491 8452 236101 8480
rect 235491 8449 235503 8452
rect 235445 8443 235503 8449
rect 236089 8449 236101 8452
rect 236135 8449 236147 8483
rect 250254 8480 250260 8492
rect 236089 8443 236147 8449
rect 244246 8452 250260 8480
rect 230032 8384 232544 8412
rect 224770 8344 224776 8356
rect 219216 8316 220860 8344
rect 220924 8316 224776 8344
rect 219216 8304 219222 8316
rect 215266 8248 219112 8276
rect 220832 8276 220860 8316
rect 224770 8304 224776 8316
rect 224828 8304 224834 8356
rect 224862 8304 224868 8356
rect 224920 8344 224926 8356
rect 228358 8344 228364 8356
rect 224920 8316 228364 8344
rect 224920 8304 224926 8316
rect 228358 8304 228364 8316
rect 228416 8304 228422 8356
rect 228450 8304 228456 8356
rect 228508 8344 228514 8356
rect 230032 8344 230060 8384
rect 233418 8372 233424 8424
rect 233476 8372 233482 8424
rect 235077 8415 235135 8421
rect 235077 8381 235089 8415
rect 235123 8412 235135 8415
rect 235810 8412 235816 8424
rect 235123 8384 235816 8412
rect 235123 8381 235135 8384
rect 235077 8375 235135 8381
rect 235810 8372 235816 8384
rect 235868 8372 235874 8424
rect 235994 8372 236000 8424
rect 236052 8412 236058 8424
rect 244246 8412 244274 8452
rect 250254 8440 250260 8452
rect 250312 8440 250318 8492
rect 256694 8440 256700 8492
rect 256752 8440 256758 8492
rect 236052 8384 244274 8412
rect 236052 8372 236058 8384
rect 256970 8372 256976 8424
rect 257028 8372 257034 8424
rect 257080 8412 257108 8520
rect 259104 8520 263876 8548
rect 258074 8440 258080 8492
rect 258132 8440 258138 8492
rect 258258 8440 258264 8492
rect 258316 8480 258322 8492
rect 259104 8489 259132 8520
rect 263870 8508 263876 8520
rect 263928 8508 263934 8560
rect 264238 8508 264244 8560
rect 264296 8548 264302 8560
rect 264514 8548 264520 8560
rect 264296 8520 264520 8548
rect 264296 8508 264302 8520
rect 264514 8508 264520 8520
rect 264572 8548 264578 8560
rect 264885 8551 264943 8557
rect 264885 8548 264897 8551
rect 264572 8520 264897 8548
rect 264572 8508 264578 8520
rect 264885 8517 264897 8520
rect 264931 8517 264943 8551
rect 264885 8511 264943 8517
rect 259089 8483 259147 8489
rect 259089 8480 259101 8483
rect 258316 8452 259101 8480
rect 258316 8440 258322 8452
rect 259089 8449 259101 8452
rect 259135 8449 259147 8483
rect 259089 8443 259147 8449
rect 259730 8440 259736 8492
rect 259788 8440 259794 8492
rect 260282 8440 260288 8492
rect 260340 8440 260346 8492
rect 260374 8440 260380 8492
rect 260432 8480 260438 8492
rect 261297 8483 261355 8489
rect 261297 8480 261309 8483
rect 260432 8452 260834 8480
rect 260432 8440 260438 8452
rect 257080 8384 260512 8412
rect 228508 8316 230060 8344
rect 228508 8304 228514 8316
rect 230566 8304 230572 8356
rect 230624 8344 230630 8356
rect 233436 8344 233464 8372
rect 230624 8316 233464 8344
rect 230624 8304 230630 8316
rect 236454 8304 236460 8356
rect 236512 8344 236518 8356
rect 260374 8344 260380 8356
rect 236512 8316 260380 8344
rect 236512 8304 236518 8316
rect 260374 8304 260380 8316
rect 260432 8304 260438 8356
rect 224586 8276 224592 8288
rect 220832 8248 224592 8276
rect 224586 8236 224592 8248
rect 224644 8236 224650 8288
rect 224678 8236 224684 8288
rect 224736 8276 224742 8288
rect 232498 8276 232504 8288
rect 224736 8248 232504 8276
rect 224736 8236 224742 8248
rect 232498 8236 232504 8248
rect 232556 8236 232562 8288
rect 232682 8236 232688 8288
rect 232740 8276 232746 8288
rect 249058 8276 249064 8288
rect 232740 8248 249064 8276
rect 232740 8236 232746 8248
rect 249058 8236 249064 8248
rect 249116 8236 249122 8288
rect 251266 8236 251272 8288
rect 251324 8276 251330 8288
rect 258718 8276 258724 8288
rect 251324 8248 258724 8276
rect 251324 8236 251330 8248
rect 258718 8236 258724 8248
rect 258776 8236 258782 8288
rect 260484 8276 260512 8384
rect 260806 8344 260834 8452
rect 260944 8452 261309 8480
rect 260944 8424 260972 8452
rect 261297 8449 261309 8452
rect 261343 8449 261355 8483
rect 261297 8443 261355 8449
rect 261478 8440 261484 8492
rect 261536 8480 261542 8492
rect 262125 8483 262183 8489
rect 262125 8480 262137 8483
rect 261536 8452 262137 8480
rect 261536 8440 261542 8452
rect 262125 8449 262137 8452
rect 262171 8449 262183 8483
rect 262125 8443 262183 8449
rect 262953 8483 263011 8489
rect 262953 8449 262965 8483
rect 262999 8480 263011 8483
rect 263042 8480 263048 8492
rect 262999 8452 263048 8480
rect 262999 8449 263011 8452
rect 262953 8443 263011 8449
rect 263042 8440 263048 8452
rect 263100 8440 263106 8492
rect 265360 8489 265388 8588
rect 265618 8576 265624 8628
rect 265676 8616 265682 8628
rect 265805 8619 265863 8625
rect 265805 8616 265817 8619
rect 265676 8588 265817 8616
rect 265676 8576 265682 8588
rect 265805 8585 265817 8588
rect 265851 8585 265863 8619
rect 265805 8579 265863 8585
rect 266262 8576 266268 8628
rect 266320 8616 266326 8628
rect 266320 8588 267044 8616
rect 266320 8576 266326 8588
rect 265894 8508 265900 8560
rect 265952 8548 265958 8560
rect 266909 8551 266967 8557
rect 266909 8548 266921 8551
rect 265952 8520 266921 8548
rect 265952 8508 265958 8520
rect 266909 8517 266921 8520
rect 266955 8517 266967 8551
rect 267016 8548 267044 8588
rect 267090 8576 267096 8628
rect 267148 8616 267154 8628
rect 270497 8619 270555 8625
rect 270497 8616 270509 8619
rect 267148 8588 270509 8616
rect 267148 8576 267154 8588
rect 270497 8585 270509 8588
rect 270543 8585 270555 8619
rect 270497 8579 270555 8585
rect 268010 8548 268016 8560
rect 267016 8520 268016 8548
rect 266909 8511 266967 8517
rect 268010 8508 268016 8520
rect 268068 8508 268074 8560
rect 268120 8520 269620 8548
rect 265345 8483 265403 8489
rect 263796 8452 264008 8480
rect 260926 8372 260932 8424
rect 260984 8372 260990 8424
rect 261386 8372 261392 8424
rect 261444 8412 261450 8424
rect 261573 8415 261631 8421
rect 261573 8412 261585 8415
rect 261444 8384 261585 8412
rect 261444 8372 261450 8384
rect 261573 8381 261585 8384
rect 261619 8381 261631 8415
rect 261573 8375 261631 8381
rect 262398 8372 262404 8424
rect 262456 8412 262462 8424
rect 263796 8412 263824 8452
rect 262456 8384 263824 8412
rect 263980 8412 264008 8452
rect 265345 8449 265357 8483
rect 265391 8480 265403 8483
rect 265710 8480 265716 8492
rect 265391 8452 265716 8480
rect 265391 8449 265403 8452
rect 265345 8443 265403 8449
rect 265710 8440 265716 8452
rect 265768 8440 265774 8492
rect 265802 8440 265808 8492
rect 265860 8480 265866 8492
rect 265860 8452 266676 8480
rect 265860 8440 265866 8452
rect 263980 8384 266492 8412
rect 262456 8372 262462 8384
rect 263870 8344 263876 8356
rect 260806 8316 263876 8344
rect 263870 8304 263876 8316
rect 263928 8304 263934 8356
rect 263962 8304 263968 8356
rect 264020 8344 264026 8356
rect 264238 8344 264244 8356
rect 264020 8316 264244 8344
rect 264020 8304 264026 8316
rect 264238 8304 264244 8316
rect 264296 8344 264302 8356
rect 264425 8347 264483 8353
rect 264425 8344 264437 8347
rect 264296 8316 264437 8344
rect 264296 8304 264302 8316
rect 264425 8313 264437 8316
rect 264471 8313 264483 8347
rect 266464 8344 266492 8384
rect 266538 8372 266544 8424
rect 266596 8372 266602 8424
rect 266648 8412 266676 8452
rect 266722 8440 266728 8492
rect 266780 8440 266786 8492
rect 266832 8452 267596 8480
rect 266832 8412 266860 8452
rect 266648 8384 266860 8412
rect 267274 8372 267280 8424
rect 267332 8412 267338 8424
rect 267461 8415 267519 8421
rect 267461 8412 267473 8415
rect 267332 8384 267473 8412
rect 267332 8372 267338 8384
rect 267461 8381 267473 8384
rect 267507 8381 267519 8415
rect 267568 8412 267596 8452
rect 267642 8440 267648 8492
rect 267700 8440 267706 8492
rect 268120 8480 268148 8520
rect 267752 8452 268148 8480
rect 267752 8412 267780 8452
rect 268378 8440 268384 8492
rect 268436 8480 268442 8492
rect 268746 8480 268752 8492
rect 268436 8452 268752 8480
rect 268436 8440 268442 8452
rect 268746 8440 268752 8452
rect 268804 8440 268810 8492
rect 269592 8489 269620 8520
rect 269577 8483 269635 8489
rect 269577 8449 269589 8483
rect 269623 8449 269635 8483
rect 269577 8443 269635 8449
rect 269758 8440 269764 8492
rect 269816 8480 269822 8492
rect 270405 8483 270463 8489
rect 270405 8480 270417 8483
rect 269816 8452 270417 8480
rect 269816 8440 269822 8452
rect 270405 8449 270417 8452
rect 270451 8449 270463 8483
rect 270405 8443 270463 8449
rect 270678 8440 270684 8492
rect 270736 8440 270742 8492
rect 267568 8384 267780 8412
rect 267829 8415 267887 8421
rect 267461 8375 267519 8381
rect 267829 8381 267841 8415
rect 267875 8412 267887 8415
rect 269298 8412 269304 8424
rect 267875 8384 269304 8412
rect 267875 8381 267887 8384
rect 267829 8375 267887 8381
rect 269298 8372 269304 8384
rect 269356 8372 269362 8424
rect 269485 8415 269543 8421
rect 269485 8381 269497 8415
rect 269531 8381 269543 8415
rect 269485 8375 269543 8381
rect 269500 8344 269528 8375
rect 270494 8344 270500 8356
rect 264425 8307 264483 8313
rect 265728 8316 265940 8344
rect 266464 8316 269528 8344
rect 269592 8316 270500 8344
rect 262950 8276 262956 8288
rect 260484 8248 262956 8276
rect 262950 8236 262956 8248
rect 263008 8276 263014 8288
rect 263045 8279 263103 8285
rect 263045 8276 263057 8279
rect 263008 8248 263057 8276
rect 263008 8236 263014 8248
rect 263045 8245 263057 8248
rect 263091 8245 263103 8279
rect 263045 8239 263103 8245
rect 263226 8236 263232 8288
rect 263284 8276 263290 8288
rect 264054 8276 264060 8288
rect 263284 8248 264060 8276
rect 263284 8236 263290 8248
rect 264054 8236 264060 8248
rect 264112 8236 264118 8288
rect 265158 8236 265164 8288
rect 265216 8276 265222 8288
rect 265728 8276 265756 8316
rect 265216 8248 265756 8276
rect 265912 8276 265940 8316
rect 268378 8276 268384 8288
rect 265912 8248 268384 8276
rect 265216 8236 265222 8248
rect 268378 8236 268384 8248
rect 268436 8236 268442 8288
rect 268470 8236 268476 8288
rect 268528 8276 268534 8288
rect 269592 8276 269620 8316
rect 270494 8304 270500 8316
rect 270552 8304 270558 8356
rect 268528 8248 269620 8276
rect 269945 8279 270003 8285
rect 268528 8236 268534 8248
rect 269945 8245 269957 8279
rect 269991 8276 270003 8279
rect 270034 8276 270040 8288
rect 269991 8248 270040 8276
rect 269991 8245 270003 8248
rect 269945 8239 270003 8245
rect 270034 8236 270040 8248
rect 270092 8236 270098 8288
rect 1104 8186 271492 8208
rect 1104 8134 34748 8186
rect 34800 8134 34812 8186
rect 34864 8134 34876 8186
rect 34928 8134 34940 8186
rect 34992 8134 35004 8186
rect 35056 8134 102345 8186
rect 102397 8134 102409 8186
rect 102461 8134 102473 8186
rect 102525 8134 102537 8186
rect 102589 8134 102601 8186
rect 102653 8134 169942 8186
rect 169994 8134 170006 8186
rect 170058 8134 170070 8186
rect 170122 8134 170134 8186
rect 170186 8134 170198 8186
rect 170250 8134 237539 8186
rect 237591 8134 237603 8186
rect 237655 8134 237667 8186
rect 237719 8134 237731 8186
rect 237783 8134 237795 8186
rect 237847 8134 271492 8186
rect 1104 8112 271492 8134
rect 9674 8032 9680 8084
rect 9732 8072 9738 8084
rect 39206 8072 39212 8084
rect 9732 8044 39212 8072
rect 9732 8032 9738 8044
rect 39206 8032 39212 8044
rect 39264 8032 39270 8084
rect 66990 8032 66996 8084
rect 67048 8072 67054 8084
rect 67269 8075 67327 8081
rect 67269 8072 67281 8075
rect 67048 8044 67281 8072
rect 67048 8032 67054 8044
rect 67269 8041 67281 8044
rect 67315 8041 67327 8075
rect 67269 8035 67327 8041
rect 77570 8032 77576 8084
rect 77628 8072 77634 8084
rect 84102 8072 84108 8084
rect 77628 8044 84108 8072
rect 77628 8032 77634 8044
rect 84102 8032 84108 8044
rect 84160 8032 84166 8084
rect 86678 8032 86684 8084
rect 86736 8072 86742 8084
rect 100478 8072 100484 8084
rect 86736 8044 100484 8072
rect 86736 8032 86742 8044
rect 100478 8032 100484 8044
rect 100536 8032 100542 8084
rect 100849 8075 100907 8081
rect 100849 8041 100861 8075
rect 100895 8072 100907 8075
rect 101030 8072 101036 8084
rect 100895 8044 101036 8072
rect 100895 8041 100907 8044
rect 100849 8035 100907 8041
rect 101030 8032 101036 8044
rect 101088 8032 101094 8084
rect 109586 8072 109592 8084
rect 101140 8044 109592 8072
rect 21910 7964 21916 8016
rect 21968 7964 21974 8016
rect 22922 7964 22928 8016
rect 22980 7964 22986 8016
rect 23658 7964 23664 8016
rect 23716 7964 23722 8016
rect 25222 7964 25228 8016
rect 25280 7964 25286 8016
rect 25314 7964 25320 8016
rect 25372 8004 25378 8016
rect 48958 8004 48964 8016
rect 25372 7976 48964 8004
rect 25372 7964 25378 7976
rect 48958 7964 48964 7976
rect 49016 7964 49022 8016
rect 74994 7964 75000 8016
rect 75052 8004 75058 8016
rect 95142 8004 95148 8016
rect 75052 7976 95148 8004
rect 75052 7964 75058 7976
rect 95142 7964 95148 7976
rect 95200 7964 95206 8016
rect 100662 7964 100668 8016
rect 100720 8004 100726 8016
rect 101140 8004 101168 8044
rect 109586 8032 109592 8044
rect 109644 8032 109650 8084
rect 116854 8072 116860 8084
rect 109788 8044 116860 8072
rect 100720 7976 101168 8004
rect 100720 7964 100726 7976
rect 101490 7964 101496 8016
rect 101548 8004 101554 8016
rect 109788 8004 109816 8044
rect 116854 8032 116860 8044
rect 116912 8032 116918 8084
rect 129274 8032 129280 8084
rect 129332 8032 129338 8084
rect 132954 8032 132960 8084
rect 133012 8032 133018 8084
rect 148594 8032 148600 8084
rect 148652 8072 148658 8084
rect 153562 8072 153568 8084
rect 148652 8044 153568 8072
rect 148652 8032 148658 8044
rect 153562 8032 153568 8044
rect 153620 8032 153626 8084
rect 157242 8032 157248 8084
rect 157300 8032 157306 8084
rect 158714 8032 158720 8084
rect 158772 8032 158778 8084
rect 159450 8032 159456 8084
rect 159508 8072 159514 8084
rect 160189 8075 160247 8081
rect 160189 8072 160201 8075
rect 159508 8044 160201 8072
rect 159508 8032 159514 8044
rect 160189 8041 160201 8044
rect 160235 8041 160247 8075
rect 160189 8035 160247 8041
rect 160922 8032 160928 8084
rect 160980 8032 160986 8084
rect 161014 8032 161020 8084
rect 161072 8072 161078 8084
rect 161661 8075 161719 8081
rect 161661 8072 161673 8075
rect 161072 8044 161673 8072
rect 161072 8032 161078 8044
rect 161661 8041 161673 8044
rect 161707 8041 161719 8075
rect 161661 8035 161719 8041
rect 162394 8032 162400 8084
rect 162452 8032 162458 8084
rect 163866 8032 163872 8084
rect 163924 8032 163930 8084
rect 163958 8032 163964 8084
rect 164016 8072 164022 8084
rect 164605 8075 164663 8081
rect 164605 8072 164617 8075
rect 164016 8044 164617 8072
rect 164016 8032 164022 8044
rect 164605 8041 164617 8044
rect 164651 8041 164663 8075
rect 164605 8035 164663 8041
rect 165338 8032 165344 8084
rect 165396 8072 165402 8084
rect 166077 8075 166135 8081
rect 166077 8072 166089 8075
rect 165396 8044 166089 8072
rect 165396 8032 165402 8044
rect 166077 8041 166089 8044
rect 166123 8041 166135 8075
rect 177666 8072 177672 8084
rect 166077 8035 166135 8041
rect 166184 8044 177672 8072
rect 101548 7976 109816 8004
rect 109865 8007 109923 8013
rect 101548 7964 101554 7976
rect 109865 7973 109877 8007
rect 109911 7973 109923 8007
rect 117866 8004 117872 8016
rect 109865 7967 109923 7973
rect 109972 7976 117872 8004
rect 16482 7896 16488 7948
rect 16540 7936 16546 7948
rect 16540 7908 25176 7936
rect 16540 7896 16546 7908
rect 21634 7828 21640 7880
rect 21692 7868 21698 7880
rect 21729 7871 21787 7877
rect 21729 7868 21741 7871
rect 21692 7840 21741 7868
rect 21692 7828 21698 7840
rect 21729 7837 21741 7840
rect 21775 7837 21787 7871
rect 21729 7831 21787 7837
rect 22738 7828 22744 7880
rect 22796 7828 22802 7880
rect 23474 7828 23480 7880
rect 23532 7828 23538 7880
rect 25038 7828 25044 7880
rect 25096 7828 25102 7880
rect 25148 7868 25176 7908
rect 32858 7896 32864 7948
rect 32916 7896 32922 7948
rect 46106 7936 46112 7948
rect 33888 7908 46112 7936
rect 33888 7868 33916 7908
rect 46106 7896 46112 7908
rect 46164 7896 46170 7948
rect 66901 7939 66959 7945
rect 66901 7905 66913 7939
rect 66947 7936 66959 7939
rect 67729 7939 67787 7945
rect 67729 7936 67741 7939
rect 66947 7908 67741 7936
rect 66947 7905 66959 7908
rect 66901 7899 66959 7905
rect 67729 7905 67741 7908
rect 67775 7905 67787 7939
rect 67729 7899 67787 7905
rect 73706 7896 73712 7948
rect 73764 7936 73770 7948
rect 88518 7936 88524 7948
rect 73764 7908 88524 7936
rect 73764 7896 73770 7908
rect 88518 7896 88524 7908
rect 88576 7896 88582 7948
rect 92566 7896 92572 7948
rect 92624 7936 92630 7948
rect 96614 7936 96620 7948
rect 92624 7908 96620 7936
rect 92624 7896 92630 7908
rect 96614 7896 96620 7908
rect 96672 7896 96678 7948
rect 100481 7939 100539 7945
rect 100481 7905 100493 7939
rect 100527 7936 100539 7939
rect 101950 7936 101956 7948
rect 100527 7908 101956 7936
rect 100527 7905 100539 7908
rect 100481 7899 100539 7905
rect 101950 7896 101956 7908
rect 102008 7896 102014 7948
rect 104434 7896 104440 7948
rect 104492 7936 104498 7948
rect 109880 7936 109908 7967
rect 104492 7908 109908 7936
rect 104492 7896 104498 7908
rect 25148 7840 33916 7868
rect 33962 7828 33968 7880
rect 34020 7868 34026 7880
rect 51718 7868 51724 7880
rect 34020 7840 51724 7868
rect 34020 7828 34026 7840
rect 51718 7828 51724 7840
rect 51776 7828 51782 7880
rect 67082 7828 67088 7880
rect 67140 7828 67146 7880
rect 89533 7871 89591 7877
rect 89533 7837 89545 7871
rect 89579 7868 89591 7871
rect 90082 7868 90088 7880
rect 89579 7840 90088 7868
rect 89579 7837 89591 7840
rect 89533 7831 89591 7837
rect 90082 7828 90088 7840
rect 90140 7828 90146 7880
rect 91480 7840 91692 7868
rect 18414 7760 18420 7812
rect 18472 7800 18478 7812
rect 25314 7800 25320 7812
rect 18472 7772 25320 7800
rect 18472 7760 18478 7772
rect 25314 7760 25320 7772
rect 25372 7760 25378 7812
rect 51626 7800 51632 7812
rect 26896 7772 34100 7800
rect 19150 7692 19156 7744
rect 19208 7732 19214 7744
rect 26896 7732 26924 7772
rect 19208 7704 26924 7732
rect 19208 7692 19214 7704
rect 27614 7692 27620 7744
rect 27672 7732 27678 7744
rect 33962 7732 33968 7744
rect 27672 7704 33968 7732
rect 27672 7692 27678 7704
rect 33962 7692 33968 7704
rect 34020 7692 34026 7744
rect 34072 7732 34100 7772
rect 41386 7772 51632 7800
rect 41386 7732 41414 7772
rect 51626 7760 51632 7772
rect 51684 7760 51690 7812
rect 83274 7760 83280 7812
rect 83332 7800 83338 7812
rect 91480 7800 91508 7840
rect 83332 7772 91508 7800
rect 91664 7800 91692 7840
rect 91922 7828 91928 7880
rect 91980 7868 91986 7880
rect 99282 7868 99288 7880
rect 91980 7840 99288 7868
rect 91980 7828 91986 7840
rect 99282 7828 99288 7840
rect 99340 7828 99346 7880
rect 100665 7871 100723 7877
rect 100665 7837 100677 7871
rect 100711 7868 100723 7871
rect 100938 7868 100944 7880
rect 100711 7840 100944 7868
rect 100711 7837 100723 7840
rect 100665 7831 100723 7837
rect 100938 7828 100944 7840
rect 100996 7828 101002 7880
rect 107746 7868 107752 7880
rect 103624 7840 107752 7868
rect 103624 7800 103652 7840
rect 107746 7828 107752 7840
rect 107804 7828 107810 7880
rect 109310 7828 109316 7880
rect 109368 7828 109374 7880
rect 109586 7828 109592 7880
rect 109644 7868 109650 7880
rect 109972 7868 110000 7976
rect 117866 7964 117872 7976
rect 117924 7964 117930 8016
rect 156598 7964 156604 8016
rect 156656 8004 156662 8016
rect 164694 8004 164700 8016
rect 156656 7976 164700 8004
rect 156656 7964 156662 7976
rect 164694 7964 164700 7976
rect 164752 7964 164758 8016
rect 112806 7896 112812 7948
rect 112864 7936 112870 7948
rect 120902 7936 120908 7948
rect 112864 7908 120908 7936
rect 112864 7896 112870 7908
rect 120902 7896 120908 7908
rect 120960 7896 120966 7948
rect 134242 7896 134248 7948
rect 134300 7896 134306 7948
rect 143994 7896 144000 7948
rect 144052 7936 144058 7948
rect 161934 7936 161940 7948
rect 144052 7908 161940 7936
rect 144052 7896 144058 7908
rect 161934 7896 161940 7908
rect 161992 7896 161998 7948
rect 166184 7936 166212 8044
rect 177666 8032 177672 8044
rect 177724 8032 177730 8084
rect 197170 8032 197176 8084
rect 197228 8072 197234 8084
rect 219066 8072 219072 8084
rect 197228 8044 219072 8072
rect 197228 8032 197234 8044
rect 219066 8032 219072 8044
rect 219124 8032 219130 8084
rect 221090 8032 221096 8084
rect 221148 8072 221154 8084
rect 249794 8072 249800 8084
rect 221148 8044 249800 8072
rect 221148 8032 221154 8044
rect 249794 8032 249800 8044
rect 249852 8032 249858 8084
rect 259546 8032 259552 8084
rect 259604 8032 259610 8084
rect 259730 8032 259736 8084
rect 259788 8072 259794 8084
rect 260837 8075 260895 8081
rect 260837 8072 260849 8075
rect 259788 8044 260849 8072
rect 259788 8032 259794 8044
rect 260837 8041 260849 8044
rect 260883 8041 260895 8075
rect 260837 8035 260895 8041
rect 261754 8032 261760 8084
rect 261812 8032 261818 8084
rect 262490 8032 262496 8084
rect 262548 8032 262554 8084
rect 263318 8032 263324 8084
rect 263376 8032 263382 8084
rect 264072 8044 264836 8072
rect 166626 8004 166632 8016
rect 162044 7908 166212 7936
rect 166552 7976 166632 8004
rect 109644 7840 110000 7868
rect 109644 7828 109650 7840
rect 110046 7828 110052 7880
rect 110104 7828 110110 7880
rect 114925 7871 114983 7877
rect 114925 7837 114937 7871
rect 114971 7868 114983 7871
rect 115382 7868 115388 7880
rect 114971 7840 115388 7868
rect 114971 7837 114983 7840
rect 114925 7831 114983 7837
rect 115382 7828 115388 7840
rect 115440 7828 115446 7880
rect 116121 7871 116179 7877
rect 116121 7837 116133 7871
rect 116167 7868 116179 7871
rect 117498 7868 117504 7880
rect 116167 7840 117504 7868
rect 116167 7837 116179 7840
rect 116121 7831 116179 7837
rect 117498 7828 117504 7840
rect 117556 7828 117562 7880
rect 129090 7828 129096 7880
rect 129148 7828 129154 7880
rect 132770 7828 132776 7880
rect 132828 7828 132834 7880
rect 146478 7828 146484 7880
rect 146536 7868 146542 7880
rect 154574 7868 154580 7880
rect 146536 7840 154580 7868
rect 146536 7828 146542 7840
rect 154574 7828 154580 7840
rect 154632 7828 154638 7880
rect 157058 7828 157064 7880
rect 157116 7828 157122 7880
rect 158530 7828 158536 7880
rect 158588 7828 158594 7880
rect 159266 7828 159272 7880
rect 159324 7828 159330 7880
rect 160002 7828 160008 7880
rect 160060 7828 160066 7880
rect 160738 7828 160744 7880
rect 160796 7828 160802 7880
rect 161474 7828 161480 7880
rect 161532 7828 161538 7880
rect 91664 7772 103652 7800
rect 83332 7760 83338 7772
rect 104158 7760 104164 7812
rect 104216 7800 104222 7812
rect 104216 7772 114968 7800
rect 104216 7760 104222 7772
rect 114940 7744 114968 7772
rect 115290 7760 115296 7812
rect 115348 7800 115354 7812
rect 115750 7800 115756 7812
rect 115348 7772 115756 7800
rect 115348 7760 115354 7772
rect 115750 7760 115756 7772
rect 115808 7800 115814 7812
rect 116213 7803 116271 7809
rect 116213 7800 116225 7803
rect 115808 7772 116225 7800
rect 115808 7760 115814 7772
rect 116213 7769 116225 7772
rect 116259 7769 116271 7803
rect 116213 7763 116271 7769
rect 151998 7760 152004 7812
rect 152056 7800 152062 7812
rect 162044 7800 162072 7908
rect 162210 7828 162216 7880
rect 162268 7828 162274 7880
rect 163682 7828 163688 7880
rect 163740 7828 163746 7880
rect 164418 7828 164424 7880
rect 164476 7828 164482 7880
rect 165154 7828 165160 7880
rect 165212 7828 165218 7880
rect 165890 7828 165896 7880
rect 165948 7828 165954 7880
rect 166552 7868 166580 7976
rect 166626 7964 166632 7976
rect 166684 7964 166690 8016
rect 168193 8007 168251 8013
rect 168193 7973 168205 8007
rect 168239 8004 168251 8007
rect 169018 8004 169024 8016
rect 168239 7976 169024 8004
rect 168239 7973 168251 7976
rect 168193 7967 168251 7973
rect 169018 7964 169024 7976
rect 169076 7964 169082 8016
rect 169202 7964 169208 8016
rect 169260 7964 169266 8016
rect 169662 7964 169668 8016
rect 169720 8004 169726 8016
rect 169720 7976 169892 8004
rect 169720 7964 169726 7976
rect 166810 7896 166816 7948
rect 166868 7936 166874 7948
rect 168837 7939 168895 7945
rect 166868 7908 168052 7936
rect 166868 7896 166874 7908
rect 166617 7871 166675 7877
rect 166617 7868 166629 7871
rect 166552 7840 166629 7868
rect 166617 7837 166629 7840
rect 166663 7837 166675 7871
rect 166617 7831 166675 7837
rect 167822 7828 167828 7880
rect 167880 7828 167886 7880
rect 168024 7877 168052 7908
rect 168837 7905 168849 7939
rect 168883 7936 168895 7939
rect 169754 7936 169760 7948
rect 168883 7908 169760 7936
rect 168883 7905 168895 7908
rect 168837 7899 168895 7905
rect 169754 7896 169760 7908
rect 169812 7896 169818 7948
rect 169864 7936 169892 7976
rect 171778 7964 171784 8016
rect 171836 8004 171842 8016
rect 182082 8004 182088 8016
rect 171836 7976 182088 8004
rect 171836 7964 171842 7976
rect 182082 7964 182088 7976
rect 182140 7964 182146 8016
rect 198734 7964 198740 8016
rect 198792 8004 198798 8016
rect 199378 8004 199384 8016
rect 198792 7976 199384 8004
rect 198792 7964 198798 7976
rect 199378 7964 199384 7976
rect 199436 8004 199442 8016
rect 211246 8004 211252 8016
rect 199436 7976 211252 8004
rect 199436 7964 199442 7976
rect 211246 7964 211252 7976
rect 211304 7964 211310 8016
rect 218974 7964 218980 8016
rect 219032 8004 219038 8016
rect 226058 8004 226064 8016
rect 219032 7976 226064 8004
rect 219032 7964 219038 7976
rect 226058 7964 226064 7976
rect 226116 7964 226122 8016
rect 226334 7964 226340 8016
rect 226392 8004 226398 8016
rect 256878 8004 256884 8016
rect 226392 7976 256884 8004
rect 226392 7964 226398 7976
rect 256878 7964 256884 7976
rect 256936 7964 256942 8016
rect 258718 7964 258724 8016
rect 258776 8004 258782 8016
rect 263226 8004 263232 8016
rect 258776 7976 263232 8004
rect 258776 7964 258782 7976
rect 263226 7964 263232 7976
rect 263284 7964 263290 8016
rect 213546 7936 213552 7948
rect 169864 7908 213552 7936
rect 213546 7896 213552 7908
rect 213604 7896 213610 7948
rect 223850 7896 223856 7948
rect 223908 7936 223914 7948
rect 255314 7936 255320 7948
rect 223908 7908 255320 7936
rect 223908 7896 223914 7908
rect 255314 7896 255320 7908
rect 255372 7896 255378 7948
rect 264072 7936 264100 8044
rect 264808 8004 264836 8044
rect 264882 8032 264888 8084
rect 264940 8072 264946 8084
rect 264977 8075 265035 8081
rect 264977 8072 264989 8075
rect 264940 8044 264989 8072
rect 264940 8032 264946 8044
rect 264977 8041 264989 8044
rect 265023 8041 265035 8075
rect 264977 8035 265035 8041
rect 265250 8032 265256 8084
rect 265308 8072 265314 8084
rect 266354 8072 266360 8084
rect 265308 8044 266360 8072
rect 265308 8032 265314 8044
rect 266354 8032 266360 8044
rect 266412 8032 266418 8084
rect 267461 8075 267519 8081
rect 266924 8044 267412 8072
rect 266924 8004 266952 8044
rect 264808 7976 266952 8004
rect 266998 7964 267004 8016
rect 267056 8004 267062 8016
rect 267384 8004 267412 8044
rect 267461 8041 267473 8075
rect 267507 8072 267519 8075
rect 267507 8044 268792 8072
rect 267507 8041 267519 8044
rect 267461 8035 267519 8041
rect 268010 8004 268016 8016
rect 267056 7976 267136 8004
rect 267384 7976 268016 8004
rect 267056 7964 267062 7976
rect 267108 7945 267136 7976
rect 268010 7964 268016 7976
rect 268068 7964 268074 8016
rect 268764 8004 268792 8044
rect 268838 8032 268844 8084
rect 268896 8032 268902 8084
rect 269574 8032 269580 8084
rect 269632 8072 269638 8084
rect 270034 8072 270040 8084
rect 269632 8044 270040 8072
rect 269632 8032 269638 8044
rect 270034 8032 270040 8044
rect 270092 8032 270098 8084
rect 271046 8072 271052 8084
rect 270144 8044 271052 8072
rect 270144 8004 270172 8044
rect 271046 8032 271052 8044
rect 271104 8032 271110 8084
rect 271138 8032 271144 8084
rect 271196 8072 271202 8084
rect 272150 8072 272156 8084
rect 271196 8044 272156 8072
rect 271196 8032 271202 8044
rect 272150 8032 272156 8044
rect 272208 8032 272214 8084
rect 268764 7976 270172 8004
rect 270221 8007 270279 8013
rect 270221 7973 270233 8007
rect 270267 8004 270279 8007
rect 270310 8004 270316 8016
rect 270267 7976 270316 8004
rect 270267 7973 270279 7976
rect 270221 7967 270279 7973
rect 270310 7964 270316 7976
rect 270368 7964 270374 8016
rect 267093 7939 267151 7945
rect 261036 7908 264100 7936
rect 264164 7908 265756 7936
rect 168009 7871 168067 7877
rect 168009 7837 168021 7871
rect 168055 7868 168067 7871
rect 168926 7868 168932 7880
rect 168055 7840 168932 7868
rect 168055 7837 168067 7840
rect 168009 7831 168067 7837
rect 168926 7828 168932 7840
rect 168984 7868 168990 7880
rect 169021 7871 169079 7877
rect 169021 7868 169033 7871
rect 168984 7840 169033 7868
rect 168984 7828 168990 7840
rect 169021 7837 169033 7840
rect 169067 7837 169079 7871
rect 169021 7831 169079 7837
rect 170582 7828 170588 7880
rect 170640 7868 170646 7880
rect 172606 7868 172612 7880
rect 170640 7840 172612 7868
rect 170640 7828 170646 7840
rect 172606 7828 172612 7840
rect 172664 7828 172670 7880
rect 202966 7828 202972 7880
rect 203024 7828 203030 7880
rect 211154 7828 211160 7880
rect 211212 7868 211218 7880
rect 219250 7868 219256 7880
rect 211212 7840 219256 7868
rect 211212 7828 211218 7840
rect 219250 7828 219256 7840
rect 219308 7828 219314 7880
rect 224034 7828 224040 7880
rect 224092 7868 224098 7880
rect 224092 7840 224954 7868
rect 224092 7828 224098 7840
rect 152056 7772 162072 7800
rect 152056 7760 152062 7772
rect 162118 7760 162124 7812
rect 162176 7800 162182 7812
rect 210326 7800 210332 7812
rect 162176 7772 210332 7800
rect 162176 7760 162182 7772
rect 210326 7760 210332 7772
rect 210384 7760 210390 7812
rect 213822 7760 213828 7812
rect 213880 7800 213886 7812
rect 213880 7772 222240 7800
rect 213880 7760 213886 7772
rect 34072 7704 41414 7732
rect 89714 7692 89720 7744
rect 89772 7692 89778 7744
rect 95970 7692 95976 7744
rect 96028 7732 96034 7744
rect 97813 7735 97871 7741
rect 97813 7732 97825 7735
rect 96028 7704 97825 7732
rect 96028 7692 96034 7704
rect 97813 7701 97825 7704
rect 97859 7701 97871 7735
rect 97813 7695 97871 7701
rect 97994 7692 98000 7744
rect 98052 7732 98058 7744
rect 109034 7732 109040 7744
rect 98052 7704 109040 7732
rect 98052 7692 98058 7704
rect 109034 7692 109040 7704
rect 109092 7692 109098 7744
rect 109129 7735 109187 7741
rect 109129 7701 109141 7735
rect 109175 7732 109187 7735
rect 109494 7732 109500 7744
rect 109175 7704 109500 7732
rect 109175 7701 109187 7704
rect 109129 7695 109187 7701
rect 109494 7692 109500 7704
rect 109552 7692 109558 7744
rect 114922 7692 114928 7744
rect 114980 7692 114986 7744
rect 115106 7692 115112 7744
rect 115164 7692 115170 7744
rect 115198 7692 115204 7744
rect 115256 7692 115262 7744
rect 115474 7692 115480 7744
rect 115532 7692 115538 7744
rect 151814 7692 151820 7744
rect 151872 7732 151878 7744
rect 158070 7732 158076 7744
rect 151872 7704 158076 7732
rect 151872 7692 151878 7704
rect 158070 7692 158076 7704
rect 158128 7692 158134 7744
rect 159358 7692 159364 7744
rect 159416 7732 159422 7744
rect 159453 7735 159511 7741
rect 159453 7732 159465 7735
rect 159416 7704 159465 7732
rect 159416 7692 159422 7704
rect 159453 7701 159465 7704
rect 159499 7701 159511 7735
rect 159453 7695 159511 7701
rect 165246 7692 165252 7744
rect 165304 7732 165310 7744
rect 165341 7735 165399 7741
rect 165341 7732 165353 7735
rect 165304 7704 165353 7732
rect 165304 7692 165310 7704
rect 165341 7701 165353 7704
rect 165387 7701 165399 7735
rect 165341 7695 165399 7701
rect 166534 7692 166540 7744
rect 166592 7732 166598 7744
rect 166813 7735 166871 7741
rect 166813 7732 166825 7735
rect 166592 7704 166825 7732
rect 166592 7692 166598 7704
rect 166813 7701 166825 7704
rect 166859 7701 166871 7735
rect 166813 7695 166871 7701
rect 169662 7692 169668 7744
rect 169720 7732 169726 7744
rect 189718 7732 189724 7744
rect 169720 7704 189724 7732
rect 169720 7692 169726 7704
rect 189718 7692 189724 7704
rect 189776 7692 189782 7744
rect 210418 7692 210424 7744
rect 210476 7732 210482 7744
rect 220814 7732 220820 7744
rect 210476 7704 220820 7732
rect 210476 7692 210482 7704
rect 220814 7692 220820 7704
rect 220872 7692 220878 7744
rect 222212 7732 222240 7772
rect 223666 7760 223672 7812
rect 223724 7800 223730 7812
rect 224405 7803 224463 7809
rect 224405 7800 224417 7803
rect 223724 7772 224417 7800
rect 223724 7760 223730 7772
rect 224405 7769 224417 7772
rect 224451 7800 224463 7803
rect 224770 7800 224776 7812
rect 224451 7772 224776 7800
rect 224451 7769 224463 7772
rect 224405 7763 224463 7769
rect 224770 7760 224776 7772
rect 224828 7760 224834 7812
rect 224926 7800 224954 7840
rect 225506 7828 225512 7880
rect 225564 7828 225570 7880
rect 227346 7828 227352 7880
rect 227404 7868 227410 7880
rect 234522 7868 234528 7880
rect 227404 7840 234528 7868
rect 227404 7828 227410 7840
rect 234522 7828 234528 7840
rect 234580 7828 234586 7880
rect 234706 7828 234712 7880
rect 234764 7828 234770 7880
rect 234798 7828 234804 7880
rect 234856 7868 234862 7880
rect 253106 7868 253112 7880
rect 234856 7840 253112 7868
rect 234856 7828 234862 7840
rect 253106 7828 253112 7840
rect 253164 7828 253170 7880
rect 261036 7877 261064 7908
rect 260377 7871 260435 7877
rect 260377 7837 260389 7871
rect 260423 7837 260435 7871
rect 260377 7831 260435 7837
rect 261021 7871 261079 7877
rect 261021 7837 261033 7871
rect 261067 7837 261079 7871
rect 261021 7831 261079 7837
rect 234430 7800 234436 7812
rect 224926 7772 234436 7800
rect 234430 7760 234436 7772
rect 234488 7760 234494 7812
rect 236638 7760 236644 7812
rect 236696 7800 236702 7812
rect 256970 7800 256976 7812
rect 236696 7772 256976 7800
rect 236696 7760 236702 7772
rect 256970 7760 256976 7772
rect 257028 7760 257034 7812
rect 259917 7803 259975 7809
rect 259917 7769 259929 7803
rect 259963 7800 259975 7803
rect 260392 7800 260420 7831
rect 261570 7828 261576 7880
rect 261628 7828 261634 7880
rect 262306 7828 262312 7880
rect 262364 7828 262370 7880
rect 263134 7828 263140 7880
rect 263192 7828 263198 7880
rect 263870 7828 263876 7880
rect 263928 7868 263934 7880
rect 264164 7877 264192 7908
rect 263965 7871 264023 7877
rect 263965 7868 263977 7871
rect 263928 7840 263977 7868
rect 263928 7828 263934 7840
rect 263965 7837 263977 7840
rect 264011 7837 264023 7871
rect 263965 7831 264023 7837
rect 264149 7871 264207 7877
rect 264149 7837 264161 7871
rect 264195 7837 264207 7871
rect 264149 7831 264207 7837
rect 264333 7871 264391 7877
rect 264333 7837 264345 7871
rect 264379 7868 264391 7871
rect 264793 7871 264851 7877
rect 264793 7868 264805 7871
rect 264379 7840 264805 7868
rect 264379 7837 264391 7840
rect 264333 7831 264391 7837
rect 264793 7837 264805 7840
rect 264839 7837 264851 7871
rect 264793 7831 264851 7837
rect 265618 7828 265624 7880
rect 265676 7828 265682 7880
rect 265728 7877 265756 7908
rect 267093 7905 267105 7939
rect 267139 7905 267151 7939
rect 267093 7899 267151 7905
rect 267734 7896 267740 7948
rect 267792 7936 267798 7948
rect 267792 7908 270816 7936
rect 267792 7896 267798 7908
rect 265713 7871 265771 7877
rect 265713 7837 265725 7871
rect 265759 7868 265771 7871
rect 267277 7871 267335 7877
rect 267277 7868 267289 7871
rect 265759 7840 267289 7868
rect 265759 7837 265771 7840
rect 265713 7831 265771 7837
rect 267277 7837 267289 7840
rect 267323 7868 267335 7871
rect 267550 7868 267556 7880
rect 267323 7840 267556 7868
rect 267323 7837 267335 7840
rect 267277 7831 267335 7837
rect 267550 7828 267556 7840
rect 267608 7828 267614 7880
rect 268013 7871 268071 7877
rect 268013 7837 268025 7871
rect 268059 7837 268071 7871
rect 268013 7831 268071 7837
rect 268105 7871 268163 7877
rect 268105 7837 268117 7871
rect 268151 7868 268163 7871
rect 268194 7868 268200 7880
rect 268151 7840 268200 7868
rect 268151 7837 268163 7840
rect 268105 7831 268163 7837
rect 264882 7800 264888 7812
rect 259963 7772 264888 7800
rect 259963 7769 259975 7772
rect 259917 7763 259975 7769
rect 264882 7760 264888 7772
rect 264940 7760 264946 7812
rect 268028 7800 268056 7831
rect 268194 7828 268200 7840
rect 268252 7868 268258 7880
rect 268378 7868 268384 7880
rect 268252 7840 268384 7868
rect 268252 7828 268258 7840
rect 268378 7828 268384 7840
rect 268436 7828 268442 7880
rect 268470 7828 268476 7880
rect 268528 7868 268534 7880
rect 268749 7871 268807 7877
rect 268749 7868 268761 7871
rect 268528 7840 268761 7868
rect 268528 7828 268534 7840
rect 268749 7837 268761 7840
rect 268795 7868 268807 7871
rect 268930 7868 268936 7880
rect 268795 7840 268936 7868
rect 268795 7837 268807 7840
rect 268749 7831 268807 7837
rect 268930 7828 268936 7840
rect 268988 7828 268994 7880
rect 269669 7871 269727 7877
rect 269669 7837 269681 7871
rect 269715 7837 269727 7871
rect 269669 7831 269727 7837
rect 265728 7772 268056 7800
rect 224497 7735 224555 7741
rect 224497 7732 224509 7735
rect 222212 7704 224509 7732
rect 224497 7701 224509 7704
rect 224543 7732 224555 7735
rect 224954 7732 224960 7744
rect 224543 7704 224960 7732
rect 224543 7701 224555 7704
rect 224497 7695 224555 7701
rect 224954 7692 224960 7704
rect 225012 7692 225018 7744
rect 225690 7692 225696 7744
rect 225748 7692 225754 7744
rect 234522 7692 234528 7744
rect 234580 7732 234586 7744
rect 234798 7732 234804 7744
rect 234580 7704 234804 7732
rect 234580 7692 234586 7704
rect 234798 7692 234804 7704
rect 234856 7692 234862 7744
rect 234890 7692 234896 7744
rect 234948 7692 234954 7744
rect 235810 7692 235816 7744
rect 235868 7692 235874 7744
rect 237190 7692 237196 7744
rect 237248 7732 237254 7744
rect 240134 7732 240140 7744
rect 237248 7704 240140 7732
rect 237248 7692 237254 7704
rect 240134 7692 240140 7704
rect 240192 7692 240198 7744
rect 248874 7692 248880 7744
rect 248932 7732 248938 7744
rect 249794 7732 249800 7744
rect 248932 7704 249800 7732
rect 248932 7692 248938 7704
rect 249794 7692 249800 7704
rect 249852 7692 249858 7744
rect 260193 7735 260251 7741
rect 260193 7701 260205 7735
rect 260239 7732 260251 7735
rect 262214 7732 262220 7744
rect 260239 7704 262220 7732
rect 260239 7701 260251 7704
rect 260193 7695 260251 7701
rect 262214 7692 262220 7704
rect 262272 7692 262278 7744
rect 262766 7692 262772 7744
rect 262824 7732 262830 7744
rect 265728 7732 265756 7772
rect 262824 7704 265756 7732
rect 265897 7735 265955 7741
rect 262824 7692 262830 7704
rect 265897 7701 265909 7735
rect 265943 7732 265955 7735
rect 265986 7732 265992 7744
rect 265943 7704 265992 7732
rect 265943 7701 265955 7704
rect 265897 7695 265955 7701
rect 265986 7692 265992 7704
rect 266044 7692 266050 7744
rect 268010 7692 268016 7744
rect 268068 7732 268074 7744
rect 268289 7735 268347 7741
rect 268289 7732 268301 7735
rect 268068 7704 268301 7732
rect 268068 7692 268074 7704
rect 268289 7701 268301 7704
rect 268335 7701 268347 7735
rect 268289 7695 268347 7701
rect 269206 7692 269212 7744
rect 269264 7692 269270 7744
rect 269684 7732 269712 7831
rect 269850 7828 269856 7880
rect 269908 7828 269914 7880
rect 270126 7877 270132 7880
rect 270089 7871 270132 7877
rect 270089 7837 270101 7871
rect 270089 7831 270132 7837
rect 270126 7828 270132 7831
rect 270184 7828 270190 7880
rect 270788 7877 270816 7908
rect 270773 7871 270831 7877
rect 270773 7837 270785 7871
rect 270819 7837 270831 7871
rect 270773 7831 270831 7837
rect 269945 7803 270003 7809
rect 269945 7769 269957 7803
rect 269991 7800 270003 7803
rect 270218 7800 270224 7812
rect 269991 7772 270224 7800
rect 269991 7769 270003 7772
rect 269945 7763 270003 7769
rect 270218 7760 270224 7772
rect 270276 7760 270282 7812
rect 270034 7732 270040 7744
rect 269684 7704 270040 7732
rect 270034 7692 270040 7704
rect 270092 7732 270098 7744
rect 270865 7735 270923 7741
rect 270865 7732 270877 7735
rect 270092 7704 270877 7732
rect 270092 7692 270098 7704
rect 270865 7701 270877 7704
rect 270911 7701 270923 7735
rect 270865 7695 270923 7701
rect 1104 7642 271651 7664
rect 1104 7590 68546 7642
rect 68598 7590 68610 7642
rect 68662 7590 68674 7642
rect 68726 7590 68738 7642
rect 68790 7590 68802 7642
rect 68854 7590 136143 7642
rect 136195 7590 136207 7642
rect 136259 7590 136271 7642
rect 136323 7590 136335 7642
rect 136387 7590 136399 7642
rect 136451 7590 203740 7642
rect 203792 7590 203804 7642
rect 203856 7590 203868 7642
rect 203920 7590 203932 7642
rect 203984 7590 203996 7642
rect 204048 7590 271337 7642
rect 271389 7590 271401 7642
rect 271453 7590 271465 7642
rect 271517 7590 271529 7642
rect 271581 7590 271593 7642
rect 271645 7590 271651 7642
rect 1104 7568 271651 7590
rect 4062 7488 4068 7540
rect 4120 7528 4126 7540
rect 24946 7528 24952 7540
rect 4120 7500 24952 7528
rect 4120 7488 4126 7500
rect 24946 7488 24952 7500
rect 25004 7488 25010 7540
rect 76374 7488 76380 7540
rect 76432 7488 76438 7540
rect 88518 7488 88524 7540
rect 88576 7528 88582 7540
rect 95694 7528 95700 7540
rect 88576 7500 95700 7528
rect 88576 7488 88582 7500
rect 95694 7488 95700 7500
rect 95752 7488 95758 7540
rect 95878 7488 95884 7540
rect 95936 7528 95942 7540
rect 100570 7528 100576 7540
rect 95936 7500 100576 7528
rect 95936 7488 95942 7500
rect 100570 7488 100576 7500
rect 100628 7488 100634 7540
rect 100754 7488 100760 7540
rect 100812 7528 100818 7540
rect 101309 7531 101367 7537
rect 101309 7528 101321 7531
rect 100812 7500 101321 7528
rect 100812 7488 100818 7500
rect 101309 7497 101321 7500
rect 101355 7497 101367 7531
rect 101309 7491 101367 7497
rect 107838 7488 107844 7540
rect 107896 7528 107902 7540
rect 110601 7531 110659 7537
rect 110601 7528 110613 7531
rect 107896 7500 110613 7528
rect 107896 7488 107902 7500
rect 110601 7497 110613 7500
rect 110647 7497 110659 7531
rect 110601 7491 110659 7497
rect 111518 7488 111524 7540
rect 111576 7488 111582 7540
rect 111610 7488 111616 7540
rect 111668 7528 111674 7540
rect 113082 7528 113088 7540
rect 111668 7500 113088 7528
rect 111668 7488 111674 7500
rect 113082 7488 113088 7500
rect 113140 7528 113146 7540
rect 113140 7500 113588 7528
rect 113140 7488 113146 7500
rect 24394 7420 24400 7472
rect 24452 7460 24458 7472
rect 42978 7460 42984 7472
rect 24452 7432 42984 7460
rect 24452 7420 24458 7432
rect 42978 7420 42984 7432
rect 43036 7420 43042 7472
rect 97258 7420 97264 7472
rect 97316 7460 97322 7472
rect 99190 7460 99196 7472
rect 97316 7432 99196 7460
rect 97316 7420 97322 7432
rect 99190 7420 99196 7432
rect 99248 7420 99254 7472
rect 99282 7420 99288 7472
rect 99340 7460 99346 7472
rect 104158 7460 104164 7472
rect 99340 7432 104164 7460
rect 99340 7420 99346 7432
rect 104158 7420 104164 7432
rect 104216 7420 104222 7472
rect 108850 7420 108856 7472
rect 108908 7460 108914 7472
rect 111536 7460 111564 7488
rect 113560 7460 113588 7500
rect 115290 7488 115296 7540
rect 115348 7488 115354 7540
rect 115382 7488 115388 7540
rect 115440 7488 115446 7540
rect 117498 7488 117504 7540
rect 117556 7488 117562 7540
rect 119893 7531 119951 7537
rect 119893 7497 119905 7531
rect 119939 7528 119951 7531
rect 120994 7528 121000 7540
rect 119939 7500 121000 7528
rect 119939 7497 119951 7500
rect 119893 7491 119951 7497
rect 120994 7488 121000 7500
rect 121052 7488 121058 7540
rect 151538 7528 151544 7540
rect 137986 7500 151544 7528
rect 116578 7460 116584 7472
rect 108908 7432 109816 7460
rect 111536 7432 112116 7460
rect 113560 7432 116584 7460
rect 108908 7420 108914 7432
rect 76558 7352 76564 7404
rect 76616 7352 76622 7404
rect 78766 7352 78772 7404
rect 78824 7352 78830 7404
rect 84194 7352 84200 7404
rect 84252 7392 84258 7404
rect 95878 7401 95884 7404
rect 94961 7395 95019 7401
rect 94961 7392 94973 7395
rect 84252 7364 94973 7392
rect 84252 7352 84258 7364
rect 94961 7361 94973 7364
rect 95007 7361 95019 7395
rect 94961 7355 95019 7361
rect 95835 7395 95884 7401
rect 95835 7361 95847 7395
rect 95881 7361 95884 7395
rect 95835 7355 95884 7361
rect 95878 7352 95884 7355
rect 95936 7352 95942 7404
rect 97350 7352 97356 7404
rect 97408 7352 97414 7404
rect 97534 7352 97540 7404
rect 97592 7352 97598 7404
rect 98641 7395 98699 7401
rect 98641 7361 98653 7395
rect 98687 7361 98699 7395
rect 98641 7355 98699 7361
rect 93946 7284 93952 7336
rect 94004 7324 94010 7336
rect 94777 7327 94835 7333
rect 94777 7324 94789 7327
rect 94004 7296 94789 7324
rect 94004 7284 94010 7296
rect 94777 7293 94789 7296
rect 94823 7293 94835 7327
rect 95697 7327 95755 7333
rect 95697 7324 95709 7327
rect 94777 7287 94835 7293
rect 95528 7296 95709 7324
rect 78953 7259 79011 7265
rect 78953 7256 78965 7259
rect 64846 7228 78965 7256
rect 33686 7148 33692 7200
rect 33744 7188 33750 7200
rect 64846 7188 64874 7228
rect 78953 7225 78965 7228
rect 78999 7225 79011 7259
rect 78953 7219 79011 7225
rect 93854 7216 93860 7268
rect 93912 7256 93918 7268
rect 95421 7259 95479 7265
rect 95421 7256 95433 7259
rect 93912 7228 95433 7256
rect 93912 7216 93918 7228
rect 95421 7225 95433 7228
rect 95467 7225 95479 7259
rect 95421 7219 95479 7225
rect 33744 7160 64874 7188
rect 95528 7188 95556 7296
rect 95697 7293 95709 7296
rect 95743 7293 95755 7327
rect 95697 7287 95755 7293
rect 95973 7327 96031 7333
rect 95973 7293 95985 7327
rect 96019 7324 96031 7327
rect 96154 7324 96160 7336
rect 96019 7296 96160 7324
rect 96019 7293 96031 7296
rect 95973 7287 96031 7293
rect 96154 7284 96160 7296
rect 96212 7284 96218 7336
rect 96522 7284 96528 7336
rect 96580 7324 96586 7336
rect 98546 7324 98552 7336
rect 96580 7296 98552 7324
rect 96580 7284 96586 7296
rect 98546 7284 98552 7296
rect 98604 7284 98610 7336
rect 98656 7324 98684 7355
rect 98730 7352 98736 7404
rect 98788 7392 98794 7404
rect 99469 7395 99527 7401
rect 99469 7392 99481 7395
rect 98788 7364 99481 7392
rect 98788 7352 98794 7364
rect 99469 7361 99481 7364
rect 99515 7361 99527 7395
rect 99469 7355 99527 7361
rect 100113 7395 100171 7401
rect 100113 7361 100125 7395
rect 100159 7392 100171 7395
rect 101398 7392 101404 7404
rect 100159 7364 101404 7392
rect 100159 7361 100171 7364
rect 100113 7355 100171 7361
rect 101398 7352 101404 7364
rect 101456 7352 101462 7404
rect 101490 7352 101496 7404
rect 101548 7352 101554 7404
rect 107102 7352 107108 7404
rect 107160 7352 107166 7404
rect 108393 7395 108451 7401
rect 108393 7361 108405 7395
rect 108439 7361 108451 7395
rect 108393 7355 108451 7361
rect 99006 7324 99012 7336
rect 98656 7296 99012 7324
rect 99006 7284 99012 7296
rect 99064 7284 99070 7336
rect 108408 7324 108436 7355
rect 109034 7352 109040 7404
rect 109092 7352 109098 7404
rect 109788 7401 109816 7432
rect 109773 7395 109831 7401
rect 109773 7361 109785 7395
rect 109819 7361 109831 7395
rect 109773 7355 109831 7361
rect 110690 7352 110696 7404
rect 110748 7392 110754 7404
rect 110785 7395 110843 7401
rect 110785 7392 110797 7395
rect 110748 7364 110797 7392
rect 110748 7352 110754 7364
rect 110785 7361 110797 7364
rect 110831 7361 110843 7395
rect 110785 7355 110843 7361
rect 111242 7352 111248 7404
rect 111300 7352 111306 7404
rect 111334 7352 111340 7404
rect 111392 7392 111398 7404
rect 112088 7401 112116 7432
rect 116578 7420 116584 7432
rect 116636 7420 116642 7472
rect 118510 7420 118516 7472
rect 118568 7460 118574 7472
rect 137986 7460 138014 7500
rect 151538 7488 151544 7500
rect 151596 7488 151602 7540
rect 152550 7488 152556 7540
rect 152608 7528 152614 7540
rect 162118 7528 162124 7540
rect 152608 7500 162124 7528
rect 152608 7488 152614 7500
rect 162118 7488 162124 7500
rect 162176 7488 162182 7540
rect 162394 7488 162400 7540
rect 162452 7528 162458 7540
rect 163133 7531 163191 7537
rect 163133 7528 163145 7531
rect 162452 7500 163145 7528
rect 162452 7488 162458 7500
rect 163133 7497 163145 7500
rect 163179 7497 163191 7531
rect 163133 7491 163191 7497
rect 166902 7488 166908 7540
rect 166960 7488 166966 7540
rect 168561 7531 168619 7537
rect 168561 7497 168573 7531
rect 168607 7528 168619 7531
rect 168650 7528 168656 7540
rect 168607 7500 168656 7528
rect 168607 7497 168619 7500
rect 168561 7491 168619 7497
rect 154666 7460 154672 7472
rect 118568 7432 138014 7460
rect 139872 7432 154672 7460
rect 118568 7420 118574 7432
rect 111889 7395 111947 7401
rect 111889 7392 111901 7395
rect 111392 7364 111901 7392
rect 111392 7352 111398 7364
rect 111889 7361 111901 7364
rect 111935 7361 111947 7395
rect 111889 7355 111947 7361
rect 112073 7395 112131 7401
rect 112073 7361 112085 7395
rect 112119 7361 112131 7395
rect 112073 7355 112131 7361
rect 112806 7352 112812 7404
rect 112864 7352 112870 7404
rect 113082 7352 113088 7404
rect 113140 7352 113146 7404
rect 115017 7395 115075 7401
rect 115017 7361 115029 7395
rect 115063 7392 115075 7395
rect 115198 7392 115204 7404
rect 115063 7364 115204 7392
rect 115063 7361 115075 7364
rect 115017 7355 115075 7361
rect 115198 7352 115204 7364
rect 115256 7392 115262 7404
rect 115566 7392 115572 7404
rect 115256 7364 115572 7392
rect 115256 7352 115262 7364
rect 115566 7352 115572 7364
rect 115624 7352 115630 7404
rect 116302 7352 116308 7404
rect 116360 7352 116366 7404
rect 116762 7352 116768 7404
rect 116820 7392 116826 7404
rect 117409 7395 117467 7401
rect 117409 7392 117421 7395
rect 116820 7364 117421 7392
rect 116820 7352 116826 7364
rect 117409 7361 117421 7364
rect 117455 7361 117467 7395
rect 117409 7355 117467 7361
rect 118050 7352 118056 7404
rect 118108 7352 118114 7404
rect 120074 7352 120080 7404
rect 120132 7352 120138 7404
rect 124214 7352 124220 7404
rect 124272 7392 124278 7404
rect 124766 7392 124772 7404
rect 124272 7364 124772 7392
rect 124272 7352 124278 7364
rect 124766 7352 124772 7364
rect 124824 7392 124830 7404
rect 139872 7392 139900 7432
rect 154666 7420 154672 7432
rect 154724 7420 154730 7472
rect 162305 7463 162363 7469
rect 162305 7429 162317 7463
rect 162351 7460 162363 7463
rect 168576 7460 168604 7491
rect 168650 7488 168656 7500
rect 168708 7488 168714 7540
rect 179414 7488 179420 7540
rect 179472 7528 179478 7540
rect 210418 7528 210424 7540
rect 179472 7500 210424 7528
rect 179472 7488 179478 7500
rect 210418 7488 210424 7500
rect 210476 7488 210482 7540
rect 221458 7488 221464 7540
rect 221516 7488 221522 7540
rect 221918 7488 221924 7540
rect 221976 7528 221982 7540
rect 224678 7528 224684 7540
rect 221976 7500 224684 7528
rect 221976 7488 221982 7500
rect 224678 7488 224684 7500
rect 224736 7488 224742 7540
rect 227346 7528 227352 7540
rect 225432 7500 227352 7528
rect 210510 7460 210516 7472
rect 162351 7432 168604 7460
rect 176626 7432 210516 7460
rect 162351 7429 162363 7432
rect 162305 7423 162363 7429
rect 151722 7392 151728 7404
rect 124824 7364 139900 7392
rect 147646 7364 151728 7392
rect 124824 7352 124830 7364
rect 109126 7324 109132 7336
rect 108408 7296 109132 7324
rect 109126 7284 109132 7296
rect 109184 7284 109190 7336
rect 112947 7327 113005 7333
rect 112947 7293 112959 7327
rect 112993 7324 113005 7327
rect 112993 7296 115060 7324
rect 112993 7293 113005 7296
rect 112947 7287 113005 7293
rect 99098 7256 99104 7268
rect 96540 7228 99104 7256
rect 96540 7188 96568 7228
rect 99098 7216 99104 7228
rect 99156 7216 99162 7268
rect 99466 7216 99472 7268
rect 99524 7256 99530 7268
rect 106921 7259 106979 7265
rect 106921 7256 106933 7259
rect 99524 7228 106933 7256
rect 99524 7216 99530 7228
rect 106921 7225 106933 7228
rect 106967 7225 106979 7259
rect 106921 7219 106979 7225
rect 108853 7259 108911 7265
rect 108853 7225 108865 7259
rect 108899 7256 108911 7259
rect 109770 7256 109776 7268
rect 108899 7228 109776 7256
rect 108899 7225 108911 7228
rect 108853 7219 108911 7225
rect 109770 7216 109776 7228
rect 109828 7216 109834 7268
rect 112530 7216 112536 7268
rect 112588 7216 112594 7268
rect 115032 7256 115060 7296
rect 115106 7284 115112 7336
rect 115164 7324 115170 7336
rect 115474 7324 115480 7336
rect 115164 7296 115480 7324
rect 115164 7284 115170 7296
rect 115474 7284 115480 7296
rect 115532 7284 115538 7336
rect 117682 7324 117688 7336
rect 115584 7296 117688 7324
rect 115584 7256 115612 7296
rect 117682 7284 117688 7296
rect 117740 7284 117746 7336
rect 139210 7284 139216 7336
rect 139268 7324 139274 7336
rect 147646 7324 147674 7364
rect 151722 7352 151728 7364
rect 151780 7352 151786 7404
rect 151814 7352 151820 7404
rect 151872 7352 151878 7404
rect 152734 7352 152740 7404
rect 152792 7352 152798 7404
rect 160462 7392 160468 7404
rect 152844 7364 160468 7392
rect 139268 7296 147674 7324
rect 139268 7284 139274 7296
rect 151630 7284 151636 7336
rect 151688 7324 151694 7336
rect 152001 7327 152059 7333
rect 152001 7324 152013 7327
rect 151688 7296 152013 7324
rect 151688 7284 151694 7296
rect 152001 7293 152013 7296
rect 152047 7293 152059 7327
rect 152001 7287 152059 7293
rect 113468 7228 113864 7256
rect 115032 7228 115612 7256
rect 95528 7160 96568 7188
rect 96617 7191 96675 7197
rect 33744 7148 33750 7160
rect 96617 7157 96629 7191
rect 96663 7188 96675 7191
rect 97074 7188 97080 7200
rect 96663 7160 97080 7188
rect 96663 7157 96675 7160
rect 96617 7151 96675 7157
rect 97074 7148 97080 7160
rect 97132 7148 97138 7200
rect 97442 7148 97448 7200
rect 97500 7148 97506 7200
rect 97718 7148 97724 7200
rect 97776 7148 97782 7200
rect 97810 7148 97816 7200
rect 97868 7188 97874 7200
rect 98457 7191 98515 7197
rect 98457 7188 98469 7191
rect 97868 7160 98469 7188
rect 97868 7148 97874 7160
rect 98457 7157 98469 7160
rect 98503 7157 98515 7191
rect 98457 7151 98515 7157
rect 99282 7148 99288 7200
rect 99340 7148 99346 7200
rect 99926 7148 99932 7200
rect 99984 7148 99990 7200
rect 100570 7148 100576 7200
rect 100628 7188 100634 7200
rect 103422 7188 103428 7200
rect 100628 7160 103428 7188
rect 100628 7148 100634 7160
rect 103422 7148 103428 7160
rect 103480 7148 103486 7200
rect 103882 7148 103888 7200
rect 103940 7188 103946 7200
rect 108209 7191 108267 7197
rect 108209 7188 108221 7191
rect 103940 7160 108221 7188
rect 103940 7148 103946 7160
rect 108209 7157 108221 7160
rect 108255 7157 108267 7191
rect 108209 7151 108267 7157
rect 109218 7148 109224 7200
rect 109276 7188 109282 7200
rect 109589 7191 109647 7197
rect 109589 7188 109601 7191
rect 109276 7160 109601 7188
rect 109276 7148 109282 7160
rect 109589 7157 109601 7160
rect 109635 7157 109647 7191
rect 109589 7151 109647 7157
rect 111058 7148 111064 7200
rect 111116 7148 111122 7200
rect 113266 7148 113272 7200
rect 113324 7188 113330 7200
rect 113468 7188 113496 7228
rect 113324 7160 113496 7188
rect 113324 7148 113330 7160
rect 113726 7148 113732 7200
rect 113784 7148 113790 7200
rect 113836 7188 113864 7228
rect 115658 7216 115664 7268
rect 115716 7216 115722 7268
rect 118602 7256 118608 7268
rect 115768 7228 118608 7256
rect 115768 7188 115796 7228
rect 118602 7216 118608 7228
rect 118660 7216 118666 7268
rect 149330 7216 149336 7268
rect 149388 7256 149394 7268
rect 152844 7256 152872 7364
rect 160462 7352 160468 7364
rect 160520 7352 160526 7404
rect 161290 7352 161296 7404
rect 161348 7392 161354 7404
rect 162489 7395 162547 7401
rect 162489 7392 162501 7395
rect 161348 7364 162501 7392
rect 161348 7352 161354 7364
rect 162489 7361 162501 7364
rect 162535 7361 162547 7395
rect 162489 7355 162547 7361
rect 162946 7352 162952 7404
rect 163004 7352 163010 7404
rect 166718 7352 166724 7404
rect 166776 7352 166782 7404
rect 168745 7395 168803 7401
rect 168745 7361 168757 7395
rect 168791 7392 168803 7395
rect 169018 7392 169024 7404
rect 168791 7364 169024 7392
rect 168791 7361 168803 7364
rect 168745 7355 168803 7361
rect 169018 7352 169024 7364
rect 169076 7352 169082 7404
rect 154666 7284 154672 7336
rect 154724 7324 154730 7336
rect 171778 7324 171784 7336
rect 154724 7296 171784 7324
rect 154724 7284 154730 7296
rect 171778 7284 171784 7296
rect 171836 7284 171842 7336
rect 149388 7228 152872 7256
rect 149388 7216 149394 7228
rect 153654 7216 153660 7268
rect 153712 7256 153718 7268
rect 176626 7256 176654 7432
rect 210510 7420 210516 7432
rect 210568 7420 210574 7472
rect 211430 7420 211436 7472
rect 211488 7460 211494 7472
rect 219158 7460 219164 7472
rect 211488 7432 219164 7460
rect 211488 7420 211494 7432
rect 219158 7420 219164 7432
rect 219216 7420 219222 7472
rect 219250 7420 219256 7472
rect 219308 7460 219314 7472
rect 223574 7460 223580 7472
rect 219308 7432 223580 7460
rect 219308 7420 219314 7432
rect 223574 7420 223580 7432
rect 223632 7420 223638 7472
rect 225432 7460 225460 7500
rect 227346 7488 227352 7500
rect 227404 7488 227410 7540
rect 227530 7488 227536 7540
rect 227588 7528 227594 7540
rect 256786 7528 256792 7540
rect 227588 7500 256792 7528
rect 227588 7488 227594 7500
rect 256786 7488 256792 7500
rect 256844 7488 256850 7540
rect 261481 7531 261539 7537
rect 261481 7497 261493 7531
rect 261527 7497 261539 7531
rect 261481 7491 261539 7497
rect 262125 7531 262183 7537
rect 262125 7497 262137 7531
rect 262171 7528 262183 7531
rect 262398 7528 262404 7540
rect 262171 7500 262404 7528
rect 262171 7497 262183 7500
rect 262125 7491 262183 7497
rect 223960 7432 225460 7460
rect 213454 7352 213460 7404
rect 213512 7352 213518 7404
rect 216858 7352 216864 7404
rect 216916 7392 216922 7404
rect 223960 7401 223988 7432
rect 225506 7420 225512 7472
rect 225564 7460 225570 7472
rect 226337 7463 226395 7469
rect 226337 7460 226349 7463
rect 225564 7432 226349 7460
rect 225564 7420 225570 7432
rect 226337 7429 226349 7432
rect 226383 7429 226395 7463
rect 226337 7423 226395 7429
rect 229738 7420 229744 7472
rect 229796 7460 229802 7472
rect 249610 7460 249616 7472
rect 229796 7432 249616 7460
rect 229796 7420 229802 7432
rect 249610 7420 249616 7432
rect 249668 7420 249674 7472
rect 252094 7420 252100 7472
rect 252152 7420 252158 7472
rect 252204 7432 252968 7460
rect 218517 7395 218575 7401
rect 218517 7392 218529 7395
rect 216916 7364 218529 7392
rect 216916 7352 216922 7364
rect 218517 7361 218529 7364
rect 218563 7361 218575 7395
rect 218517 7355 218575 7361
rect 221645 7395 221703 7401
rect 221645 7361 221657 7395
rect 221691 7361 221703 7395
rect 221645 7355 221703 7361
rect 223945 7395 224003 7401
rect 223945 7361 223957 7395
rect 223991 7361 224003 7395
rect 223945 7355 224003 7361
rect 213362 7284 213368 7336
rect 213420 7324 213426 7336
rect 213641 7327 213699 7333
rect 213641 7324 213653 7327
rect 213420 7296 213653 7324
rect 213420 7284 213426 7296
rect 213641 7293 213653 7296
rect 213687 7293 213699 7327
rect 213641 7287 213699 7293
rect 217962 7284 217968 7336
rect 218020 7324 218026 7336
rect 221660 7324 221688 7355
rect 224586 7352 224592 7404
rect 224644 7352 224650 7404
rect 225969 7395 226027 7401
rect 225969 7392 225981 7395
rect 224880 7364 225981 7392
rect 224880 7324 224908 7364
rect 225969 7361 225981 7364
rect 226015 7361 226027 7395
rect 225969 7355 226027 7361
rect 234430 7352 234436 7404
rect 234488 7392 234494 7404
rect 236638 7392 236644 7404
rect 234488 7364 236644 7392
rect 234488 7352 234494 7364
rect 236638 7352 236644 7364
rect 236696 7352 236702 7404
rect 250165 7395 250223 7401
rect 250165 7361 250177 7395
rect 250211 7392 250223 7395
rect 250993 7395 251051 7401
rect 250993 7392 251005 7395
rect 250211 7364 251005 7392
rect 250211 7361 250223 7364
rect 250165 7355 250223 7361
rect 250993 7361 251005 7364
rect 251039 7392 251051 7395
rect 251450 7392 251456 7404
rect 251039 7364 251456 7392
rect 251039 7361 251051 7364
rect 250993 7355 251051 7361
rect 251450 7352 251456 7364
rect 251508 7392 251514 7404
rect 251913 7395 251971 7401
rect 251913 7392 251925 7395
rect 251508 7364 251925 7392
rect 251508 7352 251514 7364
rect 251913 7361 251925 7364
rect 251959 7392 251971 7395
rect 252204 7392 252232 7432
rect 251959 7364 252232 7392
rect 251959 7361 251971 7364
rect 251913 7355 251971 7361
rect 252830 7352 252836 7404
rect 252888 7352 252894 7404
rect 252940 7401 252968 7432
rect 253106 7420 253112 7472
rect 253164 7420 253170 7472
rect 261496 7460 261524 7491
rect 262398 7488 262404 7500
rect 262456 7488 262462 7540
rect 262766 7488 262772 7540
rect 262824 7488 262830 7540
rect 263410 7488 263416 7540
rect 263468 7488 263474 7540
rect 264330 7488 264336 7540
rect 264388 7488 264394 7540
rect 265342 7488 265348 7540
rect 265400 7528 265406 7540
rect 265437 7531 265495 7537
rect 265437 7528 265449 7531
rect 265400 7500 265449 7528
rect 265400 7488 265406 7500
rect 265437 7497 265449 7500
rect 265483 7497 265495 7531
rect 265437 7491 265495 7497
rect 266170 7488 266176 7540
rect 266228 7488 266234 7540
rect 268028 7500 268424 7528
rect 267918 7460 267924 7472
rect 261496 7432 262904 7460
rect 252925 7395 252983 7401
rect 252925 7361 252937 7395
rect 252971 7392 252983 7395
rect 253198 7392 253204 7404
rect 252971 7364 253204 7392
rect 252971 7361 252983 7364
rect 252925 7355 252983 7361
rect 253198 7352 253204 7364
rect 253256 7352 253262 7404
rect 260377 7395 260435 7401
rect 260377 7361 260389 7395
rect 260423 7361 260435 7395
rect 260377 7355 260435 7361
rect 260837 7395 260895 7401
rect 260837 7361 260849 7395
rect 260883 7392 260895 7395
rect 261570 7392 261576 7404
rect 260883 7364 261576 7392
rect 260883 7361 260895 7364
rect 260837 7355 260895 7361
rect 218020 7296 221688 7324
rect 223776 7296 224908 7324
rect 218020 7284 218026 7296
rect 214282 7256 214288 7268
rect 153712 7228 176654 7256
rect 195946 7228 214288 7256
rect 153712 7216 153718 7228
rect 113836 7160 115796 7188
rect 116394 7148 116400 7200
rect 116452 7188 116458 7200
rect 116578 7188 116584 7200
rect 116452 7160 116584 7188
rect 116452 7148 116458 7160
rect 116578 7148 116584 7160
rect 116636 7188 116642 7200
rect 117130 7188 117136 7200
rect 116636 7160 117136 7188
rect 116636 7148 116642 7160
rect 117130 7148 117136 7160
rect 117188 7148 117194 7200
rect 118142 7148 118148 7200
rect 118200 7148 118206 7200
rect 119430 7148 119436 7200
rect 119488 7188 119494 7200
rect 146294 7188 146300 7200
rect 119488 7160 146300 7188
rect 119488 7148 119494 7160
rect 146294 7148 146300 7160
rect 146352 7148 146358 7200
rect 146386 7148 146392 7200
rect 146444 7188 146450 7200
rect 151446 7188 151452 7200
rect 146444 7160 151452 7188
rect 146444 7148 146450 7160
rect 151446 7148 151452 7160
rect 151504 7148 151510 7200
rect 152182 7148 152188 7200
rect 152240 7188 152246 7200
rect 152921 7191 152979 7197
rect 152921 7188 152933 7191
rect 152240 7160 152933 7188
rect 152240 7148 152246 7160
rect 152921 7157 152933 7160
rect 152967 7157 152979 7191
rect 152921 7151 152979 7157
rect 172514 7148 172520 7200
rect 172572 7188 172578 7200
rect 195946 7188 195974 7228
rect 214282 7216 214288 7228
rect 214340 7256 214346 7268
rect 218701 7259 218759 7265
rect 214340 7228 215432 7256
rect 214340 7216 214346 7228
rect 172572 7160 195974 7188
rect 172572 7148 172578 7160
rect 210418 7148 210424 7200
rect 210476 7188 210482 7200
rect 215294 7188 215300 7200
rect 210476 7160 215300 7188
rect 210476 7148 210482 7160
rect 215294 7148 215300 7160
rect 215352 7148 215358 7200
rect 215404 7188 215432 7228
rect 218701 7225 218713 7259
rect 218747 7256 218759 7259
rect 219434 7256 219440 7268
rect 218747 7228 219440 7256
rect 218747 7225 218759 7228
rect 218701 7219 218759 7225
rect 219434 7216 219440 7228
rect 219492 7216 219498 7268
rect 223776 7265 223804 7296
rect 225046 7284 225052 7336
rect 225104 7284 225110 7336
rect 249978 7284 249984 7336
rect 250036 7284 250042 7336
rect 250809 7327 250867 7333
rect 250809 7293 250821 7327
rect 250855 7293 250867 7327
rect 250809 7287 250867 7293
rect 223761 7259 223819 7265
rect 223761 7225 223773 7259
rect 223807 7225 223819 7259
rect 250824 7256 250852 7287
rect 251174 7284 251180 7336
rect 251232 7284 251238 7336
rect 251729 7327 251787 7333
rect 251729 7293 251741 7327
rect 251775 7293 251787 7327
rect 260392 7324 260420 7355
rect 261570 7352 261576 7364
rect 261628 7352 261634 7404
rect 261662 7352 261668 7404
rect 261720 7352 261726 7404
rect 262306 7352 262312 7404
rect 262364 7352 262370 7404
rect 261205 7327 261263 7333
rect 260392 7296 261156 7324
rect 251729 7287 251787 7293
rect 251634 7256 251640 7268
rect 250824 7228 251640 7256
rect 223761 7219 223819 7225
rect 251634 7216 251640 7228
rect 251692 7216 251698 7268
rect 251744 7256 251772 7287
rect 260653 7259 260711 7265
rect 260653 7256 260665 7259
rect 251744 7228 260665 7256
rect 260653 7225 260665 7228
rect 260699 7225 260711 7259
rect 261128 7256 261156 7296
rect 261205 7293 261217 7327
rect 261251 7324 261263 7327
rect 261680 7324 261708 7352
rect 261251 7296 261708 7324
rect 261251 7293 261263 7296
rect 261205 7287 261263 7293
rect 262876 7256 262904 7432
rect 262968 7432 267924 7460
rect 262968 7401 262996 7432
rect 267918 7420 267924 7432
rect 267976 7420 267982 7472
rect 262953 7395 263011 7401
rect 262953 7361 262965 7395
rect 262999 7361 263011 7395
rect 262953 7355 263011 7361
rect 263597 7395 263655 7401
rect 263597 7361 263609 7395
rect 263643 7392 263655 7395
rect 264054 7392 264060 7404
rect 263643 7364 264060 7392
rect 263643 7361 263655 7364
rect 263597 7355 263655 7361
rect 264054 7352 264060 7364
rect 264112 7352 264118 7404
rect 264146 7352 264152 7404
rect 264204 7352 264210 7404
rect 264330 7352 264336 7404
rect 264388 7392 264394 7404
rect 264790 7392 264796 7404
rect 264388 7364 264796 7392
rect 264388 7352 264394 7364
rect 264790 7352 264796 7364
rect 264848 7352 264854 7404
rect 265250 7352 265256 7404
rect 265308 7352 265314 7404
rect 265986 7352 265992 7404
rect 266044 7401 266050 7404
rect 266044 7392 266053 7401
rect 266044 7364 266089 7392
rect 266044 7355 266053 7364
rect 266044 7352 266050 7355
rect 267274 7352 267280 7404
rect 267332 7352 267338 7404
rect 268028 7392 268056 7500
rect 267844 7364 268056 7392
rect 268105 7395 268163 7401
rect 267090 7284 267096 7336
rect 267148 7284 267154 7336
rect 267844 7324 267872 7364
rect 268105 7361 268117 7395
rect 268151 7390 268163 7395
rect 268194 7390 268200 7404
rect 268151 7362 268200 7390
rect 268151 7361 268163 7362
rect 268105 7355 268163 7361
rect 268194 7352 268200 7362
rect 268252 7352 268258 7404
rect 267200 7296 267872 7324
rect 267921 7327 267979 7333
rect 267200 7256 267228 7296
rect 267921 7293 267933 7327
rect 267967 7324 267979 7327
rect 268396 7324 268424 7500
rect 268470 7488 268476 7540
rect 268528 7528 268534 7540
rect 270310 7528 270316 7540
rect 268528 7500 270316 7528
rect 268528 7488 268534 7500
rect 270310 7488 270316 7500
rect 270368 7488 270374 7540
rect 270678 7488 270684 7540
rect 270736 7528 270742 7540
rect 270865 7531 270923 7537
rect 270865 7528 270877 7531
rect 270736 7500 270877 7528
rect 270736 7488 270742 7500
rect 270865 7497 270877 7500
rect 270911 7497 270923 7531
rect 270865 7491 270923 7497
rect 271138 7488 271144 7540
rect 271196 7528 271202 7540
rect 272150 7528 272156 7540
rect 271196 7500 272156 7528
rect 271196 7488 271202 7500
rect 272150 7488 272156 7500
rect 272208 7488 272214 7540
rect 268838 7420 268844 7472
rect 268896 7460 268902 7472
rect 269853 7463 269911 7469
rect 268896 7432 269713 7460
rect 268896 7420 268902 7432
rect 269574 7401 269580 7404
rect 269565 7395 269580 7401
rect 269565 7361 269577 7395
rect 269565 7355 269580 7361
rect 269574 7352 269580 7355
rect 269632 7352 269638 7404
rect 269685 7401 269713 7432
rect 269853 7429 269865 7463
rect 269899 7460 269911 7463
rect 270402 7460 270408 7472
rect 269899 7432 270408 7460
rect 269899 7429 269911 7432
rect 269853 7423 269911 7429
rect 270402 7420 270408 7432
rect 270460 7420 270466 7472
rect 269670 7395 269728 7401
rect 269670 7361 269682 7395
rect 269716 7361 269728 7395
rect 269670 7355 269728 7361
rect 269758 7352 269764 7404
rect 269816 7392 269822 7404
rect 269945 7395 270003 7401
rect 269945 7392 269957 7395
rect 269816 7364 269957 7392
rect 269816 7352 269822 7364
rect 269945 7361 269957 7364
rect 269991 7361 270003 7395
rect 269945 7355 270003 7361
rect 270083 7395 270141 7401
rect 270083 7361 270095 7395
rect 270129 7392 270141 7395
rect 270696 7392 270724 7488
rect 270129 7364 270724 7392
rect 270773 7395 270831 7401
rect 270129 7361 270141 7364
rect 270083 7355 270141 7361
rect 270773 7361 270785 7395
rect 270819 7361 270831 7395
rect 270773 7355 270831 7361
rect 270788 7324 270816 7355
rect 267967 7296 268148 7324
rect 268396 7296 270816 7324
rect 267967 7293 267979 7296
rect 267921 7287 267979 7293
rect 261128 7228 262260 7256
rect 262876 7228 267228 7256
rect 268120 7256 268148 7296
rect 270770 7256 270776 7268
rect 268120 7228 270776 7256
rect 260653 7219 260711 7225
rect 223666 7188 223672 7200
rect 215404 7160 223672 7188
rect 223666 7148 223672 7160
rect 223724 7148 223730 7200
rect 224586 7148 224592 7200
rect 224644 7188 224650 7200
rect 226978 7188 226984 7200
rect 224644 7160 226984 7188
rect 224644 7148 224650 7160
rect 226978 7148 226984 7160
rect 227036 7148 227042 7200
rect 248414 7148 248420 7200
rect 248472 7188 248478 7200
rect 250349 7191 250407 7197
rect 250349 7188 250361 7191
rect 248472 7160 250361 7188
rect 248472 7148 248478 7160
rect 250349 7157 250361 7160
rect 250395 7157 250407 7191
rect 250349 7151 250407 7157
rect 252830 7148 252836 7200
rect 252888 7188 252894 7200
rect 260193 7191 260251 7197
rect 260193 7188 260205 7191
rect 252888 7160 260205 7188
rect 252888 7148 252894 7160
rect 260193 7157 260205 7160
rect 260239 7157 260251 7191
rect 262232 7188 262260 7228
rect 270770 7216 270776 7228
rect 270828 7216 270834 7268
rect 266262 7188 266268 7200
rect 262232 7160 266268 7188
rect 260193 7151 260251 7157
rect 266262 7148 266268 7160
rect 266320 7148 266326 7200
rect 266906 7148 266912 7200
rect 266964 7188 266970 7200
rect 267461 7191 267519 7197
rect 267461 7188 267473 7191
rect 266964 7160 267473 7188
rect 266964 7148 266970 7160
rect 267461 7157 267473 7160
rect 267507 7157 267519 7191
rect 267461 7151 267519 7157
rect 267826 7148 267832 7200
rect 267884 7188 267890 7200
rect 268289 7191 268347 7197
rect 268289 7188 268301 7191
rect 267884 7160 268301 7188
rect 267884 7148 267890 7160
rect 268289 7157 268301 7160
rect 268335 7157 268347 7191
rect 268289 7151 268347 7157
rect 269114 7148 269120 7200
rect 269172 7188 269178 7200
rect 270221 7191 270279 7197
rect 270221 7188 270233 7191
rect 269172 7160 270233 7188
rect 269172 7148 269178 7160
rect 270221 7157 270233 7160
rect 270267 7157 270279 7191
rect 270221 7151 270279 7157
rect 1104 7098 271492 7120
rect 1104 7046 34748 7098
rect 34800 7046 34812 7098
rect 34864 7046 34876 7098
rect 34928 7046 34940 7098
rect 34992 7046 35004 7098
rect 35056 7046 102345 7098
rect 102397 7046 102409 7098
rect 102461 7046 102473 7098
rect 102525 7046 102537 7098
rect 102589 7046 102601 7098
rect 102653 7046 169942 7098
rect 169994 7046 170006 7098
rect 170058 7046 170070 7098
rect 170122 7046 170134 7098
rect 170186 7046 170198 7098
rect 170250 7046 237539 7098
rect 237591 7046 237603 7098
rect 237655 7046 237667 7098
rect 237719 7046 237731 7098
rect 237783 7046 237795 7098
rect 237847 7046 271492 7098
rect 1104 7024 271492 7046
rect 93578 6944 93584 6996
rect 93636 6984 93642 6996
rect 96522 6984 96528 6996
rect 93636 6956 96528 6984
rect 93636 6944 93642 6956
rect 96522 6944 96528 6956
rect 96580 6944 96586 6996
rect 97629 6987 97687 6993
rect 97629 6953 97641 6987
rect 97675 6953 97687 6987
rect 97629 6947 97687 6953
rect 95510 6876 95516 6928
rect 95568 6916 95574 6928
rect 96154 6916 96160 6928
rect 95568 6888 96160 6916
rect 95568 6876 95574 6888
rect 96154 6876 96160 6888
rect 96212 6876 96218 6928
rect 97166 6916 97172 6928
rect 96586 6888 97172 6916
rect 19242 6808 19248 6860
rect 19300 6848 19306 6860
rect 24762 6848 24768 6860
rect 19300 6820 24768 6848
rect 19300 6808 19306 6820
rect 24762 6808 24768 6820
rect 24820 6808 24826 6860
rect 30466 6808 30472 6860
rect 30524 6848 30530 6860
rect 40862 6848 40868 6860
rect 30524 6820 40868 6848
rect 30524 6808 30530 6820
rect 40862 6808 40868 6820
rect 40920 6808 40926 6860
rect 95234 6808 95240 6860
rect 95292 6848 95298 6860
rect 96586 6848 96614 6888
rect 97166 6876 97172 6888
rect 97224 6876 97230 6928
rect 97644 6916 97672 6947
rect 97994 6944 98000 6996
rect 98052 6984 98058 6996
rect 98273 6987 98331 6993
rect 98273 6984 98285 6987
rect 98052 6956 98285 6984
rect 98052 6944 98058 6956
rect 98273 6953 98285 6956
rect 98319 6984 98331 6987
rect 100481 6987 100539 6993
rect 100481 6984 100493 6987
rect 98319 6956 100493 6984
rect 98319 6953 98331 6956
rect 98273 6947 98331 6953
rect 100481 6953 100493 6956
rect 100527 6984 100539 6987
rect 100938 6984 100944 6996
rect 100527 6956 100944 6984
rect 100527 6953 100539 6956
rect 100481 6947 100539 6953
rect 100938 6944 100944 6956
rect 100996 6944 101002 6996
rect 106366 6944 106372 6996
rect 106424 6984 106430 6996
rect 108390 6984 108396 6996
rect 106424 6956 108396 6984
rect 106424 6944 106430 6956
rect 108390 6944 108396 6956
rect 108448 6944 108454 6996
rect 108758 6944 108764 6996
rect 108816 6944 108822 6996
rect 108945 6987 109003 6993
rect 108945 6953 108957 6987
rect 108991 6984 109003 6987
rect 109034 6984 109040 6996
rect 108991 6956 109040 6984
rect 108991 6953 109003 6956
rect 108945 6947 109003 6953
rect 109034 6944 109040 6956
rect 109092 6944 109098 6996
rect 110230 6944 110236 6996
rect 110288 6984 110294 6996
rect 110325 6987 110383 6993
rect 110325 6984 110337 6987
rect 110288 6956 110337 6984
rect 110288 6944 110294 6956
rect 110325 6953 110337 6956
rect 110371 6984 110383 6987
rect 110371 6956 112300 6984
rect 110371 6953 110383 6956
rect 110325 6947 110383 6953
rect 97902 6916 97908 6928
rect 97644 6888 97908 6916
rect 97902 6876 97908 6888
rect 97960 6916 97966 6928
rect 106185 6919 106243 6925
rect 97960 6888 100524 6916
rect 97960 6876 97966 6888
rect 95292 6820 96614 6848
rect 95292 6808 95298 6820
rect 96982 6808 96988 6860
rect 97040 6848 97046 6860
rect 97040 6820 97396 6848
rect 97040 6808 97046 6820
rect 97368 6792 97396 6820
rect 97534 6808 97540 6860
rect 97592 6848 97598 6860
rect 97592 6820 98960 6848
rect 97592 6808 97598 6820
rect 24578 6740 24584 6792
rect 24636 6780 24642 6792
rect 38838 6780 38844 6792
rect 24636 6752 38844 6780
rect 24636 6740 24642 6752
rect 38838 6740 38844 6752
rect 38896 6740 38902 6792
rect 39114 6740 39120 6792
rect 39172 6780 39178 6792
rect 55858 6780 55864 6792
rect 39172 6752 55864 6780
rect 39172 6740 39178 6752
rect 55858 6740 55864 6752
rect 55916 6740 55922 6792
rect 94498 6780 94504 6792
rect 60706 6752 94504 6780
rect 20806 6672 20812 6724
rect 20864 6712 20870 6724
rect 43990 6712 43996 6724
rect 20864 6684 43996 6712
rect 20864 6672 20870 6684
rect 43990 6672 43996 6684
rect 44048 6672 44054 6724
rect 46658 6672 46664 6724
rect 46716 6712 46722 6724
rect 60706 6712 60734 6752
rect 94498 6740 94504 6752
rect 94556 6740 94562 6792
rect 96154 6740 96160 6792
rect 96212 6740 96218 6792
rect 96893 6783 96951 6789
rect 96893 6749 96905 6783
rect 96939 6780 96951 6783
rect 96939 6752 97304 6780
rect 96939 6749 96951 6752
rect 96893 6743 96951 6749
rect 46716 6684 60734 6712
rect 46716 6672 46722 6684
rect 83182 6672 83188 6724
rect 83240 6712 83246 6724
rect 93762 6712 93768 6724
rect 83240 6684 93768 6712
rect 83240 6672 83246 6684
rect 93762 6672 93768 6684
rect 93820 6672 93826 6724
rect 94682 6672 94688 6724
rect 94740 6712 94746 6724
rect 97276 6712 97304 6752
rect 97350 6740 97356 6792
rect 97408 6780 97414 6792
rect 97445 6783 97503 6789
rect 97445 6780 97457 6783
rect 97408 6752 97457 6780
rect 97408 6740 97414 6752
rect 97445 6749 97457 6752
rect 97491 6780 97503 6783
rect 98270 6780 98276 6792
rect 97491 6752 98276 6780
rect 97491 6749 97503 6752
rect 97445 6743 97503 6749
rect 98270 6740 98276 6752
rect 98328 6740 98334 6792
rect 98454 6740 98460 6792
rect 98512 6740 98518 6792
rect 98932 6780 98960 6820
rect 99190 6808 99196 6860
rect 99248 6848 99254 6860
rect 100018 6848 100024 6860
rect 99248 6820 100024 6848
rect 99248 6808 99254 6820
rect 100018 6808 100024 6820
rect 100076 6808 100082 6860
rect 100496 6848 100524 6888
rect 106185 6885 106197 6919
rect 106231 6885 106243 6919
rect 106185 6879 106243 6885
rect 100496 6820 102180 6848
rect 99374 6780 99380 6792
rect 98932 6752 99380 6780
rect 99374 6740 99380 6752
rect 99432 6740 99438 6792
rect 99834 6740 99840 6792
rect 99892 6740 99898 6792
rect 100391 6783 100449 6789
rect 100391 6749 100403 6783
rect 100437 6780 100449 6783
rect 100496 6780 100524 6820
rect 100437 6752 100524 6780
rect 101309 6783 101367 6789
rect 100437 6749 100449 6752
rect 100391 6743 100449 6749
rect 101309 6749 101321 6783
rect 101355 6749 101367 6783
rect 101309 6743 101367 6749
rect 98086 6712 98092 6724
rect 94740 6684 97212 6712
rect 97276 6684 98092 6712
rect 94740 6672 94746 6684
rect 20714 6604 20720 6656
rect 20772 6644 20778 6656
rect 45094 6644 45100 6656
rect 20772 6616 45100 6644
rect 20772 6604 20778 6616
rect 45094 6604 45100 6616
rect 45152 6604 45158 6656
rect 82814 6604 82820 6656
rect 82872 6644 82878 6656
rect 94222 6644 94228 6656
rect 82872 6616 94228 6644
rect 82872 6604 82878 6616
rect 94222 6604 94228 6616
rect 94280 6604 94286 6656
rect 95970 6604 95976 6656
rect 96028 6604 96034 6656
rect 96706 6604 96712 6656
rect 96764 6604 96770 6656
rect 97184 6644 97212 6684
rect 98086 6672 98092 6684
rect 98144 6672 98150 6724
rect 101214 6712 101220 6724
rect 101048 6684 101220 6712
rect 97813 6647 97871 6653
rect 97813 6644 97825 6647
rect 97184 6616 97825 6644
rect 97813 6613 97825 6616
rect 97859 6613 97871 6647
rect 97813 6607 97871 6613
rect 98638 6604 98644 6656
rect 98696 6604 98702 6656
rect 99650 6604 99656 6656
rect 99708 6604 99714 6656
rect 99834 6604 99840 6656
rect 99892 6644 99898 6656
rect 101048 6644 101076 6684
rect 101214 6672 101220 6684
rect 101272 6672 101278 6724
rect 101324 6712 101352 6743
rect 101674 6740 101680 6792
rect 101732 6780 101738 6792
rect 102045 6783 102103 6789
rect 102045 6780 102057 6783
rect 101732 6752 102057 6780
rect 101732 6740 101738 6752
rect 102045 6749 102057 6752
rect 102091 6749 102103 6783
rect 102152 6780 102180 6820
rect 102226 6808 102232 6860
rect 102284 6848 102290 6860
rect 106200 6848 106228 6879
rect 107194 6876 107200 6928
rect 107252 6916 107258 6928
rect 110601 6919 110659 6925
rect 107252 6888 108344 6916
rect 107252 6876 107258 6888
rect 102284 6820 106228 6848
rect 102284 6808 102290 6820
rect 106274 6808 106280 6860
rect 106332 6848 106338 6860
rect 108316 6848 108344 6888
rect 110601 6885 110613 6919
rect 110647 6916 110659 6919
rect 110966 6916 110972 6928
rect 110647 6888 110972 6916
rect 110647 6885 110659 6888
rect 110601 6879 110659 6885
rect 110966 6876 110972 6888
rect 111024 6876 111030 6928
rect 112165 6919 112223 6925
rect 112165 6885 112177 6919
rect 112211 6885 112223 6919
rect 112165 6879 112223 6885
rect 109681 6851 109739 6857
rect 109681 6848 109693 6851
rect 106332 6820 108252 6848
rect 108316 6820 109693 6848
rect 106332 6808 106338 6820
rect 102152 6752 102456 6780
rect 102045 6743 102103 6749
rect 102318 6712 102324 6724
rect 101324 6684 102324 6712
rect 102318 6672 102324 6684
rect 102376 6672 102382 6724
rect 102428 6712 102456 6752
rect 102686 6740 102692 6792
rect 102744 6740 102750 6792
rect 106182 6740 106188 6792
rect 106240 6780 106246 6792
rect 106369 6783 106427 6789
rect 106369 6780 106381 6783
rect 106240 6752 106381 6780
rect 106240 6740 106246 6752
rect 106369 6749 106381 6752
rect 106415 6749 106427 6783
rect 106369 6743 106427 6749
rect 107473 6783 107531 6789
rect 107473 6749 107485 6783
rect 107519 6780 107531 6783
rect 107562 6780 107568 6792
rect 107519 6752 107568 6780
rect 107519 6749 107531 6752
rect 107473 6743 107531 6749
rect 107562 6740 107568 6752
rect 107620 6740 107626 6792
rect 108117 6783 108175 6789
rect 108117 6749 108129 6783
rect 108163 6749 108175 6783
rect 108117 6743 108175 6749
rect 107010 6712 107016 6724
rect 102428 6684 107016 6712
rect 107010 6672 107016 6684
rect 107068 6672 107074 6724
rect 108132 6712 108160 6743
rect 107488 6684 108160 6712
rect 108224 6712 108252 6820
rect 109681 6817 109693 6820
rect 109727 6817 109739 6851
rect 109681 6811 109739 6817
rect 110138 6808 110144 6860
rect 110196 6848 110202 6860
rect 112180 6848 112208 6879
rect 110196 6820 112208 6848
rect 112272 6848 112300 6956
rect 114572 6956 118556 6984
rect 112530 6876 112536 6928
rect 112588 6916 112594 6928
rect 113542 6916 113548 6928
rect 112588 6888 113548 6916
rect 112588 6876 112594 6888
rect 113542 6876 113548 6888
rect 113600 6876 113606 6928
rect 114572 6916 114600 6956
rect 113652 6888 113864 6916
rect 113652 6848 113680 6888
rect 112272 6820 113680 6848
rect 110196 6808 110202 6820
rect 113726 6808 113732 6860
rect 113784 6808 113790 6860
rect 113836 6848 113864 6888
rect 114480 6888 114600 6916
rect 114480 6848 114508 6888
rect 114646 6876 114652 6928
rect 114704 6916 114710 6928
rect 116578 6916 116584 6928
rect 114704 6888 116584 6916
rect 114704 6876 114710 6888
rect 116578 6876 116584 6888
rect 116636 6876 116642 6928
rect 116673 6919 116731 6925
rect 116673 6885 116685 6919
rect 116719 6916 116731 6919
rect 116854 6916 116860 6928
rect 116719 6888 116860 6916
rect 116719 6885 116731 6888
rect 116673 6879 116731 6885
rect 116854 6876 116860 6888
rect 116912 6876 116918 6928
rect 118528 6916 118556 6956
rect 118602 6944 118608 6996
rect 118660 6984 118666 6996
rect 144914 6984 144920 6996
rect 118660 6956 144920 6984
rect 118660 6944 118666 6956
rect 144914 6944 144920 6956
rect 144972 6944 144978 6996
rect 150894 6944 150900 6996
rect 150952 6984 150958 6996
rect 151081 6987 151139 6993
rect 151081 6984 151093 6987
rect 150952 6956 151093 6984
rect 150952 6944 150958 6956
rect 151081 6953 151093 6956
rect 151127 6953 151139 6987
rect 151081 6947 151139 6953
rect 151538 6944 151544 6996
rect 151596 6984 151602 6996
rect 151817 6987 151875 6993
rect 151817 6984 151829 6987
rect 151596 6956 151829 6984
rect 151596 6944 151602 6956
rect 151817 6953 151829 6956
rect 151863 6984 151875 6987
rect 152090 6984 152096 6996
rect 151863 6956 152096 6984
rect 151863 6953 151875 6956
rect 151817 6947 151875 6953
rect 152090 6944 152096 6956
rect 152148 6944 152154 6996
rect 153381 6987 153439 6993
rect 153381 6984 153393 6987
rect 153304 6956 153393 6984
rect 118528 6888 118648 6916
rect 113836 6820 114508 6848
rect 114554 6808 114560 6860
rect 114612 6808 114618 6860
rect 116305 6851 116363 6857
rect 116305 6817 116317 6851
rect 116351 6848 116363 6851
rect 118142 6848 118148 6860
rect 116351 6820 118148 6848
rect 116351 6817 116363 6820
rect 116305 6811 116363 6817
rect 118142 6808 118148 6820
rect 118200 6808 118206 6860
rect 118620 6848 118648 6888
rect 145006 6876 145012 6928
rect 145064 6916 145070 6928
rect 148962 6916 148968 6928
rect 145064 6888 148968 6916
rect 145064 6876 145070 6888
rect 148962 6876 148968 6888
rect 149020 6876 149026 6928
rect 150434 6876 150440 6928
rect 150492 6916 150498 6928
rect 150492 6888 152872 6916
rect 150492 6876 150498 6888
rect 133230 6848 133236 6860
rect 118620 6820 133236 6848
rect 133230 6808 133236 6820
rect 133288 6808 133294 6860
rect 151078 6808 151084 6860
rect 151136 6848 151142 6860
rect 151814 6848 151820 6860
rect 151136 6820 151820 6848
rect 151136 6808 151142 6820
rect 151814 6808 151820 6820
rect 151872 6848 151878 6860
rect 152274 6848 152280 6860
rect 151872 6820 152280 6848
rect 151872 6808 151878 6820
rect 152274 6808 152280 6820
rect 152332 6808 152338 6860
rect 108574 6740 108580 6792
rect 108632 6740 108638 6792
rect 108666 6740 108672 6792
rect 108724 6740 108730 6792
rect 109954 6740 109960 6792
rect 110012 6780 110018 6792
rect 110233 6783 110291 6789
rect 110233 6780 110245 6783
rect 110012 6752 110245 6780
rect 110012 6740 110018 6752
rect 110233 6749 110245 6752
rect 110279 6749 110291 6783
rect 110233 6743 110291 6749
rect 110414 6740 110420 6792
rect 110472 6740 110478 6792
rect 110966 6740 110972 6792
rect 111024 6780 111030 6792
rect 111245 6783 111303 6789
rect 111245 6780 111257 6783
rect 111024 6752 111257 6780
rect 111024 6740 111030 6752
rect 111245 6749 111257 6752
rect 111291 6749 111303 6783
rect 111245 6743 111303 6749
rect 112346 6740 112352 6792
rect 112404 6740 112410 6792
rect 112990 6740 112996 6792
rect 113048 6740 113054 6792
rect 115658 6740 115664 6792
rect 115716 6780 115722 6792
rect 116029 6783 116087 6789
rect 116029 6780 116041 6783
rect 115716 6752 116041 6780
rect 115716 6740 115722 6752
rect 116029 6749 116041 6752
rect 116075 6780 116087 6783
rect 116210 6780 116216 6792
rect 116075 6752 116216 6780
rect 116075 6749 116087 6752
rect 116029 6743 116087 6749
rect 116210 6740 116216 6752
rect 116268 6740 116274 6792
rect 118418 6780 118424 6792
rect 116412 6752 118424 6780
rect 109402 6712 109408 6724
rect 108224 6684 109408 6712
rect 107488 6656 107516 6684
rect 109402 6672 109408 6684
rect 109460 6672 109466 6724
rect 109497 6715 109555 6721
rect 109497 6681 109509 6715
rect 109543 6712 109555 6715
rect 113082 6712 113088 6724
rect 109543 6684 113088 6712
rect 109543 6681 109555 6684
rect 109497 6675 109555 6681
rect 113082 6672 113088 6684
rect 113140 6672 113146 6724
rect 113910 6672 113916 6724
rect 113968 6672 113974 6724
rect 99892 6616 101076 6644
rect 99892 6604 99898 6616
rect 101122 6604 101128 6656
rect 101180 6604 101186 6656
rect 101582 6604 101588 6656
rect 101640 6644 101646 6656
rect 101861 6647 101919 6653
rect 101861 6644 101873 6647
rect 101640 6616 101873 6644
rect 101640 6604 101646 6616
rect 101861 6613 101873 6616
rect 101907 6613 101919 6647
rect 101861 6607 101919 6613
rect 102134 6604 102140 6656
rect 102192 6644 102198 6656
rect 102505 6647 102563 6653
rect 102505 6644 102517 6647
rect 102192 6616 102517 6644
rect 102192 6604 102198 6616
rect 102505 6613 102517 6616
rect 102551 6613 102563 6647
rect 102505 6607 102563 6613
rect 103330 6604 103336 6656
rect 103388 6644 103394 6656
rect 107289 6647 107347 6653
rect 107289 6644 107301 6647
rect 103388 6616 107301 6644
rect 103388 6604 103394 6616
rect 107289 6613 107301 6616
rect 107335 6613 107347 6647
rect 107289 6607 107347 6613
rect 107470 6604 107476 6656
rect 107528 6604 107534 6656
rect 107930 6604 107936 6656
rect 107988 6604 107994 6656
rect 108022 6604 108028 6656
rect 108080 6644 108086 6656
rect 109954 6644 109960 6656
rect 108080 6616 109960 6644
rect 108080 6604 108086 6616
rect 109954 6604 109960 6616
rect 110012 6604 110018 6656
rect 110966 6604 110972 6656
rect 111024 6644 111030 6656
rect 111061 6647 111119 6653
rect 111061 6644 111073 6647
rect 111024 6616 111073 6644
rect 111024 6604 111030 6616
rect 111061 6613 111073 6616
rect 111107 6613 111119 6647
rect 111061 6607 111119 6613
rect 111334 6604 111340 6656
rect 111392 6644 111398 6656
rect 112530 6644 112536 6656
rect 111392 6616 112536 6644
rect 111392 6604 111398 6616
rect 112530 6604 112536 6616
rect 112588 6604 112594 6656
rect 112806 6604 112812 6656
rect 112864 6604 112870 6656
rect 115106 6604 115112 6656
rect 115164 6644 115170 6656
rect 115382 6644 115388 6656
rect 115164 6616 115388 6644
rect 115164 6604 115170 6616
rect 115382 6604 115388 6616
rect 115440 6644 115446 6656
rect 116412 6653 116440 6752
rect 118418 6740 118424 6752
rect 118476 6740 118482 6792
rect 150618 6740 150624 6792
rect 150676 6780 150682 6792
rect 150989 6783 151047 6789
rect 150989 6780 151001 6783
rect 150676 6752 151001 6780
rect 150676 6740 150682 6752
rect 150989 6749 151001 6752
rect 151035 6749 151047 6783
rect 150989 6743 151047 6749
rect 151357 6783 151415 6789
rect 151357 6749 151369 6783
rect 151403 6780 151415 6783
rect 151538 6780 151544 6792
rect 151403 6752 151544 6780
rect 151403 6749 151415 6752
rect 151357 6743 151415 6749
rect 151538 6740 151544 6752
rect 151596 6740 151602 6792
rect 152090 6740 152096 6792
rect 152148 6780 152154 6792
rect 152185 6783 152243 6789
rect 152185 6780 152197 6783
rect 152148 6752 152197 6780
rect 152148 6740 152154 6752
rect 152185 6749 152197 6752
rect 152231 6780 152243 6783
rect 152844 6780 152872 6888
rect 153304 6848 153332 6956
rect 153381 6953 153393 6956
rect 153427 6953 153439 6987
rect 153381 6947 153439 6953
rect 180766 6956 190454 6984
rect 161290 6916 161296 6928
rect 154592 6888 161296 6916
rect 153378 6848 153384 6860
rect 153304 6820 153384 6848
rect 153378 6808 153384 6820
rect 153436 6808 153442 6860
rect 153838 6808 153844 6860
rect 153896 6848 153902 6860
rect 154592 6848 154620 6888
rect 161290 6876 161296 6888
rect 161348 6876 161354 6928
rect 161382 6876 161388 6928
rect 161440 6916 161446 6928
rect 180766 6916 180794 6956
rect 161440 6888 180794 6916
rect 161440 6876 161446 6888
rect 190178 6876 190184 6928
rect 190236 6876 190242 6928
rect 190426 6916 190454 6956
rect 213914 6944 213920 6996
rect 213972 6984 213978 6996
rect 220814 6984 220820 6996
rect 213972 6956 220820 6984
rect 213972 6944 213978 6956
rect 220814 6944 220820 6956
rect 220872 6944 220878 6996
rect 221274 6944 221280 6996
rect 221332 6984 221338 6996
rect 229738 6984 229744 6996
rect 221332 6956 229744 6984
rect 221332 6944 221338 6956
rect 229738 6944 229744 6956
rect 229796 6944 229802 6996
rect 249978 6944 249984 6996
rect 250036 6984 250042 6996
rect 259730 6984 259736 6996
rect 250036 6956 259736 6984
rect 250036 6944 250042 6956
rect 259730 6944 259736 6956
rect 259788 6944 259794 6996
rect 261570 6944 261576 6996
rect 261628 6984 261634 6996
rect 261628 6956 263594 6984
rect 261628 6944 261634 6956
rect 210418 6916 210424 6928
rect 190426 6888 210424 6916
rect 210418 6876 210424 6888
rect 210476 6876 210482 6928
rect 210510 6876 210516 6928
rect 210568 6916 210574 6928
rect 223485 6919 223543 6925
rect 210568 6888 219296 6916
rect 210568 6876 210574 6888
rect 153896 6820 154620 6848
rect 153896 6808 153902 6820
rect 155034 6808 155040 6860
rect 155092 6848 155098 6860
rect 157242 6848 157248 6860
rect 155092 6820 157248 6848
rect 155092 6808 155098 6820
rect 157242 6808 157248 6820
rect 157300 6808 157306 6860
rect 188816 6820 216076 6848
rect 188816 6792 188844 6820
rect 153565 6783 153623 6789
rect 152231 6752 152780 6780
rect 152844 6776 153332 6780
rect 153565 6776 153577 6783
rect 152844 6752 153577 6776
rect 152231 6749 152243 6752
rect 152185 6743 152243 6749
rect 116514 6715 116572 6721
rect 116514 6681 116526 6715
rect 116560 6712 116572 6715
rect 116854 6712 116860 6724
rect 116560 6684 116860 6712
rect 116560 6681 116572 6684
rect 116514 6675 116572 6681
rect 116854 6672 116860 6684
rect 116912 6672 116918 6724
rect 117409 6715 117467 6721
rect 117409 6681 117421 6715
rect 117455 6712 117467 6715
rect 117774 6712 117780 6724
rect 117455 6684 117780 6712
rect 117455 6681 117467 6684
rect 117409 6675 117467 6681
rect 117774 6672 117780 6684
rect 117832 6672 117838 6724
rect 118142 6672 118148 6724
rect 118200 6712 118206 6724
rect 118329 6715 118387 6721
rect 118329 6712 118341 6715
rect 118200 6684 118341 6712
rect 118200 6672 118206 6684
rect 118329 6681 118341 6684
rect 118375 6681 118387 6715
rect 118329 6675 118387 6681
rect 142798 6672 142804 6724
rect 142856 6712 142862 6724
rect 152458 6712 152464 6724
rect 142856 6684 152464 6712
rect 142856 6672 142862 6684
rect 152458 6672 152464 6684
rect 152516 6672 152522 6724
rect 152752 6712 152780 6752
rect 153304 6749 153577 6752
rect 153611 6749 153623 6783
rect 153304 6748 153623 6749
rect 153565 6743 153623 6748
rect 153746 6740 153752 6792
rect 153804 6780 153810 6792
rect 188798 6780 188804 6792
rect 153804 6752 188804 6780
rect 153804 6740 153810 6752
rect 188798 6740 188804 6752
rect 188856 6740 188862 6792
rect 189718 6740 189724 6792
rect 189776 6780 189782 6792
rect 190365 6783 190423 6789
rect 190365 6780 190377 6783
rect 189776 6752 190377 6780
rect 189776 6740 189782 6752
rect 190365 6749 190377 6752
rect 190411 6749 190423 6783
rect 190365 6743 190423 6749
rect 213178 6740 213184 6792
rect 213236 6740 213242 6792
rect 213546 6740 213552 6792
rect 213604 6780 213610 6792
rect 213604 6752 215294 6780
rect 213604 6740 213610 6752
rect 152752 6684 153424 6712
rect 116397 6647 116455 6653
rect 116397 6644 116409 6647
rect 115440 6616 116409 6644
rect 115440 6604 115446 6616
rect 116397 6613 116409 6616
rect 116443 6613 116455 6647
rect 116397 6607 116455 6613
rect 116670 6604 116676 6656
rect 116728 6644 116734 6656
rect 117501 6647 117559 6653
rect 117501 6644 117513 6647
rect 116728 6616 117513 6644
rect 116728 6604 116734 6616
rect 117501 6613 117513 6616
rect 117547 6613 117559 6647
rect 117501 6607 117559 6613
rect 117590 6604 117596 6656
rect 117648 6644 117654 6656
rect 118050 6644 118056 6656
rect 117648 6616 118056 6644
rect 117648 6604 117654 6616
rect 118050 6604 118056 6616
rect 118108 6644 118114 6656
rect 118421 6647 118479 6653
rect 118421 6644 118433 6647
rect 118108 6616 118433 6644
rect 118108 6604 118114 6616
rect 118421 6613 118433 6616
rect 118467 6613 118479 6647
rect 118421 6607 118479 6613
rect 119982 6604 119988 6656
rect 120040 6644 120046 6656
rect 128078 6644 128084 6656
rect 120040 6616 128084 6644
rect 120040 6604 120046 6616
rect 128078 6604 128084 6616
rect 128136 6644 128142 6656
rect 140314 6644 140320 6656
rect 128136 6616 140320 6644
rect 128136 6604 128142 6616
rect 140314 6604 140320 6616
rect 140372 6604 140378 6656
rect 148962 6604 148968 6656
rect 149020 6644 149026 6656
rect 151446 6644 151452 6656
rect 149020 6616 151452 6644
rect 149020 6604 149026 6616
rect 151446 6604 151452 6616
rect 151504 6604 151510 6656
rect 151541 6647 151599 6653
rect 151541 6613 151553 6647
rect 151587 6644 151599 6647
rect 151722 6644 151728 6656
rect 151587 6616 151728 6644
rect 151587 6613 151599 6616
rect 151541 6607 151599 6613
rect 151722 6604 151728 6616
rect 151780 6604 151786 6656
rect 153396 6644 153424 6684
rect 153838 6672 153844 6724
rect 153896 6712 153902 6724
rect 189350 6712 189356 6724
rect 153896 6684 189356 6712
rect 153896 6672 153902 6684
rect 189350 6672 189356 6684
rect 189408 6712 189414 6724
rect 189810 6712 189816 6724
rect 189408 6684 189816 6712
rect 189408 6672 189414 6684
rect 189810 6672 189816 6684
rect 189868 6672 189874 6724
rect 213638 6712 213644 6724
rect 195946 6684 213644 6712
rect 167730 6644 167736 6656
rect 153396 6616 167736 6644
rect 167730 6604 167736 6616
rect 167788 6604 167794 6656
rect 168834 6604 168840 6656
rect 168892 6644 168898 6656
rect 195946 6644 195974 6684
rect 213638 6672 213644 6684
rect 213696 6712 213702 6724
rect 213825 6715 213883 6721
rect 213825 6712 213837 6715
rect 213696 6684 213837 6712
rect 213696 6672 213702 6684
rect 213825 6681 213837 6684
rect 213871 6681 213883 6715
rect 213825 6675 213883 6681
rect 168892 6616 195974 6644
rect 168892 6604 168898 6616
rect 210326 6604 210332 6656
rect 210384 6644 210390 6656
rect 213914 6644 213920 6656
rect 210384 6616 213920 6644
rect 210384 6604 210390 6616
rect 213914 6604 213920 6616
rect 213972 6604 213978 6656
rect 215266 6644 215294 6752
rect 216048 6721 216076 6820
rect 216858 6808 216864 6860
rect 216916 6808 216922 6860
rect 217244 6820 217456 6848
rect 216122 6740 216128 6792
rect 216180 6780 216186 6792
rect 216585 6783 216643 6789
rect 216585 6780 216597 6783
rect 216180 6752 216597 6780
rect 216180 6740 216186 6752
rect 216585 6749 216597 6752
rect 216631 6780 216643 6783
rect 217244 6780 217272 6820
rect 216631 6752 217272 6780
rect 216631 6749 216643 6752
rect 216585 6743 216643 6749
rect 217318 6740 217324 6792
rect 217376 6740 217382 6792
rect 217428 6780 217456 6820
rect 217870 6808 217876 6860
rect 217928 6848 217934 6860
rect 218238 6848 218244 6860
rect 217928 6820 218244 6848
rect 217928 6808 217934 6820
rect 218238 6808 218244 6820
rect 218296 6808 218302 6860
rect 219268 6848 219296 6888
rect 223485 6885 223497 6919
rect 223531 6885 223543 6919
rect 223485 6879 223543 6885
rect 219618 6848 219624 6860
rect 219268 6820 219624 6848
rect 219618 6808 219624 6820
rect 219676 6808 219682 6860
rect 223500 6848 223528 6879
rect 224862 6876 224868 6928
rect 224920 6916 224926 6928
rect 227622 6916 227628 6928
rect 224920 6888 227628 6916
rect 224920 6876 224926 6888
rect 227622 6876 227628 6888
rect 227680 6876 227686 6928
rect 236454 6876 236460 6928
rect 236512 6916 236518 6928
rect 261757 6919 261815 6925
rect 236512 6888 241514 6916
rect 236512 6876 236518 6888
rect 224310 6848 224316 6860
rect 223500 6820 224316 6848
rect 224310 6808 224316 6820
rect 224368 6848 224374 6860
rect 226610 6848 226616 6860
rect 224368 6820 226616 6848
rect 224368 6808 224374 6820
rect 226610 6808 226616 6820
rect 226668 6808 226674 6860
rect 226978 6808 226984 6860
rect 227036 6808 227042 6860
rect 241238 6848 241244 6860
rect 231826 6820 241244 6848
rect 219158 6780 219164 6792
rect 217428 6752 219164 6780
rect 219158 6740 219164 6752
rect 219216 6780 219222 6792
rect 223301 6783 223359 6789
rect 223301 6780 223313 6783
rect 219216 6752 223313 6780
rect 219216 6740 219222 6752
rect 223301 6749 223313 6752
rect 223347 6780 223359 6783
rect 224218 6780 224224 6792
rect 223347 6752 224224 6780
rect 223347 6749 223359 6752
rect 223301 6743 223359 6749
rect 224218 6740 224224 6752
rect 224276 6780 224282 6792
rect 224770 6780 224776 6792
rect 224276 6752 224776 6780
rect 224276 6740 224282 6752
rect 224770 6740 224776 6752
rect 224828 6740 224834 6792
rect 224954 6740 224960 6792
rect 225012 6780 225018 6792
rect 225601 6783 225659 6789
rect 225601 6780 225613 6783
rect 225012 6752 225613 6780
rect 225012 6740 225018 6752
rect 225601 6749 225613 6752
rect 225647 6749 225659 6783
rect 225601 6743 225659 6749
rect 226705 6783 226763 6789
rect 226705 6749 226717 6783
rect 226751 6780 226763 6783
rect 231826 6780 231854 6820
rect 241238 6808 241244 6820
rect 241296 6808 241302 6860
rect 241486 6848 241514 6888
rect 261757 6885 261769 6919
rect 261803 6885 261815 6919
rect 263566 6916 263594 6956
rect 264606 6944 264612 6996
rect 264664 6984 264670 6996
rect 267642 6984 267648 6996
rect 264664 6956 267648 6984
rect 264664 6944 264670 6956
rect 267642 6944 267648 6956
rect 267700 6944 267706 6996
rect 267734 6944 267740 6996
rect 267792 6984 267798 6996
rect 269209 6987 269267 6993
rect 269209 6984 269221 6987
rect 267792 6956 269221 6984
rect 267792 6944 267798 6956
rect 269209 6953 269221 6956
rect 269255 6953 269267 6987
rect 269209 6947 269267 6953
rect 270494 6944 270500 6996
rect 270552 6944 270558 6996
rect 268286 6916 268292 6928
rect 263566 6888 268292 6916
rect 261757 6879 261815 6885
rect 250070 6848 250076 6860
rect 241486 6820 250076 6848
rect 250070 6808 250076 6820
rect 250128 6808 250134 6860
rect 251634 6808 251640 6860
rect 251692 6848 251698 6860
rect 261772 6848 261800 6879
rect 268286 6876 268292 6888
rect 268344 6876 268350 6928
rect 270512 6916 270540 6944
rect 268396 6888 270540 6916
rect 263597 6851 263655 6857
rect 263597 6848 263609 6851
rect 251692 6820 261800 6848
rect 262416 6820 263609 6848
rect 251692 6808 251698 6820
rect 226751 6752 231854 6780
rect 238389 6783 238447 6789
rect 226751 6749 226763 6752
rect 226705 6743 226763 6749
rect 238389 6749 238401 6783
rect 238435 6780 238447 6783
rect 238435 6752 239168 6780
rect 238435 6749 238447 6752
rect 238389 6743 238447 6749
rect 216033 6715 216091 6721
rect 216033 6681 216045 6715
rect 216079 6712 216091 6715
rect 216306 6712 216312 6724
rect 216079 6684 216312 6712
rect 216079 6681 216091 6684
rect 216033 6675 216091 6681
rect 216306 6672 216312 6684
rect 216364 6672 216370 6724
rect 219250 6712 219256 6724
rect 216416 6684 219256 6712
rect 216416 6644 216444 6684
rect 219250 6672 219256 6684
rect 219308 6672 219314 6724
rect 224126 6712 224132 6724
rect 219360 6684 224132 6712
rect 215266 6616 216444 6644
rect 216490 6604 216496 6656
rect 216548 6604 216554 6656
rect 216677 6647 216735 6653
rect 216677 6613 216689 6647
rect 216723 6644 216735 6647
rect 217042 6644 217048 6656
rect 216723 6616 217048 6644
rect 216723 6613 216735 6616
rect 216677 6607 216735 6613
rect 217042 6604 217048 6616
rect 217100 6644 217106 6656
rect 217413 6647 217471 6653
rect 217413 6644 217425 6647
rect 217100 6616 217425 6644
rect 217100 6604 217106 6616
rect 217413 6613 217425 6616
rect 217459 6613 217471 6647
rect 217413 6607 217471 6613
rect 218698 6604 218704 6656
rect 218756 6644 218762 6656
rect 219360 6644 219388 6684
rect 224126 6672 224132 6684
rect 224184 6712 224190 6724
rect 224184 6684 224954 6712
rect 224184 6672 224190 6684
rect 218756 6616 219388 6644
rect 218756 6604 218762 6616
rect 219526 6604 219532 6656
rect 219584 6644 219590 6656
rect 221090 6644 221096 6656
rect 219584 6616 221096 6644
rect 219584 6604 219590 6616
rect 221090 6604 221096 6616
rect 221148 6604 221154 6656
rect 223482 6604 223488 6656
rect 223540 6644 223546 6656
rect 224221 6647 224279 6653
rect 224221 6644 224233 6647
rect 223540 6616 224233 6644
rect 223540 6604 223546 6616
rect 224221 6613 224233 6616
rect 224267 6613 224279 6647
rect 224926 6644 224954 6684
rect 225782 6672 225788 6724
rect 225840 6712 225846 6724
rect 233050 6712 233056 6724
rect 225840 6684 233056 6712
rect 225840 6672 225846 6684
rect 233050 6672 233056 6684
rect 233108 6672 233114 6724
rect 239030 6672 239036 6724
rect 239088 6672 239094 6724
rect 239140 6712 239168 6752
rect 241330 6740 241336 6792
rect 241388 6780 241394 6792
rect 248414 6780 248420 6792
rect 241388 6752 248420 6780
rect 241388 6740 241394 6752
rect 248414 6740 248420 6752
rect 248472 6740 248478 6792
rect 248506 6740 248512 6792
rect 248564 6780 248570 6792
rect 248693 6783 248751 6789
rect 248693 6780 248705 6783
rect 248564 6752 248705 6780
rect 248564 6740 248570 6752
rect 248693 6749 248705 6752
rect 248739 6749 248751 6783
rect 248693 6743 248751 6749
rect 249334 6740 249340 6792
rect 249392 6740 249398 6792
rect 251358 6740 251364 6792
rect 251416 6740 251422 6792
rect 251450 6740 251456 6792
rect 251508 6740 251514 6792
rect 253014 6740 253020 6792
rect 253072 6740 253078 6792
rect 253198 6740 253204 6792
rect 253256 6780 253262 6792
rect 253293 6783 253351 6789
rect 253293 6780 253305 6783
rect 253256 6752 253305 6780
rect 253256 6740 253262 6752
rect 253293 6749 253305 6752
rect 253339 6749 253351 6783
rect 253293 6743 253351 6749
rect 256605 6783 256663 6789
rect 256605 6749 256617 6783
rect 256651 6780 256663 6783
rect 256694 6780 256700 6792
rect 256651 6752 256700 6780
rect 256651 6749 256663 6752
rect 256605 6743 256663 6749
rect 256694 6740 256700 6752
rect 256752 6740 256758 6792
rect 261021 6783 261079 6789
rect 261021 6749 261033 6783
rect 261067 6780 261079 6783
rect 261938 6780 261944 6792
rect 261067 6752 261944 6780
rect 261067 6749 261079 6752
rect 261021 6743 261079 6749
rect 261938 6740 261944 6752
rect 261996 6740 262002 6792
rect 262416 6789 262444 6820
rect 263597 6817 263609 6820
rect 263643 6848 263655 6851
rect 263962 6848 263968 6860
rect 263643 6820 263968 6848
rect 263643 6817 263655 6820
rect 263597 6811 263655 6817
rect 263962 6808 263968 6820
rect 264020 6808 264026 6860
rect 264054 6808 264060 6860
rect 264112 6848 264118 6860
rect 267918 6848 267924 6860
rect 264112 6820 267924 6848
rect 264112 6808 264118 6820
rect 267918 6808 267924 6820
rect 267976 6808 267982 6860
rect 262401 6783 262459 6789
rect 262401 6749 262413 6783
rect 262447 6749 262459 6783
rect 262401 6743 262459 6749
rect 262769 6783 262827 6789
rect 262769 6749 262781 6783
rect 262815 6780 262827 6783
rect 263226 6780 263232 6792
rect 262815 6752 263232 6780
rect 262815 6749 262827 6752
rect 262769 6743 262827 6749
rect 263226 6740 263232 6752
rect 263284 6740 263290 6792
rect 263686 6740 263692 6792
rect 263744 6740 263750 6792
rect 264425 6783 264483 6789
rect 264425 6749 264437 6783
rect 264471 6780 264483 6783
rect 264471 6752 265848 6780
rect 264471 6749 264483 6752
rect 264425 6743 264483 6749
rect 253106 6712 253112 6724
rect 239140 6684 241514 6712
rect 225693 6647 225751 6653
rect 225693 6644 225705 6647
rect 224926 6616 225705 6644
rect 224221 6607 224279 6613
rect 225693 6613 225705 6616
rect 225739 6613 225751 6647
rect 225693 6607 225751 6613
rect 226150 6604 226156 6656
rect 226208 6644 226214 6656
rect 226794 6644 226800 6656
rect 226208 6616 226800 6644
rect 226208 6604 226214 6616
rect 226794 6604 226800 6616
rect 226852 6604 226858 6656
rect 241486 6644 241514 6684
rect 244246 6684 253112 6712
rect 244246 6644 244274 6684
rect 253106 6672 253112 6684
rect 253164 6672 253170 6724
rect 255685 6715 255743 6721
rect 255685 6712 255697 6715
rect 253216 6684 255697 6712
rect 241486 6616 244274 6644
rect 248509 6647 248567 6653
rect 248509 6613 248521 6647
rect 248555 6644 248567 6647
rect 248874 6644 248880 6656
rect 248555 6616 248880 6644
rect 248555 6613 248567 6616
rect 248509 6607 248567 6613
rect 248874 6604 248880 6616
rect 248932 6604 248938 6656
rect 249153 6647 249211 6653
rect 249153 6613 249165 6647
rect 249199 6644 249211 6647
rect 249242 6644 249248 6656
rect 249199 6616 249248 6644
rect 249199 6613 249211 6616
rect 249153 6607 249211 6613
rect 249242 6604 249248 6616
rect 249300 6604 249306 6656
rect 251634 6604 251640 6656
rect 251692 6604 251698 6656
rect 251726 6604 251732 6656
rect 251784 6644 251790 6656
rect 253216 6644 253244 6684
rect 255685 6681 255697 6684
rect 255731 6712 255743 6715
rect 260834 6712 260840 6724
rect 255731 6684 260840 6712
rect 255731 6681 255743 6684
rect 255685 6675 255743 6681
rect 260834 6672 260840 6684
rect 260892 6672 260898 6724
rect 262232 6684 264836 6712
rect 251784 6616 253244 6644
rect 251784 6604 251790 6616
rect 253842 6604 253848 6656
rect 253900 6644 253906 6656
rect 255590 6644 255596 6656
rect 253900 6616 255596 6644
rect 253900 6604 253906 6616
rect 255590 6604 255596 6616
rect 255648 6604 255654 6656
rect 255774 6604 255780 6656
rect 255832 6604 255838 6656
rect 256421 6647 256479 6653
rect 256421 6613 256433 6647
rect 256467 6644 256479 6647
rect 256602 6644 256608 6656
rect 256467 6616 256608 6644
rect 256467 6613 256479 6616
rect 256421 6607 256479 6613
rect 256602 6604 256608 6616
rect 256660 6604 256666 6656
rect 262232 6653 262260 6684
rect 262217 6647 262275 6653
rect 262217 6613 262229 6647
rect 262263 6613 262275 6647
rect 262217 6607 262275 6613
rect 263042 6604 263048 6656
rect 263100 6604 263106 6656
rect 263778 6604 263784 6656
rect 263836 6604 263842 6656
rect 264808 6644 264836 6684
rect 264882 6672 264888 6724
rect 264940 6672 264946 6724
rect 265820 6712 265848 6752
rect 265894 6740 265900 6792
rect 265952 6740 265958 6792
rect 266814 6740 266820 6792
rect 266872 6740 266878 6792
rect 266909 6783 266967 6789
rect 266909 6749 266921 6783
rect 266955 6780 266967 6783
rect 267274 6780 267280 6792
rect 266955 6752 267280 6780
rect 266955 6749 266967 6752
rect 266909 6743 266967 6749
rect 267274 6740 267280 6752
rect 267332 6740 267338 6792
rect 267550 6740 267556 6792
rect 267608 6780 267614 6792
rect 267608 6752 267872 6780
rect 267608 6740 267614 6752
rect 267734 6712 267740 6724
rect 265820 6684 267740 6712
rect 267734 6672 267740 6684
rect 267792 6672 267798 6724
rect 267844 6712 267872 6752
rect 268010 6740 268016 6792
rect 268068 6740 268074 6792
rect 268396 6712 268424 6888
rect 268565 6851 268623 6857
rect 268565 6817 268577 6851
rect 268611 6848 268623 6851
rect 268746 6848 268752 6860
rect 268611 6820 268752 6848
rect 268611 6817 268623 6820
rect 268565 6811 268623 6817
rect 268746 6808 268752 6820
rect 268804 6808 268810 6860
rect 270218 6808 270224 6860
rect 270276 6848 270282 6860
rect 270497 6851 270555 6857
rect 270497 6848 270509 6851
rect 270276 6820 270509 6848
rect 270276 6808 270282 6820
rect 270497 6817 270509 6820
rect 270543 6817 270555 6851
rect 270497 6811 270555 6817
rect 269206 6740 269212 6792
rect 269264 6740 269270 6792
rect 269850 6740 269856 6792
rect 269908 6740 269914 6792
rect 270034 6740 270040 6792
rect 270092 6740 270098 6792
rect 270589 6783 270647 6789
rect 270589 6749 270601 6783
rect 270635 6749 270647 6783
rect 270589 6743 270647 6749
rect 267844 6684 268424 6712
rect 265986 6644 265992 6656
rect 264808 6616 265992 6644
rect 265986 6604 265992 6616
rect 266044 6604 266050 6656
rect 266081 6647 266139 6653
rect 266081 6613 266093 6647
rect 266127 6644 266139 6647
rect 266354 6644 266360 6656
rect 266127 6616 266360 6644
rect 266127 6613 266139 6616
rect 266081 6607 266139 6613
rect 266354 6604 266360 6616
rect 266412 6604 266418 6656
rect 266630 6604 266636 6656
rect 266688 6644 266694 6656
rect 267093 6647 267151 6653
rect 267093 6644 267105 6647
rect 266688 6616 267105 6644
rect 266688 6604 266694 6616
rect 267093 6613 267105 6616
rect 267139 6613 267151 6647
rect 267093 6607 267151 6613
rect 267642 6604 267648 6656
rect 267700 6644 267706 6656
rect 270126 6644 270132 6656
rect 267700 6616 270132 6644
rect 267700 6604 267706 6616
rect 270126 6604 270132 6616
rect 270184 6644 270190 6656
rect 270604 6644 270632 6743
rect 270184 6616 270632 6644
rect 270184 6604 270190 6616
rect 1104 6554 271651 6576
rect 1104 6502 68546 6554
rect 68598 6502 68610 6554
rect 68662 6502 68674 6554
rect 68726 6502 68738 6554
rect 68790 6502 68802 6554
rect 68854 6502 136143 6554
rect 136195 6502 136207 6554
rect 136259 6502 136271 6554
rect 136323 6502 136335 6554
rect 136387 6502 136399 6554
rect 136451 6502 203740 6554
rect 203792 6502 203804 6554
rect 203856 6502 203868 6554
rect 203920 6502 203932 6554
rect 203984 6502 203996 6554
rect 204048 6502 271337 6554
rect 271389 6502 271401 6554
rect 271453 6502 271465 6554
rect 271517 6502 271529 6554
rect 271581 6502 271593 6554
rect 271645 6502 271651 6554
rect 1104 6480 271651 6502
rect 12894 6400 12900 6452
rect 12952 6440 12958 6452
rect 42702 6440 42708 6452
rect 12952 6412 42708 6440
rect 12952 6400 12958 6412
rect 42702 6400 42708 6412
rect 42760 6400 42766 6452
rect 72326 6400 72332 6452
rect 72384 6440 72390 6452
rect 93946 6440 93952 6452
rect 72384 6412 93952 6440
rect 72384 6400 72390 6412
rect 93946 6400 93952 6412
rect 94004 6400 94010 6452
rect 95326 6400 95332 6452
rect 95384 6440 95390 6452
rect 97718 6440 97724 6452
rect 95384 6412 97724 6440
rect 95384 6400 95390 6412
rect 97718 6400 97724 6412
rect 97776 6400 97782 6452
rect 98362 6400 98368 6452
rect 98420 6400 98426 6452
rect 98730 6400 98736 6452
rect 98788 6400 98794 6452
rect 100021 6443 100079 6449
rect 100021 6440 100033 6443
rect 98840 6412 100033 6440
rect 8478 6332 8484 6384
rect 8536 6372 8542 6384
rect 38746 6372 38752 6384
rect 8536 6344 38752 6372
rect 8536 6332 8542 6344
rect 38746 6332 38752 6344
rect 38804 6332 38810 6384
rect 55766 6372 55772 6384
rect 51368 6344 55772 6372
rect 15562 6264 15568 6316
rect 15620 6304 15626 6316
rect 49510 6304 49516 6316
rect 15620 6276 49516 6304
rect 15620 6264 15626 6276
rect 49510 6264 49516 6276
rect 49568 6264 49574 6316
rect 13630 6196 13636 6248
rect 13688 6236 13694 6248
rect 47486 6236 47492 6248
rect 13688 6208 47492 6236
rect 13688 6196 13694 6208
rect 47486 6196 47492 6208
rect 47544 6196 47550 6248
rect 48866 6236 48872 6248
rect 47596 6208 48872 6236
rect 13722 6128 13728 6180
rect 13780 6168 13786 6180
rect 47596 6168 47624 6208
rect 48866 6196 48872 6208
rect 48924 6196 48930 6248
rect 13780 6140 47624 6168
rect 13780 6128 13786 6140
rect 48038 6128 48044 6180
rect 48096 6168 48102 6180
rect 51368 6168 51396 6344
rect 55766 6332 55772 6344
rect 55824 6332 55830 6384
rect 95513 6375 95571 6381
rect 95513 6341 95525 6375
rect 95559 6372 95571 6375
rect 96706 6372 96712 6384
rect 95559 6344 96712 6372
rect 95559 6341 95571 6344
rect 95513 6335 95571 6341
rect 96706 6332 96712 6344
rect 96764 6332 96770 6384
rect 96798 6332 96804 6384
rect 96856 6372 96862 6384
rect 98380 6372 98408 6400
rect 96856 6344 98408 6372
rect 96856 6332 96862 6344
rect 98546 6332 98552 6384
rect 98604 6372 98610 6384
rect 98840 6372 98868 6412
rect 100021 6409 100033 6412
rect 100067 6409 100079 6443
rect 100021 6403 100079 6409
rect 101030 6400 101036 6452
rect 101088 6440 101094 6452
rect 101858 6440 101864 6452
rect 101088 6412 101864 6440
rect 101088 6400 101094 6412
rect 101858 6400 101864 6412
rect 101916 6400 101922 6452
rect 102318 6400 102324 6452
rect 102376 6400 102382 6452
rect 108022 6440 108028 6452
rect 102428 6412 108028 6440
rect 102428 6372 102456 6412
rect 108022 6400 108028 6412
rect 108080 6400 108086 6452
rect 108117 6443 108175 6449
rect 108117 6409 108129 6443
rect 108163 6440 108175 6443
rect 109310 6440 109316 6452
rect 108163 6412 109316 6440
rect 108163 6409 108175 6412
rect 108117 6403 108175 6409
rect 109310 6400 109316 6412
rect 109368 6400 109374 6452
rect 110414 6440 110420 6452
rect 109696 6412 110420 6440
rect 98604 6344 98868 6372
rect 98932 6344 102456 6372
rect 102873 6375 102931 6381
rect 98604 6332 98610 6344
rect 51442 6264 51448 6316
rect 51500 6304 51506 6316
rect 52362 6304 52368 6316
rect 51500 6276 52368 6304
rect 51500 6264 51506 6276
rect 52362 6264 52368 6276
rect 52420 6264 52426 6316
rect 52917 6307 52975 6313
rect 52917 6273 52929 6307
rect 52963 6273 52975 6307
rect 52917 6267 52975 6273
rect 48096 6140 51396 6168
rect 52932 6168 52960 6267
rect 80238 6264 80244 6316
rect 80296 6304 80302 6316
rect 91925 6307 91983 6313
rect 91925 6304 91937 6307
rect 80296 6276 91937 6304
rect 80296 6264 80302 6276
rect 91925 6273 91937 6276
rect 91971 6273 91983 6307
rect 91925 6267 91983 6273
rect 92934 6264 92940 6316
rect 92992 6264 92998 6316
rect 94869 6307 94927 6313
rect 94869 6273 94881 6307
rect 94915 6304 94927 6307
rect 95234 6304 95240 6316
rect 94915 6276 95240 6304
rect 94915 6273 94927 6276
rect 94869 6267 94927 6273
rect 95234 6264 95240 6276
rect 95292 6264 95298 6316
rect 97902 6264 97908 6316
rect 97960 6264 97966 6316
rect 98270 6264 98276 6316
rect 98328 6304 98334 6316
rect 98365 6307 98423 6313
rect 98365 6304 98377 6307
rect 98328 6276 98377 6304
rect 98328 6264 98334 6276
rect 98365 6273 98377 6276
rect 98411 6304 98423 6307
rect 98932 6304 98960 6344
rect 102873 6341 102885 6375
rect 102919 6372 102931 6375
rect 105998 6372 106004 6384
rect 102919 6344 106004 6372
rect 102919 6341 102931 6344
rect 102873 6335 102931 6341
rect 105998 6332 106004 6344
rect 106056 6332 106062 6384
rect 107105 6375 107163 6381
rect 107105 6341 107117 6375
rect 107151 6372 107163 6375
rect 109696 6372 109724 6412
rect 110414 6400 110420 6412
rect 110472 6400 110478 6452
rect 112809 6443 112867 6449
rect 112809 6409 112821 6443
rect 112855 6440 112867 6443
rect 113910 6440 113916 6452
rect 112855 6412 113916 6440
rect 112855 6409 112867 6412
rect 112809 6403 112867 6409
rect 113910 6400 113916 6412
rect 113968 6400 113974 6452
rect 115198 6400 115204 6452
rect 115256 6440 115262 6452
rect 115474 6440 115480 6452
rect 115256 6412 115480 6440
rect 115256 6400 115262 6412
rect 115474 6400 115480 6412
rect 115532 6440 115538 6452
rect 116854 6440 116860 6452
rect 115532 6412 116860 6440
rect 115532 6400 115538 6412
rect 116854 6400 116860 6412
rect 116912 6400 116918 6452
rect 117866 6400 117872 6452
rect 117924 6440 117930 6452
rect 118050 6440 118056 6452
rect 117924 6412 118056 6440
rect 117924 6400 117930 6412
rect 118050 6400 118056 6412
rect 118108 6400 118114 6452
rect 118142 6400 118148 6452
rect 118200 6400 118206 6452
rect 118234 6400 118240 6452
rect 118292 6440 118298 6452
rect 118973 6443 119031 6449
rect 118973 6440 118985 6443
rect 118292 6412 118985 6440
rect 118292 6400 118298 6412
rect 118973 6409 118985 6412
rect 119019 6409 119031 6443
rect 118973 6403 119031 6409
rect 119157 6443 119215 6449
rect 119157 6409 119169 6443
rect 119203 6440 119215 6443
rect 120074 6440 120080 6452
rect 119203 6412 120080 6440
rect 119203 6409 119215 6412
rect 119157 6403 119215 6409
rect 120074 6400 120080 6412
rect 120132 6400 120138 6452
rect 130378 6400 130384 6452
rect 130436 6440 130442 6452
rect 148134 6440 148140 6452
rect 130436 6412 148140 6440
rect 130436 6400 130442 6412
rect 148134 6400 148140 6412
rect 148192 6400 148198 6452
rect 149054 6400 149060 6452
rect 149112 6440 149118 6452
rect 150250 6440 150256 6452
rect 149112 6412 150256 6440
rect 149112 6400 149118 6412
rect 150250 6400 150256 6412
rect 150308 6440 150314 6452
rect 150986 6440 150992 6452
rect 150308 6412 150992 6440
rect 150308 6400 150314 6412
rect 150986 6400 150992 6412
rect 151044 6400 151050 6452
rect 151262 6400 151268 6452
rect 151320 6440 151326 6452
rect 151357 6443 151415 6449
rect 151357 6440 151369 6443
rect 151320 6412 151369 6440
rect 151320 6400 151326 6412
rect 151357 6409 151369 6412
rect 151403 6409 151415 6443
rect 151357 6403 151415 6409
rect 151446 6400 151452 6452
rect 151504 6440 151510 6452
rect 152366 6440 152372 6452
rect 151504 6412 152372 6440
rect 151504 6400 151510 6412
rect 152366 6400 152372 6412
rect 152424 6400 152430 6452
rect 153562 6400 153568 6452
rect 153620 6440 153626 6452
rect 156322 6440 156328 6452
rect 153620 6412 156328 6440
rect 153620 6400 153626 6412
rect 156322 6400 156328 6412
rect 156380 6400 156386 6452
rect 159450 6400 159456 6452
rect 159508 6440 159514 6452
rect 184842 6440 184848 6452
rect 159508 6412 184848 6440
rect 159508 6400 159514 6412
rect 184842 6400 184848 6412
rect 184900 6400 184906 6452
rect 188798 6400 188804 6452
rect 188856 6440 188862 6452
rect 188856 6412 189212 6440
rect 188856 6400 188862 6412
rect 107151 6344 109724 6372
rect 107151 6341 107163 6344
rect 107105 6335 107163 6341
rect 98411 6276 98960 6304
rect 99469 6307 99527 6313
rect 98411 6273 98423 6276
rect 98365 6267 98423 6273
rect 99469 6273 99481 6307
rect 99515 6304 99527 6307
rect 99558 6304 99564 6316
rect 99515 6276 99564 6304
rect 99515 6273 99527 6276
rect 99469 6267 99527 6273
rect 99558 6264 99564 6276
rect 99616 6264 99622 6316
rect 99837 6307 99895 6313
rect 99837 6273 99849 6307
rect 99883 6304 99895 6307
rect 100386 6304 100392 6316
rect 99883 6276 100392 6304
rect 99883 6273 99895 6276
rect 99837 6267 99895 6273
rect 100386 6264 100392 6276
rect 100444 6264 100450 6316
rect 100662 6264 100668 6316
rect 100720 6264 100726 6316
rect 101030 6264 101036 6316
rect 101088 6304 101094 6316
rect 101125 6307 101183 6313
rect 101125 6304 101137 6307
rect 101088 6276 101137 6304
rect 101088 6264 101094 6276
rect 101125 6273 101137 6276
rect 101171 6273 101183 6307
rect 101125 6267 101183 6273
rect 101309 6307 101367 6313
rect 101309 6273 101321 6307
rect 101355 6304 101367 6307
rect 101490 6304 101496 6316
rect 101355 6276 101496 6304
rect 101355 6273 101367 6276
rect 101309 6267 101367 6273
rect 101490 6264 101496 6276
rect 101548 6264 101554 6316
rect 101858 6264 101864 6316
rect 101916 6302 101922 6316
rect 101953 6307 102011 6313
rect 101953 6302 101965 6307
rect 101916 6274 101965 6302
rect 101916 6264 101922 6274
rect 101953 6273 101965 6274
rect 101999 6273 102011 6307
rect 101953 6267 102011 6273
rect 102042 6264 102048 6316
rect 102100 6304 102106 6316
rect 103057 6307 103115 6313
rect 103057 6304 103069 6307
rect 102100 6276 103069 6304
rect 102100 6264 102106 6276
rect 103057 6273 103069 6276
rect 103103 6273 103115 6307
rect 103057 6267 103115 6273
rect 104618 6264 104624 6316
rect 104676 6264 104682 6316
rect 105630 6264 105636 6316
rect 105688 6264 105694 6316
rect 106277 6307 106335 6313
rect 106277 6273 106289 6307
rect 106323 6304 106335 6307
rect 106458 6304 106464 6316
rect 106323 6276 106464 6304
rect 106323 6273 106335 6276
rect 106277 6267 106335 6273
rect 106458 6264 106464 6276
rect 106516 6264 106522 6316
rect 53098 6196 53104 6248
rect 53156 6196 53162 6248
rect 91094 6196 91100 6248
rect 91152 6236 91158 6248
rect 91741 6239 91799 6245
rect 91741 6236 91753 6239
rect 91152 6208 91753 6236
rect 91152 6196 91158 6208
rect 91741 6205 91753 6208
rect 91787 6205 91799 6239
rect 91741 6199 91799 6205
rect 92658 6196 92664 6248
rect 92716 6196 92722 6248
rect 92799 6239 92857 6245
rect 92799 6205 92811 6239
rect 92845 6236 92857 6239
rect 93581 6239 93639 6245
rect 92845 6208 93532 6236
rect 92845 6205 92857 6208
rect 92799 6199 92857 6205
rect 53742 6168 53748 6180
rect 52932 6140 53748 6168
rect 48096 6128 48102 6140
rect 53742 6128 53748 6140
rect 53800 6128 53806 6180
rect 92385 6171 92443 6177
rect 92385 6137 92397 6171
rect 92431 6137 92443 6171
rect 93504 6168 93532 6208
rect 93581 6205 93593 6239
rect 93627 6236 93639 6239
rect 95329 6239 95387 6245
rect 95329 6236 95341 6239
rect 93627 6208 95341 6236
rect 93627 6205 93639 6208
rect 93581 6199 93639 6205
rect 95329 6205 95341 6208
rect 95375 6205 95387 6239
rect 95329 6199 95387 6205
rect 96890 6196 96896 6248
rect 96948 6196 96954 6248
rect 97350 6196 97356 6248
rect 97408 6236 97414 6248
rect 98454 6236 98460 6248
rect 97408 6208 98460 6236
rect 97408 6196 97414 6208
rect 98454 6196 98460 6208
rect 98512 6196 98518 6248
rect 99374 6196 99380 6248
rect 99432 6236 99438 6248
rect 107120 6236 107148 6335
rect 109770 6332 109776 6384
rect 109828 6332 109834 6384
rect 111429 6375 111487 6381
rect 111429 6341 111441 6375
rect 111475 6372 111487 6375
rect 113266 6372 113272 6384
rect 111475 6344 113272 6372
rect 111475 6341 111487 6344
rect 111429 6335 111487 6341
rect 113266 6332 113272 6344
rect 113324 6332 113330 6384
rect 113542 6332 113548 6384
rect 113600 6372 113606 6384
rect 132862 6372 132868 6384
rect 113600 6344 115244 6372
rect 113600 6332 113606 6344
rect 107749 6307 107807 6313
rect 107749 6273 107761 6307
rect 107795 6304 107807 6307
rect 108574 6304 108580 6316
rect 107795 6276 108580 6304
rect 107795 6273 107807 6276
rect 107749 6267 107807 6273
rect 107764 6236 107792 6267
rect 108574 6264 108580 6276
rect 108632 6264 108638 6316
rect 109586 6264 109592 6316
rect 109644 6264 109650 6316
rect 112073 6307 112131 6313
rect 112073 6304 112085 6307
rect 110984 6276 112085 6304
rect 99432 6208 107148 6236
rect 107212 6208 107792 6236
rect 107841 6239 107899 6245
rect 99432 6196 99438 6208
rect 101493 6171 101551 6177
rect 93504 6140 95372 6168
rect 92385 6131 92443 6137
rect 18690 6060 18696 6112
rect 18748 6100 18754 6112
rect 51534 6100 51540 6112
rect 18748 6072 51540 6100
rect 18748 6060 18754 6072
rect 51534 6060 51540 6072
rect 51592 6060 51598 6112
rect 92198 6060 92204 6112
rect 92256 6100 92262 6112
rect 92400 6100 92428 6131
rect 93854 6100 93860 6112
rect 92256 6072 93860 6100
rect 92256 6060 92262 6072
rect 93854 6060 93860 6072
rect 93912 6100 93918 6112
rect 94130 6100 94136 6112
rect 93912 6072 94136 6100
rect 93912 6060 93918 6072
rect 94130 6060 94136 6072
rect 94188 6060 94194 6112
rect 94685 6103 94743 6109
rect 94685 6069 94697 6103
rect 94731 6100 94743 6103
rect 94774 6100 94780 6112
rect 94731 6072 94780 6100
rect 94731 6069 94743 6072
rect 94685 6063 94743 6069
rect 94774 6060 94780 6072
rect 94832 6060 94838 6112
rect 95344 6100 95372 6140
rect 95528 6140 101444 6168
rect 95528 6100 95556 6140
rect 95344 6072 95556 6100
rect 96062 6060 96068 6112
rect 96120 6100 96126 6112
rect 97442 6100 97448 6112
rect 96120 6072 97448 6100
rect 96120 6060 96126 6072
rect 97442 6060 97448 6072
rect 97500 6060 97506 6112
rect 97718 6060 97724 6112
rect 97776 6060 97782 6112
rect 97994 6060 98000 6112
rect 98052 6100 98058 6112
rect 98365 6103 98423 6109
rect 98365 6100 98377 6103
rect 98052 6072 98377 6100
rect 98052 6060 98058 6072
rect 98365 6069 98377 6072
rect 98411 6069 98423 6103
rect 98365 6063 98423 6069
rect 99466 6060 99472 6112
rect 99524 6100 99530 6112
rect 99561 6103 99619 6109
rect 99561 6100 99573 6103
rect 99524 6072 99573 6100
rect 99524 6060 99530 6072
rect 99561 6069 99573 6072
rect 99607 6069 99619 6103
rect 99561 6063 99619 6069
rect 99742 6060 99748 6112
rect 99800 6100 99806 6112
rect 100481 6103 100539 6109
rect 100481 6100 100493 6103
rect 99800 6072 100493 6100
rect 99800 6060 99806 6072
rect 100481 6069 100493 6072
rect 100527 6069 100539 6103
rect 100481 6063 100539 6069
rect 100938 6060 100944 6112
rect 100996 6100 101002 6112
rect 101125 6103 101183 6109
rect 101125 6100 101137 6103
rect 100996 6072 101137 6100
rect 100996 6060 101002 6072
rect 101125 6069 101137 6072
rect 101171 6069 101183 6103
rect 101416 6100 101444 6140
rect 101493 6137 101505 6171
rect 101539 6168 101551 6171
rect 101674 6168 101680 6180
rect 101539 6140 101680 6168
rect 101539 6137 101551 6140
rect 101493 6131 101551 6137
rect 101674 6128 101680 6140
rect 101732 6128 101738 6180
rect 104437 6171 104495 6177
rect 104437 6168 104449 6171
rect 101784 6140 104449 6168
rect 101784 6100 101812 6140
rect 104437 6137 104449 6140
rect 104483 6137 104495 6171
rect 104437 6131 104495 6137
rect 104526 6128 104532 6180
rect 104584 6168 104590 6180
rect 107212 6168 107240 6208
rect 107841 6205 107853 6239
rect 107887 6236 107899 6239
rect 108666 6236 108672 6248
rect 107887 6208 108672 6236
rect 107887 6205 107899 6208
rect 107841 6199 107899 6205
rect 108666 6196 108672 6208
rect 108724 6196 108730 6248
rect 109310 6196 109316 6248
rect 109368 6236 109374 6248
rect 110984 6236 111012 6276
rect 112073 6273 112085 6276
rect 112119 6273 112131 6307
rect 112073 6267 112131 6273
rect 112993 6307 113051 6313
rect 112993 6273 113005 6307
rect 113039 6273 113051 6307
rect 112993 6267 113051 6273
rect 109368 6208 111012 6236
rect 113008 6236 113036 6267
rect 113450 6264 113456 6316
rect 113508 6264 113514 6316
rect 113726 6264 113732 6316
rect 113784 6264 113790 6316
rect 115014 6264 115020 6316
rect 115072 6264 115078 6316
rect 115216 6304 115244 6344
rect 117516 6344 120120 6372
rect 115216 6276 115336 6304
rect 115201 6239 115259 6245
rect 113008 6220 113772 6236
rect 113008 6208 113956 6220
rect 109368 6196 109374 6208
rect 113744 6192 113956 6208
rect 115201 6205 115213 6239
rect 115247 6205 115259 6239
rect 115308 6236 115336 6276
rect 115934 6264 115940 6316
rect 115992 6264 115998 6316
rect 117516 6304 117544 6344
rect 116780 6302 117544 6304
rect 117593 6307 117651 6313
rect 117593 6302 117605 6307
rect 116780 6276 117605 6302
rect 116118 6245 116124 6248
rect 115661 6239 115719 6245
rect 115661 6236 115673 6239
rect 115308 6208 115673 6236
rect 115201 6199 115259 6205
rect 115661 6205 115673 6208
rect 115707 6205 115719 6239
rect 115661 6199 115719 6205
rect 116075 6239 116124 6245
rect 116075 6205 116087 6239
rect 116121 6205 116124 6239
rect 116075 6199 116124 6205
rect 104584 6140 107240 6168
rect 107289 6171 107347 6177
rect 104584 6128 104590 6140
rect 107289 6137 107301 6171
rect 107335 6168 107347 6171
rect 107378 6168 107384 6180
rect 107335 6140 107384 6168
rect 107335 6137 107347 6140
rect 107289 6131 107347 6137
rect 107378 6128 107384 6140
rect 107436 6128 107442 6180
rect 108206 6128 108212 6180
rect 108264 6168 108270 6180
rect 113450 6168 113456 6180
rect 108264 6140 113456 6168
rect 108264 6128 108270 6140
rect 113450 6128 113456 6140
rect 113508 6128 113514 6180
rect 113928 6168 113956 6192
rect 114005 6171 114063 6177
rect 114005 6168 114017 6171
rect 113928 6140 114017 6168
rect 114005 6137 114017 6140
rect 114051 6137 114063 6171
rect 114005 6131 114063 6137
rect 115014 6128 115020 6180
rect 115072 6168 115078 6180
rect 115216 6168 115244 6199
rect 115072 6140 115244 6168
rect 115072 6128 115078 6140
rect 101416 6072 101812 6100
rect 101125 6063 101183 6069
rect 101858 6060 101864 6112
rect 101916 6100 101922 6112
rect 101953 6103 102011 6109
rect 101953 6100 101965 6103
rect 101916 6072 101965 6100
rect 101916 6060 101922 6072
rect 101953 6069 101965 6072
rect 101999 6069 102011 6103
rect 101953 6063 102011 6069
rect 103514 6060 103520 6112
rect 103572 6100 103578 6112
rect 103701 6103 103759 6109
rect 103701 6100 103713 6103
rect 103572 6072 103713 6100
rect 103572 6060 103578 6072
rect 103701 6069 103713 6072
rect 103747 6069 103759 6103
rect 103701 6063 103759 6069
rect 103790 6060 103796 6112
rect 103848 6100 103854 6112
rect 105449 6103 105507 6109
rect 105449 6100 105461 6103
rect 103848 6072 105461 6100
rect 103848 6060 103854 6072
rect 105449 6069 105461 6072
rect 105495 6069 105507 6103
rect 105449 6063 105507 6069
rect 105906 6060 105912 6112
rect 105964 6100 105970 6112
rect 106093 6103 106151 6109
rect 106093 6100 106105 6103
rect 105964 6072 106105 6100
rect 105964 6060 105970 6072
rect 106093 6069 106105 6072
rect 106139 6069 106151 6103
rect 106093 6063 106151 6069
rect 107933 6103 107991 6109
rect 107933 6069 107945 6103
rect 107979 6100 107991 6103
rect 108758 6100 108764 6112
rect 107979 6072 108764 6100
rect 107979 6069 107991 6072
rect 107933 6063 107991 6069
rect 108758 6060 108764 6072
rect 108816 6060 108822 6112
rect 108942 6060 108948 6112
rect 109000 6060 109006 6112
rect 111889 6103 111947 6109
rect 111889 6069 111901 6103
rect 111935 6100 111947 6103
rect 112254 6100 112260 6112
rect 111935 6072 112260 6100
rect 111935 6069 111947 6072
rect 111889 6063 111947 6069
rect 112254 6060 112260 6072
rect 112312 6060 112318 6112
rect 112714 6060 112720 6112
rect 112772 6100 112778 6112
rect 113545 6103 113603 6109
rect 113545 6100 113557 6103
rect 112772 6072 113557 6100
rect 112772 6060 112778 6072
rect 113545 6069 113557 6072
rect 113591 6100 113603 6103
rect 114646 6100 114652 6112
rect 113591 6072 114652 6100
rect 113591 6069 113603 6072
rect 113545 6063 113603 6069
rect 114646 6060 114652 6072
rect 114704 6060 114710 6112
rect 115676 6100 115704 6199
rect 116118 6196 116124 6199
rect 116176 6196 116182 6248
rect 116223 6239 116281 6245
rect 116223 6205 116235 6239
rect 116269 6236 116281 6239
rect 116394 6236 116400 6248
rect 116269 6208 116400 6236
rect 116269 6205 116281 6208
rect 116223 6199 116281 6205
rect 116394 6196 116400 6208
rect 116452 6196 116458 6248
rect 116578 6196 116584 6248
rect 116636 6236 116642 6248
rect 116780 6236 116808 6276
rect 117516 6274 117605 6276
rect 117593 6273 117605 6274
rect 117639 6273 117651 6307
rect 118789 6307 118847 6313
rect 118789 6304 118801 6307
rect 117593 6267 117651 6273
rect 117700 6276 118801 6304
rect 116636 6208 116808 6236
rect 116636 6196 116642 6208
rect 116854 6196 116860 6248
rect 116912 6236 116918 6248
rect 117700 6236 117728 6276
rect 118789 6273 118801 6276
rect 118835 6273 118847 6307
rect 118789 6267 118847 6273
rect 116912 6208 117728 6236
rect 116912 6196 116918 6208
rect 117866 6196 117872 6248
rect 117924 6196 117930 6248
rect 118418 6196 118424 6248
rect 118476 6236 118482 6248
rect 118605 6239 118663 6245
rect 118605 6236 118617 6239
rect 118476 6208 118617 6236
rect 118476 6196 118482 6208
rect 118605 6205 118617 6208
rect 118651 6236 118663 6239
rect 118694 6236 118700 6248
rect 118651 6208 118700 6236
rect 118651 6205 118663 6208
rect 118605 6199 118663 6205
rect 118694 6196 118700 6208
rect 118752 6196 118758 6248
rect 116596 6140 118004 6168
rect 116210 6100 116216 6112
rect 115676 6072 116216 6100
rect 116210 6060 116216 6072
rect 116268 6060 116274 6112
rect 116394 6060 116400 6112
rect 116452 6100 116458 6112
rect 116596 6100 116624 6140
rect 116452 6072 116624 6100
rect 116857 6103 116915 6109
rect 116452 6060 116458 6072
rect 116857 6069 116869 6103
rect 116903 6100 116915 6103
rect 117314 6100 117320 6112
rect 116903 6072 117320 6100
rect 116903 6069 116915 6072
rect 116857 6063 116915 6069
rect 117314 6060 117320 6072
rect 117372 6060 117378 6112
rect 117976 6109 118004 6140
rect 117961 6103 118019 6109
rect 117961 6069 117973 6103
rect 118007 6100 118019 6103
rect 118142 6100 118148 6112
rect 118007 6072 118148 6100
rect 118007 6069 118019 6072
rect 117961 6063 118019 6069
rect 118142 6060 118148 6072
rect 118200 6060 118206 6112
rect 118804 6100 118832 6267
rect 118878 6264 118884 6316
rect 118936 6304 118942 6316
rect 120092 6304 120120 6344
rect 125566 6344 132868 6372
rect 125566 6304 125594 6344
rect 132862 6332 132868 6344
rect 132920 6372 132926 6384
rect 141513 6375 141571 6381
rect 141513 6372 141525 6375
rect 132920 6344 141525 6372
rect 132920 6332 132926 6344
rect 141513 6341 141525 6344
rect 141559 6372 141571 6375
rect 162118 6372 162124 6384
rect 141559 6344 162124 6372
rect 141559 6341 141571 6344
rect 141513 6335 141571 6341
rect 162118 6332 162124 6344
rect 162176 6332 162182 6384
rect 168006 6332 168012 6384
rect 168064 6372 168070 6384
rect 189184 6381 189212 6412
rect 189350 6400 189356 6452
rect 189408 6400 189414 6452
rect 189442 6400 189448 6452
rect 189500 6400 189506 6452
rect 189718 6400 189724 6452
rect 189776 6400 189782 6452
rect 189810 6400 189816 6452
rect 189868 6440 189874 6452
rect 216401 6443 216459 6449
rect 216401 6440 216413 6443
rect 189868 6412 216413 6440
rect 189868 6400 189874 6412
rect 216401 6409 216413 6412
rect 216447 6440 216459 6443
rect 216490 6440 216496 6452
rect 216447 6412 216496 6440
rect 216447 6409 216459 6412
rect 216401 6403 216459 6409
rect 216490 6400 216496 6412
rect 216548 6400 216554 6452
rect 216582 6400 216588 6452
rect 216640 6440 216646 6452
rect 222194 6440 222200 6452
rect 216640 6412 222200 6440
rect 216640 6400 216646 6412
rect 222194 6400 222200 6412
rect 222252 6400 222258 6452
rect 224957 6443 225015 6449
rect 224957 6409 224969 6443
rect 225003 6440 225015 6443
rect 226150 6440 226156 6452
rect 225003 6412 226156 6440
rect 225003 6409 225015 6412
rect 224957 6403 225015 6409
rect 226150 6400 226156 6412
rect 226208 6400 226214 6452
rect 226242 6400 226248 6452
rect 226300 6440 226306 6452
rect 248322 6440 248328 6452
rect 226300 6412 248328 6440
rect 226300 6400 226306 6412
rect 248322 6400 248328 6412
rect 248380 6400 248386 6452
rect 249334 6400 249340 6452
rect 249392 6400 249398 6452
rect 253106 6400 253112 6452
rect 253164 6400 253170 6452
rect 254673 6443 254731 6449
rect 254673 6409 254685 6443
rect 254719 6440 254731 6443
rect 255314 6440 255320 6452
rect 254719 6412 255320 6440
rect 254719 6409 254731 6412
rect 254673 6403 254731 6409
rect 255314 6400 255320 6412
rect 255372 6400 255378 6452
rect 255590 6400 255596 6452
rect 255648 6440 255654 6452
rect 255777 6443 255835 6449
rect 255777 6440 255789 6443
rect 255648 6412 255789 6440
rect 255648 6400 255654 6412
rect 255777 6409 255789 6412
rect 255823 6409 255835 6443
rect 255777 6403 255835 6409
rect 256694 6400 256700 6452
rect 256752 6400 256758 6452
rect 261938 6400 261944 6452
rect 261996 6440 262002 6452
rect 264790 6440 264796 6452
rect 261996 6412 264796 6440
rect 261996 6400 262002 6412
rect 264790 6400 264796 6412
rect 264848 6400 264854 6452
rect 266814 6400 266820 6452
rect 266872 6440 266878 6452
rect 269114 6440 269120 6452
rect 266872 6412 269120 6440
rect 266872 6400 266878 6412
rect 269114 6400 269120 6412
rect 269172 6400 269178 6452
rect 270862 6440 270868 6452
rect 270420 6412 270868 6440
rect 168745 6375 168803 6381
rect 168745 6372 168757 6375
rect 168064 6344 168757 6372
rect 168064 6332 168070 6344
rect 168745 6341 168757 6344
rect 168791 6372 168803 6375
rect 169941 6375 169999 6381
rect 169941 6372 169953 6375
rect 168791 6344 169953 6372
rect 168791 6341 168803 6344
rect 168745 6335 168803 6341
rect 169941 6341 169953 6344
rect 169987 6341 169999 6375
rect 169941 6335 169999 6341
rect 189169 6375 189227 6381
rect 189169 6341 189181 6375
rect 189215 6341 189227 6375
rect 189460 6372 189488 6400
rect 189994 6372 190000 6384
rect 189460 6344 190000 6372
rect 189169 6335 189227 6341
rect 189994 6332 190000 6344
rect 190052 6332 190058 6384
rect 216030 6332 216036 6384
rect 216088 6372 216094 6384
rect 217318 6372 217324 6384
rect 216088 6344 217324 6372
rect 216088 6332 216094 6344
rect 217318 6332 217324 6344
rect 217376 6332 217382 6384
rect 221550 6332 221556 6384
rect 221608 6372 221614 6384
rect 224402 6372 224408 6384
rect 221608 6344 224408 6372
rect 221608 6332 221614 6344
rect 224402 6332 224408 6344
rect 224460 6332 224466 6384
rect 231394 6332 231400 6384
rect 231452 6372 231458 6384
rect 245102 6372 245108 6384
rect 231452 6344 245108 6372
rect 231452 6332 231458 6344
rect 245102 6332 245108 6344
rect 245160 6332 245166 6384
rect 255222 6372 255228 6384
rect 245212 6344 250668 6372
rect 118936 6276 119016 6304
rect 120092 6276 125594 6304
rect 135349 6307 135407 6313
rect 118936 6264 118942 6276
rect 118988 6168 119016 6276
rect 135349 6273 135361 6307
rect 135395 6304 135407 6307
rect 135395 6276 136956 6304
rect 135395 6273 135407 6276
rect 135349 6267 135407 6273
rect 119062 6196 119068 6248
rect 119120 6236 119126 6248
rect 130378 6236 130384 6248
rect 119120 6208 130384 6236
rect 119120 6196 119126 6208
rect 130378 6196 130384 6208
rect 130436 6196 130442 6248
rect 135530 6196 135536 6248
rect 135588 6196 135594 6248
rect 136928 6236 136956 6276
rect 137002 6264 137008 6316
rect 137060 6264 137066 6316
rect 138658 6304 138664 6316
rect 137112 6276 138664 6304
rect 137112 6236 137140 6276
rect 138658 6264 138664 6276
rect 138716 6264 138722 6316
rect 140038 6264 140044 6316
rect 140096 6304 140102 6316
rect 140501 6307 140559 6313
rect 140501 6304 140513 6307
rect 140096 6276 140513 6304
rect 140096 6264 140102 6276
rect 140501 6273 140513 6276
rect 140547 6304 140559 6307
rect 142249 6307 142307 6313
rect 142249 6304 142261 6307
rect 140547 6276 142261 6304
rect 140547 6273 140559 6276
rect 140501 6267 140559 6273
rect 142249 6273 142261 6276
rect 142295 6273 142307 6307
rect 142249 6267 142307 6273
rect 150253 6307 150311 6313
rect 150253 6273 150265 6307
rect 150299 6302 150311 6307
rect 150299 6274 150388 6302
rect 150299 6273 150311 6274
rect 150253 6267 150311 6273
rect 136928 6208 137140 6236
rect 137186 6196 137192 6248
rect 137244 6196 137250 6248
rect 139578 6196 139584 6248
rect 139636 6236 139642 6248
rect 140777 6239 140835 6245
rect 140777 6236 140789 6239
rect 139636 6208 140789 6236
rect 139636 6196 139642 6208
rect 140777 6205 140789 6208
rect 140823 6236 140835 6239
rect 150158 6236 150164 6248
rect 140823 6208 150164 6236
rect 140823 6205 140835 6208
rect 140777 6199 140835 6205
rect 150158 6196 150164 6208
rect 150216 6196 150222 6248
rect 120534 6168 120540 6180
rect 118988 6140 120540 6168
rect 120534 6128 120540 6140
rect 120592 6128 120598 6180
rect 142798 6168 142804 6180
rect 128326 6140 142804 6168
rect 119890 6100 119896 6112
rect 118804 6072 119896 6100
rect 119890 6060 119896 6072
rect 119948 6100 119954 6112
rect 128326 6100 128354 6140
rect 142798 6128 142804 6140
rect 142856 6128 142862 6180
rect 150360 6168 150388 6274
rect 150618 6264 150624 6316
rect 150676 6304 150682 6316
rect 150805 6307 150863 6313
rect 150805 6304 150817 6307
rect 150676 6276 150817 6304
rect 150676 6264 150682 6276
rect 150805 6273 150817 6276
rect 150851 6304 150863 6307
rect 151817 6307 151875 6313
rect 151817 6304 151829 6307
rect 150851 6276 151829 6304
rect 150851 6273 150863 6276
rect 150805 6267 150863 6273
rect 151817 6273 151829 6276
rect 151863 6273 151875 6307
rect 152550 6304 152556 6316
rect 151817 6267 151875 6273
rect 152108 6276 152556 6304
rect 150986 6196 150992 6248
rect 151044 6236 151050 6248
rect 151081 6239 151139 6245
rect 151081 6236 151093 6239
rect 151044 6208 151093 6236
rect 151044 6196 151050 6208
rect 151081 6205 151093 6208
rect 151127 6236 151139 6239
rect 151538 6236 151544 6248
rect 151127 6208 151544 6236
rect 151127 6205 151139 6208
rect 151081 6199 151139 6205
rect 151538 6196 151544 6208
rect 151596 6236 151602 6248
rect 152108 6245 152136 6276
rect 152550 6264 152556 6276
rect 152608 6264 152614 6316
rect 152829 6307 152887 6313
rect 152829 6273 152841 6307
rect 152875 6304 152887 6307
rect 153746 6304 153752 6316
rect 152875 6276 153752 6304
rect 152875 6273 152887 6276
rect 152829 6267 152887 6273
rect 153746 6264 153752 6276
rect 153804 6264 153810 6316
rect 153841 6307 153899 6313
rect 153841 6273 153853 6307
rect 153887 6273 153899 6307
rect 153841 6267 153899 6273
rect 152093 6239 152151 6245
rect 152093 6236 152105 6239
rect 151596 6208 152105 6236
rect 151596 6196 151602 6208
rect 152093 6205 152105 6208
rect 152139 6205 152151 6239
rect 152093 6199 152151 6205
rect 152274 6196 152280 6248
rect 152332 6236 152338 6248
rect 153013 6239 153071 6245
rect 153013 6236 153025 6239
rect 152332 6208 153025 6236
rect 152332 6196 152338 6208
rect 153013 6205 153025 6208
rect 153059 6205 153071 6239
rect 153856 6236 153884 6267
rect 154850 6264 154856 6316
rect 154908 6264 154914 6316
rect 156138 6264 156144 6316
rect 156196 6264 156202 6316
rect 161198 6304 161204 6316
rect 156248 6276 161204 6304
rect 154942 6236 154948 6248
rect 153856 6208 154948 6236
rect 153013 6199 153071 6205
rect 154942 6196 154948 6208
rect 155000 6196 155006 6248
rect 155862 6196 155868 6248
rect 155920 6236 155926 6248
rect 156248 6236 156276 6276
rect 161198 6264 161204 6276
rect 161256 6264 161262 6316
rect 161290 6264 161296 6316
rect 161348 6304 161354 6316
rect 168101 6307 168159 6313
rect 168101 6304 168113 6307
rect 161348 6276 168113 6304
rect 161348 6264 161354 6276
rect 168101 6273 168113 6276
rect 168147 6304 168159 6307
rect 168377 6307 168435 6313
rect 168377 6304 168389 6307
rect 168147 6276 168389 6304
rect 168147 6273 168159 6276
rect 168101 6267 168159 6273
rect 168377 6273 168389 6276
rect 168423 6304 168435 6307
rect 169573 6307 169631 6313
rect 168423 6276 169524 6304
rect 168423 6273 168435 6276
rect 168377 6267 168435 6273
rect 155920 6208 156276 6236
rect 155920 6196 155926 6208
rect 156322 6196 156328 6248
rect 156380 6236 156386 6248
rect 161658 6236 161664 6248
rect 156380 6208 161664 6236
rect 156380 6196 156386 6208
rect 161658 6196 161664 6208
rect 161716 6196 161722 6248
rect 162854 6196 162860 6248
rect 162912 6236 162918 6248
rect 165706 6236 165712 6248
rect 162912 6208 165712 6236
rect 162912 6196 162918 6208
rect 165706 6196 165712 6208
rect 165764 6196 165770 6248
rect 168650 6196 168656 6248
rect 168708 6196 168714 6248
rect 168862 6239 168920 6245
rect 168862 6236 168874 6239
rect 168852 6205 168874 6236
rect 168908 6236 168920 6239
rect 168908 6208 169432 6236
rect 168908 6205 168920 6208
rect 168852 6199 168920 6205
rect 152369 6171 152427 6177
rect 152369 6168 152381 6171
rect 150360 6140 152381 6168
rect 152369 6137 152381 6140
rect 152415 6137 152427 6171
rect 152369 6131 152427 6137
rect 153746 6128 153752 6180
rect 153804 6168 153810 6180
rect 155957 6171 156015 6177
rect 153804 6140 155908 6168
rect 153804 6128 153810 6140
rect 119948 6072 128354 6100
rect 119948 6060 119954 6072
rect 137002 6060 137008 6112
rect 137060 6100 137066 6112
rect 139946 6100 139952 6112
rect 137060 6072 139952 6100
rect 137060 6060 137066 6072
rect 139946 6060 139952 6072
rect 140004 6060 140010 6112
rect 141605 6103 141663 6109
rect 141605 6069 141617 6103
rect 141651 6100 141663 6103
rect 142246 6100 142252 6112
rect 141651 6072 142252 6100
rect 141651 6069 141663 6072
rect 141605 6063 141663 6069
rect 142246 6060 142252 6072
rect 142304 6060 142310 6112
rect 142341 6103 142399 6109
rect 142341 6069 142353 6103
rect 142387 6100 142399 6103
rect 143166 6100 143172 6112
rect 142387 6072 143172 6100
rect 142387 6069 142399 6072
rect 142341 6063 142399 6069
rect 143166 6060 143172 6072
rect 143224 6100 143230 6112
rect 149054 6100 149060 6112
rect 143224 6072 149060 6100
rect 143224 6060 143230 6072
rect 149054 6060 149060 6072
rect 149112 6060 149118 6112
rect 150066 6060 150072 6112
rect 150124 6060 150130 6112
rect 150894 6060 150900 6112
rect 150952 6100 150958 6112
rect 151909 6103 151967 6109
rect 151909 6100 151921 6103
rect 150952 6072 151921 6100
rect 150952 6060 150958 6072
rect 151909 6069 151921 6072
rect 151955 6069 151967 6103
rect 151909 6063 151967 6069
rect 152734 6060 152740 6112
rect 152792 6100 152798 6112
rect 153933 6103 153991 6109
rect 153933 6100 153945 6103
rect 152792 6072 153945 6100
rect 152792 6060 152798 6072
rect 153933 6069 153945 6072
rect 153979 6069 153991 6103
rect 153933 6063 153991 6069
rect 154669 6103 154727 6109
rect 154669 6069 154681 6103
rect 154715 6100 154727 6103
rect 155770 6100 155776 6112
rect 154715 6072 155776 6100
rect 154715 6069 154727 6072
rect 154669 6063 154727 6069
rect 155770 6060 155776 6072
rect 155828 6060 155834 6112
rect 155880 6100 155908 6140
rect 155957 6137 155969 6171
rect 156003 6168 156015 6171
rect 158438 6168 158444 6180
rect 156003 6140 158444 6168
rect 156003 6137 156015 6140
rect 155957 6131 156015 6137
rect 158438 6128 158444 6140
rect 158496 6128 158502 6180
rect 167730 6128 167736 6180
rect 167788 6168 167794 6180
rect 168852 6168 168880 6199
rect 167788 6140 168880 6168
rect 167788 6128 167794 6140
rect 169018 6128 169024 6180
rect 169076 6128 169082 6180
rect 156322 6100 156328 6112
rect 155880 6072 156328 6100
rect 156322 6060 156328 6072
rect 156380 6060 156386 6112
rect 156414 6060 156420 6112
rect 156472 6100 156478 6112
rect 156782 6100 156788 6112
rect 156472 6072 156788 6100
rect 156472 6060 156478 6072
rect 156782 6060 156788 6072
rect 156840 6100 156846 6112
rect 159818 6100 159824 6112
rect 156840 6072 159824 6100
rect 156840 6060 156846 6072
rect 159818 6060 159824 6072
rect 159876 6060 159882 6112
rect 169404 6100 169432 6208
rect 169496 6168 169524 6276
rect 169573 6273 169585 6307
rect 169619 6304 169631 6307
rect 169754 6304 169760 6316
rect 169619 6276 169760 6304
rect 169619 6273 169631 6276
rect 169573 6267 169631 6273
rect 169754 6264 169760 6276
rect 169812 6304 169818 6316
rect 171226 6304 171232 6316
rect 169812 6276 171232 6304
rect 169812 6264 169818 6276
rect 171226 6264 171232 6276
rect 171284 6264 171290 6316
rect 189534 6264 189540 6316
rect 189592 6264 189598 6316
rect 207474 6264 207480 6316
rect 207532 6304 207538 6316
rect 208213 6307 208271 6313
rect 208213 6304 208225 6307
rect 207532 6276 208225 6304
rect 207532 6264 207538 6276
rect 208213 6273 208225 6276
rect 208259 6273 208271 6307
rect 208213 6267 208271 6273
rect 209130 6264 209136 6316
rect 209188 6264 209194 6316
rect 209314 6313 209320 6316
rect 209271 6307 209320 6313
rect 209271 6273 209283 6307
rect 209317 6273 209320 6307
rect 209271 6267 209320 6273
rect 209314 6264 209320 6267
rect 209372 6264 209378 6316
rect 213086 6264 213092 6316
rect 213144 6264 213150 6316
rect 216125 6307 216183 6313
rect 216125 6273 216137 6307
rect 216171 6304 216183 6307
rect 216306 6304 216312 6316
rect 216171 6276 216312 6304
rect 216171 6273 216183 6276
rect 216125 6267 216183 6273
rect 216306 6264 216312 6276
rect 216364 6304 216370 6316
rect 217137 6307 217195 6313
rect 217137 6304 217149 6307
rect 216364 6276 217149 6304
rect 216364 6264 216370 6276
rect 217137 6273 217149 6276
rect 217183 6273 217195 6307
rect 217137 6267 217195 6273
rect 217870 6264 217876 6316
rect 217928 6264 217934 6316
rect 217965 6307 218023 6313
rect 217965 6273 217977 6307
rect 218011 6273 218023 6307
rect 217965 6267 218023 6273
rect 208397 6239 208455 6245
rect 185596 6208 190454 6236
rect 185486 6168 185492 6180
rect 169496 6140 185492 6168
rect 185486 6128 185492 6140
rect 185544 6128 185550 6180
rect 185596 6100 185624 6208
rect 169404 6072 185624 6100
rect 190426 6100 190454 6208
rect 208397 6205 208409 6239
rect 208443 6236 208455 6239
rect 208486 6236 208492 6248
rect 208443 6208 208492 6236
rect 208443 6205 208455 6208
rect 208397 6199 208455 6205
rect 208486 6196 208492 6208
rect 208544 6196 208550 6248
rect 209406 6196 209412 6248
rect 209464 6236 209470 6248
rect 209464 6208 212534 6236
rect 209464 6196 209470 6208
rect 207750 6128 207756 6180
rect 207808 6168 207814 6180
rect 208857 6171 208915 6177
rect 208857 6168 208869 6171
rect 207808 6140 208869 6168
rect 207808 6128 207814 6140
rect 208857 6137 208869 6140
rect 208903 6137 208915 6171
rect 212506 6168 212534 6208
rect 212810 6196 212816 6248
rect 212868 6236 212874 6248
rect 213273 6239 213331 6245
rect 213273 6236 213285 6239
rect 212868 6208 213285 6236
rect 212868 6196 212874 6208
rect 213273 6205 213285 6208
rect 213319 6205 213331 6239
rect 213273 6199 213331 6205
rect 216493 6239 216551 6245
rect 216493 6205 216505 6239
rect 216539 6205 216551 6239
rect 216493 6199 216551 6205
rect 216610 6239 216668 6245
rect 216610 6205 216622 6239
rect 216656 6236 216668 6239
rect 217042 6236 217048 6248
rect 216656 6208 217048 6236
rect 216656 6205 216668 6208
rect 216610 6199 216668 6205
rect 213454 6168 213460 6180
rect 212506 6140 213460 6168
rect 208857 6131 208915 6137
rect 213454 6128 213460 6140
rect 213512 6128 213518 6180
rect 200758 6100 200764 6112
rect 190426 6072 200764 6100
rect 200758 6060 200764 6072
rect 200816 6060 200822 6112
rect 207290 6060 207296 6112
rect 207348 6100 207354 6112
rect 210053 6103 210111 6109
rect 210053 6100 210065 6103
rect 207348 6072 210065 6100
rect 207348 6060 207354 6072
rect 210053 6069 210065 6072
rect 210099 6069 210111 6103
rect 210053 6063 210111 6069
rect 215846 6060 215852 6112
rect 215904 6100 215910 6112
rect 216508 6100 216536 6199
rect 217042 6196 217048 6208
rect 217100 6196 217106 6248
rect 217980 6236 218008 6267
rect 218054 6264 218060 6316
rect 218112 6264 218118 6316
rect 218422 6264 218428 6316
rect 218480 6304 218486 6316
rect 218793 6307 218851 6313
rect 218793 6304 218805 6307
rect 218480 6276 218805 6304
rect 218480 6264 218486 6276
rect 218793 6273 218805 6276
rect 218839 6273 218851 6307
rect 218793 6267 218851 6273
rect 221366 6264 221372 6316
rect 221424 6304 221430 6316
rect 221645 6307 221703 6313
rect 221645 6304 221657 6307
rect 221424 6276 221657 6304
rect 221424 6264 221430 6276
rect 221645 6273 221657 6276
rect 221691 6273 221703 6307
rect 221645 6267 221703 6273
rect 221734 6264 221740 6316
rect 221792 6264 221798 6316
rect 221826 6264 221832 6316
rect 221884 6264 221890 6316
rect 224586 6264 224592 6316
rect 224644 6264 224650 6316
rect 226150 6264 226156 6316
rect 226208 6264 226214 6316
rect 226426 6264 226432 6316
rect 226484 6264 226490 6316
rect 244642 6264 244648 6316
rect 244700 6304 244706 6316
rect 245212 6304 245240 6344
rect 244700 6276 245240 6304
rect 248141 6307 248199 6313
rect 244700 6264 244706 6276
rect 248141 6273 248153 6307
rect 248187 6304 248199 6307
rect 248230 6304 248236 6316
rect 248187 6276 248236 6304
rect 248187 6273 248199 6276
rect 248141 6267 248199 6273
rect 248230 6264 248236 6276
rect 248288 6264 248294 6316
rect 248322 6264 248328 6316
rect 248380 6304 248386 6316
rect 248877 6307 248935 6313
rect 248380 6276 248828 6304
rect 248380 6264 248386 6276
rect 218330 6236 218336 6248
rect 217980 6208 218336 6236
rect 218330 6196 218336 6208
rect 218388 6196 218394 6248
rect 218974 6196 218980 6248
rect 219032 6196 219038 6248
rect 219526 6196 219532 6248
rect 219584 6236 219590 6248
rect 219894 6245 219900 6248
rect 219713 6239 219771 6245
rect 219713 6236 219725 6239
rect 219584 6208 219725 6236
rect 219584 6196 219590 6208
rect 219713 6205 219725 6208
rect 219759 6205 219771 6239
rect 219713 6199 219771 6205
rect 219851 6239 219900 6245
rect 219851 6205 219863 6239
rect 219897 6205 219900 6239
rect 219851 6199 219900 6205
rect 219894 6196 219900 6199
rect 219952 6196 219958 6248
rect 219989 6239 220047 6245
rect 219989 6205 220001 6239
rect 220035 6236 220047 6239
rect 220722 6236 220728 6248
rect 220035 6208 220728 6236
rect 220035 6205 220047 6208
rect 219989 6199 220047 6205
rect 220722 6196 220728 6208
rect 220780 6236 220786 6248
rect 222286 6236 222292 6248
rect 220780 6208 222292 6236
rect 220780 6196 220786 6208
rect 222286 6196 222292 6208
rect 222344 6196 222350 6248
rect 222746 6196 222752 6248
rect 222804 6196 222810 6248
rect 222933 6239 222991 6245
rect 222933 6205 222945 6239
rect 222979 6236 222991 6239
rect 223298 6236 223304 6248
rect 222979 6208 223304 6236
rect 222979 6205 222991 6208
rect 222933 6199 222991 6205
rect 223298 6196 223304 6208
rect 223356 6196 223362 6248
rect 225230 6196 225236 6248
rect 225288 6196 225294 6248
rect 225414 6196 225420 6248
rect 225472 6196 225478 6248
rect 226242 6196 226248 6248
rect 226300 6245 226306 6248
rect 226300 6239 226328 6245
rect 226316 6205 226328 6239
rect 226300 6199 226328 6205
rect 226300 6196 226306 6199
rect 226794 6196 226800 6248
rect 226852 6236 226858 6248
rect 241514 6236 241520 6248
rect 226852 6208 241520 6236
rect 226852 6196 226858 6208
rect 241514 6196 241520 6208
rect 241572 6196 241578 6248
rect 248690 6236 248696 6248
rect 244246 6208 248696 6236
rect 216766 6128 216772 6180
rect 216824 6128 216830 6180
rect 217134 6128 217140 6180
rect 217192 6168 217198 6180
rect 217192 6140 218376 6168
rect 217192 6128 217198 6140
rect 215904 6072 216536 6100
rect 215904 6060 215910 6072
rect 218146 6060 218152 6112
rect 218204 6100 218210 6112
rect 218241 6103 218299 6109
rect 218241 6100 218253 6103
rect 218204 6072 218253 6100
rect 218204 6060 218210 6072
rect 218241 6069 218253 6072
rect 218287 6069 218299 6103
rect 218348 6100 218376 6140
rect 218606 6128 218612 6180
rect 218664 6168 218670 6180
rect 219437 6171 219495 6177
rect 219437 6168 219449 6171
rect 218664 6140 219449 6168
rect 218664 6128 218670 6140
rect 219437 6137 219449 6140
rect 219483 6137 219495 6171
rect 219437 6131 219495 6137
rect 218698 6100 218704 6112
rect 218348 6072 218704 6100
rect 218241 6063 218299 6069
rect 218698 6060 218704 6072
rect 218756 6060 218762 6112
rect 219452 6100 219480 6131
rect 220446 6128 220452 6180
rect 220504 6168 220510 6180
rect 221642 6168 221648 6180
rect 220504 6140 221648 6168
rect 220504 6128 220510 6140
rect 221642 6128 221648 6140
rect 221700 6128 221706 6180
rect 222838 6128 222844 6180
rect 222896 6168 222902 6180
rect 224770 6168 224776 6180
rect 222896 6140 224776 6168
rect 222896 6128 222902 6140
rect 224770 6128 224776 6140
rect 224828 6128 224834 6180
rect 225874 6128 225880 6180
rect 225932 6128 225938 6180
rect 226812 6140 227392 6168
rect 219802 6100 219808 6112
rect 219452 6072 219808 6100
rect 219802 6060 219808 6072
rect 219860 6060 219866 6112
rect 220170 6060 220176 6112
rect 220228 6100 220234 6112
rect 220633 6103 220691 6109
rect 220633 6100 220645 6103
rect 220228 6072 220645 6100
rect 220228 6060 220234 6072
rect 220633 6069 220645 6072
rect 220679 6069 220691 6103
rect 220633 6063 220691 6069
rect 222013 6103 222071 6109
rect 222013 6069 222025 6103
rect 222059 6100 222071 6103
rect 223114 6100 223120 6112
rect 222059 6072 223120 6100
rect 222059 6069 222071 6072
rect 222013 6063 222071 6069
rect 223114 6060 223120 6072
rect 223172 6060 223178 6112
rect 223206 6060 223212 6112
rect 223264 6100 223270 6112
rect 224862 6100 224868 6112
rect 223264 6072 224868 6100
rect 223264 6060 223270 6072
rect 224862 6060 224868 6072
rect 224920 6060 224926 6112
rect 226150 6060 226156 6112
rect 226208 6100 226214 6112
rect 226812 6100 226840 6140
rect 226208 6072 226840 6100
rect 226208 6060 226214 6072
rect 227070 6060 227076 6112
rect 227128 6060 227134 6112
rect 227364 6100 227392 6140
rect 227438 6128 227444 6180
rect 227496 6168 227502 6180
rect 244246 6168 244274 6208
rect 248690 6196 248696 6208
rect 248748 6196 248754 6248
rect 248800 6236 248828 6276
rect 248877 6273 248889 6307
rect 248923 6304 248935 6307
rect 248923 6276 249104 6304
rect 248923 6273 248935 6276
rect 248877 6267 248935 6273
rect 248969 6239 249027 6245
rect 248969 6236 248981 6239
rect 248800 6208 248981 6236
rect 248969 6205 248981 6208
rect 249015 6205 249027 6239
rect 249076 6236 249104 6276
rect 249150 6264 249156 6316
rect 249208 6264 249214 6316
rect 250640 6313 250668 6344
rect 252848 6344 255228 6372
rect 249981 6307 250039 6313
rect 249981 6273 249993 6307
rect 250027 6273 250039 6307
rect 249981 6267 250039 6273
rect 250625 6307 250683 6313
rect 250625 6273 250637 6307
rect 250671 6273 250683 6307
rect 250625 6267 250683 6273
rect 249334 6236 249340 6248
rect 249076 6208 249340 6236
rect 248969 6199 249027 6205
rect 249334 6196 249340 6208
rect 249392 6196 249398 6248
rect 227496 6140 244274 6168
rect 227496 6128 227502 6140
rect 248138 6128 248144 6180
rect 248196 6168 248202 6180
rect 249996 6168 250024 6267
rect 251358 6264 251364 6316
rect 251416 6304 251422 6316
rect 252848 6313 252876 6344
rect 255222 6332 255228 6344
rect 255280 6332 255286 6384
rect 256237 6375 256295 6381
rect 256237 6372 256249 6375
rect 255424 6344 256249 6372
rect 255424 6316 255452 6344
rect 256237 6341 256249 6344
rect 256283 6341 256295 6375
rect 256237 6335 256295 6341
rect 256326 6332 256332 6384
rect 256384 6372 256390 6384
rect 259638 6372 259644 6384
rect 256384 6344 259644 6372
rect 256384 6332 256390 6344
rect 259638 6332 259644 6344
rect 259696 6332 259702 6384
rect 261754 6332 261760 6384
rect 261812 6372 261818 6384
rect 262033 6375 262091 6381
rect 262033 6372 262045 6375
rect 261812 6344 262045 6372
rect 261812 6332 261818 6344
rect 262033 6341 262045 6344
rect 262079 6341 262091 6375
rect 262033 6335 262091 6341
rect 263778 6332 263784 6384
rect 263836 6372 263842 6384
rect 270218 6372 270224 6384
rect 263836 6344 270224 6372
rect 263836 6332 263842 6344
rect 270218 6332 270224 6344
rect 270276 6332 270282 6384
rect 252833 6307 252891 6313
rect 251416 6276 252600 6304
rect 251416 6264 251422 6276
rect 248196 6140 250024 6168
rect 250088 6208 251588 6236
rect 248196 6128 248202 6140
rect 239490 6100 239496 6112
rect 227364 6072 239496 6100
rect 239490 6060 239496 6072
rect 239548 6060 239554 6112
rect 242894 6060 242900 6112
rect 242952 6100 242958 6112
rect 247402 6100 247408 6112
rect 242952 6072 247408 6100
rect 242952 6060 242958 6072
rect 247402 6060 247408 6072
rect 247460 6060 247466 6112
rect 247957 6103 248015 6109
rect 247957 6069 247969 6103
rect 248003 6100 248015 6103
rect 248598 6100 248604 6112
rect 248003 6072 248604 6100
rect 248003 6069 248015 6072
rect 247957 6063 248015 6069
rect 248598 6060 248604 6072
rect 248656 6060 248662 6112
rect 248782 6060 248788 6112
rect 248840 6100 248846 6112
rect 248877 6103 248935 6109
rect 248877 6100 248889 6103
rect 248840 6072 248889 6100
rect 248840 6060 248846 6072
rect 248877 6069 248889 6072
rect 248923 6069 248935 6103
rect 248877 6063 248935 6069
rect 249058 6060 249064 6112
rect 249116 6100 249122 6112
rect 249797 6103 249855 6109
rect 249797 6100 249809 6103
rect 249116 6072 249809 6100
rect 249116 6060 249122 6072
rect 249797 6069 249809 6072
rect 249843 6069 249855 6103
rect 249797 6063 249855 6069
rect 249886 6060 249892 6112
rect 249944 6100 249950 6112
rect 250088 6100 250116 6208
rect 249944 6072 250116 6100
rect 250441 6103 250499 6109
rect 249944 6060 249950 6072
rect 250441 6069 250453 6103
rect 250487 6100 250499 6103
rect 251450 6100 251456 6112
rect 250487 6072 251456 6100
rect 250487 6069 250499 6072
rect 250441 6063 250499 6069
rect 251450 6060 251456 6072
rect 251508 6060 251514 6112
rect 251560 6100 251588 6208
rect 252572 6168 252600 6276
rect 252833 6273 252845 6307
rect 252879 6273 252891 6307
rect 252833 6267 252891 6273
rect 252925 6307 252983 6313
rect 252925 6273 252937 6307
rect 252971 6304 252983 6307
rect 253198 6304 253204 6316
rect 252971 6276 253204 6304
rect 252971 6273 252983 6276
rect 252925 6267 252983 6273
rect 253198 6264 253204 6276
rect 253256 6264 253262 6316
rect 254026 6264 254032 6316
rect 254084 6304 254090 6316
rect 254857 6307 254915 6313
rect 254857 6304 254869 6307
rect 254084 6276 254869 6304
rect 254084 6264 254090 6276
rect 254857 6273 254869 6276
rect 254903 6273 254915 6307
rect 254857 6267 254915 6273
rect 255317 6307 255375 6313
rect 255317 6273 255329 6307
rect 255363 6304 255375 6307
rect 255406 6304 255412 6316
rect 255363 6276 255412 6304
rect 255363 6273 255375 6276
rect 255317 6267 255375 6273
rect 255406 6264 255412 6276
rect 255464 6264 255470 6316
rect 255593 6307 255651 6313
rect 255593 6273 255605 6307
rect 255639 6304 255651 6307
rect 256513 6307 256571 6313
rect 256513 6304 256525 6307
rect 255639 6276 256525 6304
rect 255639 6273 255651 6276
rect 255593 6267 255651 6273
rect 256513 6273 256525 6276
rect 256559 6304 256571 6307
rect 256786 6304 256792 6316
rect 256559 6276 256792 6304
rect 256559 6273 256571 6276
rect 256513 6267 256571 6273
rect 256786 6264 256792 6276
rect 256844 6264 256850 6316
rect 257341 6307 257399 6313
rect 257341 6273 257353 6307
rect 257387 6304 257399 6307
rect 258902 6304 258908 6316
rect 257387 6276 258908 6304
rect 257387 6273 257399 6276
rect 257341 6267 257399 6273
rect 258902 6264 258908 6276
rect 258960 6264 258966 6316
rect 260101 6307 260159 6313
rect 260101 6273 260113 6307
rect 260147 6304 260159 6307
rect 260929 6307 260987 6313
rect 260929 6304 260941 6307
rect 260147 6276 260941 6304
rect 260147 6273 260159 6276
rect 260101 6267 260159 6273
rect 260929 6273 260941 6276
rect 260975 6304 260987 6307
rect 261570 6304 261576 6316
rect 260975 6276 261576 6304
rect 260975 6273 260987 6276
rect 260929 6267 260987 6273
rect 261570 6264 261576 6276
rect 261628 6264 261634 6316
rect 261665 6307 261723 6313
rect 261665 6273 261677 6307
rect 261711 6304 261723 6307
rect 262490 6304 262496 6316
rect 261711 6276 262496 6304
rect 261711 6273 261723 6276
rect 261665 6267 261723 6273
rect 262490 6264 262496 6276
rect 262548 6264 262554 6316
rect 262953 6307 263011 6313
rect 262953 6273 262965 6307
rect 262999 6304 263011 6307
rect 263134 6304 263140 6316
rect 262999 6276 263140 6304
rect 262999 6273 263011 6276
rect 262953 6267 263011 6273
rect 263134 6264 263140 6276
rect 263192 6264 263198 6316
rect 264241 6307 264299 6313
rect 264241 6273 264253 6307
rect 264287 6304 264299 6307
rect 265250 6304 265256 6316
rect 264287 6276 265256 6304
rect 264287 6273 264299 6276
rect 264241 6267 264299 6273
rect 265250 6264 265256 6276
rect 265308 6264 265314 6316
rect 265437 6307 265495 6313
rect 265437 6273 265449 6307
rect 265483 6304 265495 6307
rect 266538 6304 266544 6316
rect 265483 6276 266544 6304
rect 265483 6273 265495 6276
rect 265437 6267 265495 6273
rect 266538 6264 266544 6276
rect 266596 6264 266602 6316
rect 266630 6264 266636 6316
rect 266688 6264 266694 6316
rect 267182 6264 267188 6316
rect 267240 6264 267246 6316
rect 267826 6264 267832 6316
rect 267884 6264 267890 6316
rect 268930 6264 268936 6316
rect 268988 6264 268994 6316
rect 269390 6264 269396 6316
rect 269448 6264 269454 6316
rect 254578 6196 254584 6248
rect 254636 6236 254642 6248
rect 255501 6239 255559 6245
rect 255501 6236 255513 6239
rect 254636 6208 255513 6236
rect 254636 6196 254642 6208
rect 255501 6205 255513 6208
rect 255547 6236 255559 6239
rect 256421 6239 256479 6245
rect 256421 6236 256433 6239
rect 255547 6208 256433 6236
rect 255547 6205 255559 6208
rect 255501 6199 255559 6205
rect 256421 6205 256433 6208
rect 256467 6236 256479 6239
rect 256694 6236 256700 6248
rect 256467 6208 256700 6236
rect 256467 6205 256479 6208
rect 256421 6199 256479 6205
rect 256694 6196 256700 6208
rect 256752 6196 256758 6248
rect 259917 6239 259975 6245
rect 259917 6205 259929 6239
rect 259963 6205 259975 6239
rect 259917 6199 259975 6205
rect 260745 6239 260803 6245
rect 260745 6205 260757 6239
rect 260791 6236 260803 6239
rect 262122 6236 262128 6248
rect 260791 6208 262128 6236
rect 260791 6205 260803 6208
rect 260745 6199 260803 6205
rect 258810 6168 258816 6180
rect 252572 6140 258816 6168
rect 258810 6128 258816 6140
rect 258868 6128 258874 6180
rect 259932 6168 259960 6199
rect 262122 6196 262128 6208
rect 262180 6196 262186 6248
rect 263226 6196 263232 6248
rect 263284 6196 263290 6248
rect 264514 6196 264520 6248
rect 264572 6196 264578 6248
rect 265710 6196 265716 6248
rect 265768 6196 265774 6248
rect 268381 6239 268439 6245
rect 268381 6205 268393 6239
rect 268427 6236 268439 6239
rect 268948 6236 268976 6264
rect 268427 6208 268976 6236
rect 269669 6239 269727 6245
rect 268427 6205 268439 6208
rect 268381 6199 268439 6205
rect 269669 6205 269681 6239
rect 269715 6236 269727 6239
rect 270420 6236 270448 6412
rect 270862 6400 270868 6412
rect 270920 6400 270926 6452
rect 270494 6332 270500 6384
rect 270552 6372 270558 6384
rect 270552 6344 270724 6372
rect 270552 6332 270558 6344
rect 270696 6313 270724 6344
rect 270681 6307 270739 6313
rect 270681 6273 270693 6307
rect 270727 6273 270739 6307
rect 270681 6267 270739 6273
rect 269715 6208 270448 6236
rect 269715 6205 269727 6208
rect 269669 6199 269727 6205
rect 261754 6168 261760 6180
rect 259932 6140 261760 6168
rect 261754 6128 261760 6140
rect 261812 6128 261818 6180
rect 263042 6128 263048 6180
rect 263100 6168 263106 6180
rect 268838 6168 268844 6180
rect 263100 6140 268844 6168
rect 263100 6128 263106 6140
rect 268838 6128 268844 6140
rect 268896 6128 268902 6180
rect 254394 6100 254400 6112
rect 251560 6072 254400 6100
rect 254394 6060 254400 6072
rect 254452 6060 254458 6112
rect 255593 6103 255651 6109
rect 255593 6069 255605 6103
rect 255639 6100 255651 6103
rect 255774 6100 255780 6112
rect 255639 6072 255780 6100
rect 255639 6069 255651 6072
rect 255593 6063 255651 6069
rect 255774 6060 255780 6072
rect 255832 6100 255838 6112
rect 256418 6100 256424 6112
rect 255832 6072 256424 6100
rect 255832 6060 255838 6072
rect 256418 6060 256424 6072
rect 256476 6060 256482 6112
rect 256510 6060 256516 6112
rect 256568 6100 256574 6112
rect 257157 6103 257215 6109
rect 257157 6100 257169 6103
rect 256568 6072 257169 6100
rect 256568 6060 256574 6072
rect 257157 6069 257169 6072
rect 257203 6069 257215 6103
rect 257157 6063 257215 6069
rect 260285 6103 260343 6109
rect 260285 6069 260297 6103
rect 260331 6100 260343 6103
rect 260374 6100 260380 6112
rect 260331 6072 260380 6100
rect 260331 6069 260343 6072
rect 260285 6063 260343 6069
rect 260374 6060 260380 6072
rect 260432 6060 260438 6112
rect 261113 6103 261171 6109
rect 261113 6069 261125 6103
rect 261159 6100 261171 6103
rect 261662 6100 261668 6112
rect 261159 6072 261668 6100
rect 261159 6069 261171 6072
rect 261113 6063 261171 6069
rect 261662 6060 261668 6072
rect 261720 6060 261726 6112
rect 267642 6060 267648 6112
rect 267700 6100 267706 6112
rect 269684 6100 269712 6199
rect 270494 6196 270500 6248
rect 270552 6196 270558 6248
rect 267700 6072 269712 6100
rect 267700 6060 267706 6072
rect 270862 6060 270868 6112
rect 270920 6060 270926 6112
rect 1104 6010 271492 6032
rect 1104 5958 34748 6010
rect 34800 5958 34812 6010
rect 34864 5958 34876 6010
rect 34928 5958 34940 6010
rect 34992 5958 35004 6010
rect 35056 5958 102345 6010
rect 102397 5958 102409 6010
rect 102461 5958 102473 6010
rect 102525 5958 102537 6010
rect 102589 5958 102601 6010
rect 102653 5958 169942 6010
rect 169994 5958 170006 6010
rect 170058 5958 170070 6010
rect 170122 5958 170134 6010
rect 170186 5958 170198 6010
rect 170250 5958 237539 6010
rect 237591 5958 237603 6010
rect 237655 5958 237667 6010
rect 237719 5958 237731 6010
rect 237783 5958 237795 6010
rect 237847 5958 271492 6010
rect 1104 5936 271492 5958
rect 46658 5856 46664 5908
rect 46716 5856 46722 5908
rect 55766 5856 55772 5908
rect 55824 5896 55830 5908
rect 94498 5896 94504 5908
rect 55824 5868 94504 5896
rect 55824 5856 55830 5868
rect 94498 5856 94504 5868
rect 94556 5856 94562 5908
rect 95973 5899 96031 5905
rect 95973 5865 95985 5899
rect 96019 5896 96031 5899
rect 96062 5896 96068 5908
rect 96019 5868 96068 5896
rect 96019 5865 96031 5868
rect 95973 5859 96031 5865
rect 96062 5856 96068 5868
rect 96120 5856 96126 5908
rect 96154 5856 96160 5908
rect 96212 5856 96218 5908
rect 96430 5856 96436 5908
rect 96488 5896 96494 5908
rect 96709 5899 96767 5905
rect 96709 5896 96721 5899
rect 96488 5868 96721 5896
rect 96488 5856 96494 5868
rect 96709 5865 96721 5868
rect 96755 5865 96767 5899
rect 96709 5859 96767 5865
rect 97077 5899 97135 5905
rect 97077 5865 97089 5899
rect 97123 5896 97135 5899
rect 97123 5868 97672 5896
rect 97123 5865 97135 5868
rect 97077 5859 97135 5865
rect 97644 5840 97672 5868
rect 100110 5856 100116 5908
rect 100168 5856 100174 5908
rect 100938 5856 100944 5908
rect 100996 5896 101002 5908
rect 101766 5896 101772 5908
rect 100996 5868 101772 5896
rect 100996 5856 101002 5868
rect 101766 5856 101772 5868
rect 101824 5896 101830 5908
rect 101861 5899 101919 5905
rect 101861 5896 101873 5899
rect 101824 5868 101873 5896
rect 101824 5856 101830 5868
rect 101861 5865 101873 5868
rect 101907 5865 101919 5899
rect 101861 5859 101919 5865
rect 103422 5856 103428 5908
rect 103480 5896 103486 5908
rect 104345 5899 104403 5905
rect 104345 5896 104357 5899
rect 103480 5868 104357 5896
rect 103480 5856 103486 5868
rect 104345 5865 104357 5868
rect 104391 5865 104403 5899
rect 104345 5859 104403 5865
rect 106918 5856 106924 5908
rect 106976 5896 106982 5908
rect 107194 5896 107200 5908
rect 106976 5868 107200 5896
rect 106976 5856 106982 5868
rect 107194 5856 107200 5868
rect 107252 5856 107258 5908
rect 107286 5856 107292 5908
rect 107344 5896 107350 5908
rect 112162 5896 112168 5908
rect 107344 5868 112168 5896
rect 107344 5856 107350 5868
rect 112162 5856 112168 5868
rect 112220 5896 112226 5908
rect 112714 5896 112720 5908
rect 112220 5868 112720 5896
rect 112220 5856 112226 5868
rect 112714 5856 112720 5868
rect 112772 5856 112778 5908
rect 113453 5899 113511 5905
rect 113453 5896 113465 5899
rect 113008 5868 113465 5896
rect 77266 5800 86954 5828
rect 46474 5760 46480 5772
rect 46414 5732 46480 5760
rect 46474 5720 46480 5732
rect 46532 5760 46538 5772
rect 47581 5763 47639 5769
rect 47581 5760 47593 5763
rect 46532 5732 47593 5760
rect 46532 5720 46538 5732
rect 47581 5729 47593 5732
rect 47627 5729 47639 5763
rect 53098 5760 53104 5772
rect 53038 5732 53104 5760
rect 47581 5723 47639 5729
rect 53098 5720 53104 5732
rect 53156 5720 53162 5772
rect 45646 5652 45652 5704
rect 45704 5652 45710 5704
rect 46106 5652 46112 5704
rect 46164 5652 46170 5704
rect 46934 5652 46940 5704
rect 46992 5692 46998 5704
rect 47946 5692 47952 5704
rect 46992 5664 47952 5692
rect 46992 5652 46998 5664
rect 47946 5652 47952 5664
rect 48004 5692 48010 5704
rect 48133 5695 48191 5701
rect 48133 5692 48145 5695
rect 48004 5664 48145 5692
rect 48004 5652 48010 5664
rect 48133 5661 48145 5664
rect 48179 5661 48191 5695
rect 48133 5655 48191 5661
rect 51534 5652 51540 5704
rect 51592 5692 51598 5704
rect 51592 5664 52224 5692
rect 51592 5652 51598 5664
rect 35526 5584 35532 5636
rect 35584 5624 35590 5636
rect 35584 5596 45508 5624
rect 35584 5584 35590 5596
rect 45370 5516 45376 5568
rect 45428 5516 45434 5568
rect 45480 5556 45508 5596
rect 45738 5584 45744 5636
rect 45796 5584 45802 5636
rect 47210 5584 47216 5636
rect 47268 5624 47274 5636
rect 47305 5627 47363 5633
rect 47305 5624 47317 5627
rect 47268 5596 47317 5624
rect 47268 5584 47274 5596
rect 47305 5593 47317 5596
rect 47351 5593 47363 5627
rect 52196 5624 52224 5664
rect 52270 5652 52276 5704
rect 52328 5652 52334 5704
rect 52362 5652 52368 5704
rect 52420 5652 52426 5704
rect 55858 5652 55864 5704
rect 55916 5692 55922 5704
rect 77266 5692 77294 5800
rect 55916 5664 77294 5692
rect 86926 5692 86954 5800
rect 92658 5788 92664 5840
rect 92716 5828 92722 5840
rect 94038 5828 94044 5840
rect 92716 5800 94044 5828
rect 92716 5788 92722 5800
rect 94038 5788 94044 5800
rect 94096 5788 94102 5840
rect 95145 5831 95203 5837
rect 95145 5797 95157 5831
rect 95191 5828 95203 5831
rect 96614 5828 96620 5840
rect 95191 5800 96620 5828
rect 95191 5797 95203 5800
rect 95145 5791 95203 5797
rect 96614 5788 96620 5800
rect 96672 5788 96678 5840
rect 97626 5788 97632 5840
rect 97684 5788 97690 5840
rect 97902 5788 97908 5840
rect 97960 5828 97966 5840
rect 100389 5831 100447 5837
rect 100389 5828 100401 5831
rect 97960 5800 100401 5828
rect 97960 5788 97966 5800
rect 100389 5797 100401 5800
rect 100435 5797 100447 5831
rect 100389 5791 100447 5797
rect 101309 5831 101367 5837
rect 101309 5797 101321 5831
rect 101355 5828 101367 5831
rect 101674 5828 101680 5840
rect 101355 5800 101680 5828
rect 101355 5797 101367 5800
rect 101309 5791 101367 5797
rect 101674 5788 101680 5800
rect 101732 5788 101738 5840
rect 102229 5831 102287 5837
rect 102229 5797 102241 5831
rect 102275 5828 102287 5831
rect 102275 5800 102916 5828
rect 102275 5797 102287 5800
rect 102229 5791 102287 5797
rect 96982 5760 96988 5772
rect 95804 5732 96200 5760
rect 94590 5692 94596 5704
rect 86926 5664 94596 5692
rect 55916 5652 55922 5664
rect 94590 5652 94596 5664
rect 94648 5652 94654 5704
rect 94682 5652 94688 5704
rect 94740 5652 94746 5704
rect 95804 5701 95832 5732
rect 95329 5695 95387 5701
rect 95329 5661 95341 5695
rect 95375 5661 95387 5695
rect 95329 5655 95387 5661
rect 95789 5695 95847 5701
rect 95789 5661 95801 5695
rect 95835 5661 95847 5695
rect 95789 5655 95847 5661
rect 95973 5695 96031 5701
rect 95973 5661 95985 5695
rect 96019 5692 96031 5695
rect 96062 5692 96068 5704
rect 96019 5664 96068 5692
rect 96019 5661 96031 5664
rect 95973 5655 96031 5661
rect 52733 5627 52791 5633
rect 52733 5624 52745 5627
rect 52196 5596 52745 5624
rect 47305 5587 47363 5593
rect 52733 5593 52745 5596
rect 52779 5593 52791 5627
rect 52733 5587 52791 5593
rect 77478 5584 77484 5636
rect 77536 5624 77542 5636
rect 77536 5596 89714 5624
rect 77536 5584 77542 5596
rect 46477 5559 46535 5565
rect 46477 5556 46489 5559
rect 45480 5528 46489 5556
rect 46477 5525 46489 5528
rect 46523 5525 46535 5559
rect 46477 5519 46535 5525
rect 48314 5516 48320 5568
rect 48372 5516 48378 5568
rect 51169 5559 51227 5565
rect 51169 5525 51181 5559
rect 51215 5556 51227 5559
rect 51442 5556 51448 5568
rect 51215 5528 51448 5556
rect 51215 5525 51227 5528
rect 51169 5519 51227 5525
rect 51442 5516 51448 5528
rect 51500 5516 51506 5568
rect 51994 5516 52000 5568
rect 52052 5516 52058 5568
rect 52546 5516 52552 5568
rect 52604 5556 52610 5568
rect 53101 5559 53159 5565
rect 53101 5556 53113 5559
rect 52604 5528 53113 5556
rect 52604 5516 52610 5528
rect 53101 5525 53113 5528
rect 53147 5525 53159 5559
rect 53101 5519 53159 5525
rect 53282 5516 53288 5568
rect 53340 5516 53346 5568
rect 89686 5556 89714 5596
rect 92382 5584 92388 5636
rect 92440 5624 92446 5636
rect 95234 5624 95240 5636
rect 92440 5596 95240 5624
rect 92440 5584 92446 5596
rect 95234 5584 95240 5596
rect 95292 5584 95298 5636
rect 95344 5624 95372 5655
rect 96062 5652 96068 5664
rect 96120 5652 96126 5704
rect 96172 5692 96200 5732
rect 96724 5732 96988 5760
rect 96724 5701 96752 5732
rect 96982 5720 96988 5732
rect 97040 5720 97046 5772
rect 97074 5720 97080 5772
rect 97132 5760 97138 5772
rect 97537 5763 97595 5769
rect 97537 5760 97549 5763
rect 97132 5732 97549 5760
rect 97132 5720 97138 5732
rect 97537 5729 97549 5732
rect 97583 5729 97595 5763
rect 97537 5723 97595 5729
rect 97718 5720 97724 5772
rect 97776 5720 97782 5772
rect 98454 5720 98460 5772
rect 98512 5720 98518 5772
rect 98546 5720 98552 5772
rect 98604 5760 98610 5772
rect 101033 5763 101091 5769
rect 101033 5760 101045 5763
rect 98604 5732 101045 5760
rect 98604 5720 98610 5732
rect 101033 5729 101045 5732
rect 101079 5760 101091 5763
rect 101490 5760 101496 5772
rect 101079 5732 101496 5760
rect 101079 5729 101091 5732
rect 101033 5723 101091 5729
rect 101490 5720 101496 5732
rect 101548 5760 101554 5772
rect 101953 5763 102011 5769
rect 101953 5760 101965 5763
rect 101548 5732 101965 5760
rect 101548 5720 101554 5732
rect 101953 5729 101965 5732
rect 101999 5760 102011 5763
rect 102410 5760 102416 5772
rect 101999 5732 102416 5760
rect 101999 5729 102011 5732
rect 101953 5723 102011 5729
rect 102410 5720 102416 5732
rect 102468 5720 102474 5772
rect 102888 5760 102916 5800
rect 102962 5788 102968 5840
rect 103020 5828 103026 5840
rect 104526 5828 104532 5840
rect 103020 5800 104532 5828
rect 103020 5788 103026 5800
rect 104526 5788 104532 5800
rect 104584 5788 104590 5840
rect 104894 5788 104900 5840
rect 104952 5828 104958 5840
rect 107657 5831 107715 5837
rect 107657 5828 107669 5831
rect 104952 5800 107669 5828
rect 104952 5788 104958 5800
rect 107657 5797 107669 5800
rect 107703 5797 107715 5831
rect 107657 5791 107715 5797
rect 108206 5788 108212 5840
rect 108264 5828 108270 5840
rect 108393 5831 108451 5837
rect 108393 5828 108405 5831
rect 108264 5800 108405 5828
rect 108264 5788 108270 5800
rect 108393 5797 108405 5800
rect 108439 5797 108451 5831
rect 108393 5791 108451 5797
rect 108758 5788 108764 5840
rect 108816 5828 108822 5840
rect 108816 5800 109908 5828
rect 108816 5788 108822 5800
rect 108942 5760 108948 5772
rect 102888 5732 103652 5760
rect 96709 5695 96767 5701
rect 96709 5692 96721 5695
rect 96172 5664 96721 5692
rect 96709 5661 96721 5664
rect 96755 5692 96767 5695
rect 96798 5692 96804 5704
rect 96755 5664 96804 5692
rect 96755 5661 96767 5664
rect 96709 5655 96767 5661
rect 96798 5652 96804 5664
rect 96856 5652 96862 5704
rect 96893 5695 96951 5701
rect 96893 5661 96905 5695
rect 96939 5692 96951 5695
rect 97350 5692 97356 5704
rect 96939 5664 97356 5692
rect 96939 5661 96951 5664
rect 96893 5655 96951 5661
rect 97350 5652 97356 5664
rect 97408 5652 97414 5704
rect 99374 5652 99380 5704
rect 99432 5692 99438 5704
rect 99558 5692 99564 5704
rect 99432 5664 99564 5692
rect 99432 5652 99438 5664
rect 99558 5652 99564 5664
rect 99616 5692 99622 5704
rect 99837 5695 99895 5701
rect 99837 5692 99849 5695
rect 99616 5664 99849 5692
rect 99616 5652 99622 5664
rect 99837 5661 99849 5664
rect 99883 5661 99895 5695
rect 99837 5655 99895 5661
rect 100205 5695 100263 5701
rect 100205 5661 100217 5695
rect 100251 5692 100263 5695
rect 100386 5692 100392 5704
rect 100251 5664 100392 5692
rect 100251 5661 100263 5664
rect 100205 5655 100263 5661
rect 98638 5624 98644 5636
rect 95344 5596 98644 5624
rect 98638 5584 98644 5596
rect 98696 5584 98702 5636
rect 99852 5624 99880 5655
rect 100386 5652 100392 5664
rect 100444 5652 100450 5704
rect 100938 5652 100944 5704
rect 100996 5692 101002 5704
rect 101861 5695 101919 5701
rect 101861 5692 101873 5695
rect 100996 5664 101873 5692
rect 100996 5652 101002 5664
rect 101861 5661 101873 5664
rect 101907 5692 101919 5695
rect 102318 5692 102324 5704
rect 101907 5664 102324 5692
rect 101907 5661 101919 5664
rect 101861 5655 101919 5661
rect 102318 5652 102324 5664
rect 102376 5692 102382 5704
rect 102962 5692 102968 5704
rect 102376 5664 102968 5692
rect 102376 5652 102382 5664
rect 102962 5652 102968 5664
rect 103020 5652 103026 5704
rect 103624 5701 103652 5732
rect 106476 5732 108948 5760
rect 103609 5695 103667 5701
rect 103609 5661 103621 5695
rect 103655 5661 103667 5695
rect 103609 5655 103667 5661
rect 104526 5652 104532 5704
rect 104584 5652 104590 5704
rect 105173 5695 105231 5701
rect 105173 5661 105185 5695
rect 105219 5692 105231 5695
rect 105262 5692 105268 5704
rect 105219 5664 105268 5692
rect 105219 5661 105231 5664
rect 105173 5655 105231 5661
rect 105262 5652 105268 5664
rect 105320 5652 105326 5704
rect 105817 5695 105875 5701
rect 105817 5661 105829 5695
rect 105863 5692 105875 5695
rect 106366 5692 106372 5704
rect 105863 5664 106372 5692
rect 105863 5661 105875 5664
rect 105817 5655 105875 5661
rect 106366 5652 106372 5664
rect 106424 5652 106430 5704
rect 106476 5701 106504 5732
rect 108942 5720 108948 5732
rect 109000 5720 109006 5772
rect 109034 5720 109040 5772
rect 109092 5720 109098 5772
rect 109218 5720 109224 5772
rect 109276 5720 109282 5772
rect 109880 5760 109908 5800
rect 109954 5788 109960 5840
rect 110012 5828 110018 5840
rect 112441 5831 112499 5837
rect 112441 5828 112453 5831
rect 110012 5800 112453 5828
rect 110012 5788 110018 5800
rect 112441 5797 112453 5800
rect 112487 5828 112499 5831
rect 112898 5828 112904 5840
rect 112487 5800 112904 5828
rect 112487 5797 112499 5800
rect 112441 5791 112499 5797
rect 112898 5788 112904 5800
rect 112956 5788 112962 5840
rect 113008 5760 113036 5868
rect 113376 5840 113404 5868
rect 113453 5865 113465 5868
rect 113499 5896 113511 5899
rect 114281 5899 114339 5905
rect 114281 5896 114293 5899
rect 113499 5868 114293 5896
rect 113499 5865 113511 5868
rect 113453 5859 113511 5865
rect 114281 5865 114293 5868
rect 114327 5865 114339 5899
rect 114281 5859 114339 5865
rect 114830 5856 114836 5908
rect 114888 5896 114894 5908
rect 116026 5896 116032 5908
rect 114888 5868 116032 5896
rect 114888 5856 114894 5868
rect 116026 5856 116032 5868
rect 116084 5856 116090 5908
rect 116578 5856 116584 5908
rect 116636 5856 116642 5908
rect 116762 5856 116768 5908
rect 116820 5856 116826 5908
rect 148318 5896 148324 5908
rect 116872 5868 148324 5896
rect 113358 5788 113364 5840
rect 113416 5788 113422 5840
rect 113473 5800 113680 5828
rect 113473 5760 113501 5800
rect 109880 5732 113036 5760
rect 113100 5732 113501 5760
rect 113652 5760 113680 5800
rect 114646 5788 114652 5840
rect 114704 5788 114710 5840
rect 114738 5788 114744 5840
rect 114796 5828 114802 5840
rect 116872 5828 116900 5868
rect 148318 5856 148324 5868
rect 148376 5856 148382 5908
rect 149790 5856 149796 5908
rect 149848 5896 149854 5908
rect 150069 5899 150127 5905
rect 150069 5896 150081 5899
rect 149848 5868 150081 5896
rect 149848 5856 149854 5868
rect 150069 5865 150081 5868
rect 150115 5865 150127 5899
rect 154850 5896 154856 5908
rect 150069 5859 150127 5865
rect 150360 5868 154856 5896
rect 114796 5800 116900 5828
rect 116964 5800 121592 5828
rect 114796 5788 114802 5800
rect 113726 5760 113732 5772
rect 113652 5732 113732 5760
rect 106461 5695 106519 5701
rect 106461 5661 106473 5695
rect 106507 5661 106519 5695
rect 106461 5655 106519 5661
rect 107105 5695 107163 5701
rect 107105 5661 107117 5695
rect 107151 5692 107163 5695
rect 107194 5692 107200 5704
rect 107151 5664 107200 5692
rect 107151 5661 107163 5664
rect 107105 5655 107163 5661
rect 107194 5652 107200 5664
rect 107252 5652 107258 5704
rect 107378 5652 107384 5704
rect 107436 5652 107442 5704
rect 110414 5652 110420 5704
rect 110472 5692 110478 5704
rect 110472 5664 111472 5692
rect 110472 5652 110478 5664
rect 111444 5636 111472 5664
rect 112162 5652 112168 5704
rect 112220 5692 112226 5704
rect 112257 5695 112315 5701
rect 112257 5692 112269 5695
rect 112220 5664 112269 5692
rect 112220 5652 112226 5664
rect 112257 5661 112269 5664
rect 112303 5661 112315 5695
rect 113100 5692 113128 5732
rect 113726 5720 113732 5732
rect 113784 5760 113790 5772
rect 114373 5763 114431 5769
rect 114373 5760 114385 5763
rect 113784 5732 114385 5760
rect 113784 5720 113790 5732
rect 114373 5729 114385 5732
rect 114419 5729 114431 5763
rect 114373 5723 114431 5729
rect 115198 5720 115204 5772
rect 115256 5760 115262 5772
rect 115385 5763 115443 5769
rect 115385 5760 115397 5763
rect 115256 5732 115397 5760
rect 115256 5720 115262 5732
rect 115385 5729 115397 5732
rect 115431 5729 115443 5763
rect 115385 5723 115443 5729
rect 115569 5763 115627 5769
rect 115569 5729 115581 5763
rect 115615 5760 115627 5763
rect 115750 5760 115756 5772
rect 115615 5732 115756 5760
rect 115615 5729 115627 5732
rect 115569 5723 115627 5729
rect 115750 5720 115756 5732
rect 115808 5720 115814 5772
rect 116486 5720 116492 5772
rect 116544 5720 116550 5772
rect 112257 5655 112315 5661
rect 112364 5664 113128 5692
rect 113453 5695 113511 5701
rect 100294 5624 100300 5636
rect 99852 5596 100300 5624
rect 100294 5584 100300 5596
rect 100352 5584 100358 5636
rect 100662 5584 100668 5636
rect 100720 5624 100726 5636
rect 101950 5624 101956 5636
rect 100720 5596 101956 5624
rect 100720 5584 100726 5596
rect 101950 5584 101956 5596
rect 102008 5584 102014 5636
rect 102781 5627 102839 5633
rect 102781 5593 102793 5627
rect 102827 5624 102839 5627
rect 107286 5624 107292 5636
rect 102827 5596 107292 5624
rect 102827 5593 102839 5596
rect 102781 5587 102839 5593
rect 94406 5556 94412 5568
rect 89686 5528 94412 5556
rect 94406 5516 94412 5528
rect 94464 5516 94470 5568
rect 94501 5559 94559 5565
rect 94501 5525 94513 5559
rect 94547 5556 94559 5559
rect 96154 5556 96160 5568
rect 94547 5528 96160 5556
rect 94547 5525 94559 5528
rect 94501 5519 94559 5525
rect 96154 5516 96160 5528
rect 96212 5516 96218 5568
rect 96430 5516 96436 5568
rect 96488 5556 96494 5568
rect 97442 5556 97448 5568
rect 96488 5528 97448 5556
rect 96488 5516 96494 5528
rect 97442 5516 97448 5528
rect 97500 5516 97506 5568
rect 99006 5516 99012 5568
rect 99064 5556 99070 5568
rect 100018 5556 100024 5568
rect 99064 5528 100024 5556
rect 99064 5516 99070 5528
rect 100018 5516 100024 5528
rect 100076 5516 100082 5568
rect 100110 5516 100116 5568
rect 100168 5556 100174 5568
rect 102796 5556 102824 5587
rect 107286 5584 107292 5596
rect 107344 5584 107350 5636
rect 107654 5584 107660 5636
rect 107712 5624 107718 5636
rect 108209 5627 108267 5633
rect 108209 5624 108221 5627
rect 107712 5596 108221 5624
rect 107712 5584 107718 5596
rect 108209 5593 108221 5596
rect 108255 5624 108267 5627
rect 110230 5624 110236 5636
rect 108255 5596 110236 5624
rect 108255 5593 108267 5596
rect 108209 5587 108267 5593
rect 110230 5584 110236 5596
rect 110288 5584 110294 5636
rect 110874 5584 110880 5636
rect 110932 5584 110938 5636
rect 111426 5584 111432 5636
rect 111484 5584 111490 5636
rect 112364 5624 112392 5664
rect 113453 5661 113465 5695
rect 113499 5661 113511 5695
rect 113453 5655 113511 5661
rect 113637 5695 113695 5701
rect 113637 5661 113649 5695
rect 113683 5692 113695 5695
rect 113744 5692 113772 5720
rect 113683 5664 113772 5692
rect 113683 5661 113695 5664
rect 113637 5655 113695 5661
rect 111536 5596 112392 5624
rect 100168 5528 102824 5556
rect 100168 5516 100174 5528
rect 102962 5516 102968 5568
rect 103020 5556 103026 5568
rect 103425 5559 103483 5565
rect 103425 5556 103437 5559
rect 103020 5528 103437 5556
rect 103020 5516 103026 5528
rect 103425 5525 103437 5528
rect 103471 5525 103483 5559
rect 103425 5519 103483 5525
rect 104802 5516 104808 5568
rect 104860 5556 104866 5568
rect 104989 5559 105047 5565
rect 104989 5556 105001 5559
rect 104860 5528 105001 5556
rect 104860 5516 104866 5528
rect 104989 5525 105001 5528
rect 105035 5525 105047 5559
rect 104989 5519 105047 5525
rect 105446 5516 105452 5568
rect 105504 5556 105510 5568
rect 105633 5559 105691 5565
rect 105633 5556 105645 5559
rect 105504 5528 105645 5556
rect 105504 5516 105510 5528
rect 105633 5525 105645 5528
rect 105679 5525 105691 5559
rect 105633 5519 105691 5525
rect 106277 5559 106335 5565
rect 106277 5525 106289 5559
rect 106323 5556 106335 5559
rect 108114 5556 108120 5568
rect 106323 5528 108120 5556
rect 106323 5525 106335 5528
rect 106277 5519 106335 5525
rect 108114 5516 108120 5528
rect 108172 5516 108178 5568
rect 108666 5516 108672 5568
rect 108724 5556 108730 5568
rect 111536 5565 111564 5596
rect 113468 5595 113496 5655
rect 114186 5652 114192 5704
rect 114244 5692 114250 5704
rect 114281 5695 114339 5701
rect 114281 5692 114293 5695
rect 114244 5664 114293 5692
rect 114244 5652 114250 5664
rect 114281 5661 114293 5664
rect 114327 5661 114339 5695
rect 114281 5655 114339 5661
rect 115106 5652 115112 5704
rect 115164 5652 115170 5704
rect 115477 5695 115535 5701
rect 115477 5661 115489 5695
rect 115523 5692 115535 5695
rect 115658 5692 115664 5704
rect 115523 5664 115664 5692
rect 115523 5661 115535 5664
rect 115477 5655 115535 5661
rect 115658 5652 115664 5664
rect 115716 5652 115722 5704
rect 116394 5652 116400 5704
rect 116452 5652 116458 5704
rect 114204 5624 114232 5652
rect 113560 5596 114232 5624
rect 113560 5595 113588 5596
rect 113468 5567 113588 5595
rect 114462 5584 114468 5636
rect 114520 5624 114526 5636
rect 116964 5624 116992 5800
rect 117314 5720 117320 5772
rect 117372 5720 117378 5772
rect 117590 5720 117596 5772
rect 117648 5760 117654 5772
rect 119062 5760 119068 5772
rect 117648 5732 119068 5760
rect 117648 5720 117654 5732
rect 119062 5720 119068 5732
rect 119120 5720 119126 5772
rect 120102 5763 120160 5769
rect 120102 5760 120114 5763
rect 119356 5732 120114 5760
rect 119157 5695 119215 5701
rect 119157 5661 119169 5695
rect 119203 5692 119215 5695
rect 119246 5692 119252 5704
rect 119203 5664 119252 5692
rect 119203 5661 119215 5664
rect 119157 5655 119215 5661
rect 119246 5652 119252 5664
rect 119304 5652 119310 5704
rect 114520 5596 116992 5624
rect 114520 5584 114526 5596
rect 117498 5584 117504 5636
rect 117556 5584 117562 5636
rect 118234 5584 118240 5636
rect 118292 5624 118298 5636
rect 119356 5624 119384 5732
rect 120102 5729 120114 5732
rect 120148 5729 120160 5763
rect 121454 5760 121460 5772
rect 120102 5723 120160 5729
rect 120276 5732 121460 5760
rect 119617 5695 119675 5701
rect 119617 5661 119629 5695
rect 119663 5692 119675 5695
rect 119663 5688 120212 5692
rect 120276 5688 120304 5732
rect 121454 5720 121460 5732
rect 121512 5720 121518 5772
rect 121564 5760 121592 5800
rect 121638 5788 121644 5840
rect 121696 5828 121702 5840
rect 135530 5828 135536 5840
rect 121696 5800 135536 5828
rect 121696 5788 121702 5800
rect 135530 5788 135536 5800
rect 135588 5788 135594 5840
rect 138937 5831 138995 5837
rect 135916 5800 138796 5828
rect 135916 5760 135944 5800
rect 138768 5772 138796 5800
rect 138937 5797 138949 5831
rect 138983 5828 138995 5831
rect 138983 5800 140176 5828
rect 138983 5797 138995 5800
rect 138937 5791 138995 5797
rect 137186 5760 137192 5772
rect 121564 5732 135944 5760
rect 136008 5732 137192 5760
rect 121564 5701 121592 5732
rect 120997 5695 121055 5701
rect 120997 5692 121009 5695
rect 119663 5664 120304 5688
rect 119663 5661 119675 5664
rect 119617 5655 119675 5661
rect 120184 5660 120304 5664
rect 120644 5664 121009 5692
rect 118292 5596 119384 5624
rect 118292 5584 118298 5596
rect 111521 5559 111579 5565
rect 111521 5556 111533 5559
rect 108724 5528 111533 5556
rect 108724 5516 108730 5528
rect 111521 5525 111533 5528
rect 111567 5525 111579 5559
rect 111521 5519 111579 5525
rect 113634 5516 113640 5568
rect 113692 5556 113698 5568
rect 113821 5559 113879 5565
rect 113821 5556 113833 5559
rect 113692 5528 113833 5556
rect 113692 5516 113698 5528
rect 113821 5525 113833 5528
rect 113867 5525 113879 5559
rect 113821 5519 113879 5525
rect 114002 5516 114008 5568
rect 114060 5556 114066 5568
rect 115753 5559 115811 5565
rect 115753 5556 115765 5559
rect 114060 5528 115765 5556
rect 114060 5516 114066 5528
rect 115753 5525 115765 5528
rect 115799 5525 115811 5559
rect 115753 5519 115811 5525
rect 116026 5516 116032 5568
rect 116084 5556 116090 5568
rect 117590 5556 117596 5568
rect 116084 5528 117596 5556
rect 116084 5516 116090 5528
rect 117590 5516 117596 5528
rect 117648 5516 117654 5568
rect 118694 5516 118700 5568
rect 118752 5556 118758 5568
rect 119632 5556 119660 5655
rect 119890 5584 119896 5636
rect 119948 5584 119954 5636
rect 119985 5627 120043 5633
rect 119985 5593 119997 5627
rect 120031 5624 120043 5627
rect 120534 5624 120540 5636
rect 120031 5596 120540 5624
rect 120031 5593 120043 5596
rect 119985 5587 120043 5593
rect 120534 5584 120540 5596
rect 120592 5584 120598 5636
rect 118752 5528 119660 5556
rect 120261 5559 120319 5565
rect 118752 5516 118758 5528
rect 120261 5525 120273 5559
rect 120307 5556 120319 5559
rect 120644 5556 120672 5664
rect 120997 5661 121009 5664
rect 121043 5661 121055 5695
rect 120997 5655 121055 5661
rect 121549 5695 121607 5701
rect 121549 5661 121561 5695
rect 121595 5661 121607 5695
rect 121549 5655 121607 5661
rect 121914 5652 121920 5704
rect 121972 5652 121978 5704
rect 127710 5652 127716 5704
rect 127768 5652 127774 5704
rect 128078 5652 128084 5704
rect 128136 5652 128142 5704
rect 136008 5692 136036 5732
rect 137186 5720 137192 5732
rect 137244 5720 137250 5772
rect 138750 5720 138756 5772
rect 138808 5760 138814 5772
rect 140038 5760 140044 5772
rect 138808 5732 140044 5760
rect 138808 5720 138814 5732
rect 140038 5720 140044 5732
rect 140096 5720 140102 5772
rect 140148 5760 140176 5800
rect 140682 5788 140688 5840
rect 140740 5828 140746 5840
rect 148781 5831 148839 5837
rect 140740 5800 145512 5828
rect 140740 5788 140746 5800
rect 140777 5763 140835 5769
rect 140777 5760 140789 5763
rect 140148 5732 140789 5760
rect 140777 5729 140789 5732
rect 140823 5729 140835 5763
rect 145098 5760 145104 5772
rect 140777 5723 140835 5729
rect 142356 5732 145104 5760
rect 128326 5664 136036 5692
rect 120718 5584 120724 5636
rect 120776 5624 120782 5636
rect 128326 5624 128354 5664
rect 136082 5652 136088 5704
rect 136140 5652 136146 5704
rect 138106 5652 138112 5704
rect 138164 5692 138170 5704
rect 139121 5695 139179 5701
rect 139121 5692 139133 5695
rect 138164 5664 139133 5692
rect 138164 5652 138170 5664
rect 139121 5661 139133 5664
rect 139167 5661 139179 5695
rect 139121 5655 139179 5661
rect 139762 5652 139768 5704
rect 139820 5652 139826 5704
rect 140593 5695 140651 5701
rect 140593 5661 140605 5695
rect 140639 5661 140651 5695
rect 140593 5655 140651 5661
rect 120776 5596 128354 5624
rect 120776 5584 120782 5596
rect 132862 5584 132868 5636
rect 132920 5584 132926 5636
rect 133230 5584 133236 5636
rect 133288 5624 133294 5636
rect 136100 5624 136128 5652
rect 133288 5596 136128 5624
rect 140608 5624 140636 5655
rect 142356 5624 142384 5732
rect 145098 5720 145104 5732
rect 145156 5720 145162 5772
rect 145484 5760 145512 5800
rect 148781 5797 148793 5831
rect 148827 5828 148839 5831
rect 150360 5828 150388 5868
rect 154850 5856 154856 5868
rect 154908 5856 154914 5908
rect 155957 5899 156015 5905
rect 155957 5865 155969 5899
rect 156003 5896 156015 5899
rect 156414 5896 156420 5908
rect 156003 5868 156420 5896
rect 156003 5865 156015 5868
rect 155957 5859 156015 5865
rect 156414 5856 156420 5868
rect 156472 5856 156478 5908
rect 157702 5856 157708 5908
rect 157760 5856 157766 5908
rect 162118 5856 162124 5908
rect 162176 5896 162182 5908
rect 169205 5899 169263 5905
rect 169205 5896 169217 5899
rect 162176 5868 169217 5896
rect 162176 5856 162182 5868
rect 169205 5865 169217 5868
rect 169251 5896 169263 5899
rect 169251 5868 195974 5896
rect 169251 5865 169263 5868
rect 169205 5859 169263 5865
rect 148827 5800 150388 5828
rect 150529 5831 150587 5837
rect 148827 5797 148839 5800
rect 148781 5791 148839 5797
rect 150529 5797 150541 5831
rect 150575 5828 150587 5831
rect 154482 5828 154488 5840
rect 150575 5800 151768 5828
rect 150575 5797 150587 5800
rect 150529 5791 150587 5797
rect 147122 5760 147128 5772
rect 145484 5732 147128 5760
rect 142430 5652 142436 5704
rect 142488 5652 142494 5704
rect 143258 5652 143264 5704
rect 143316 5652 143322 5704
rect 143534 5652 143540 5704
rect 143592 5692 143598 5704
rect 144822 5692 144828 5704
rect 143592 5664 144828 5692
rect 143592 5652 143598 5664
rect 144822 5652 144828 5664
rect 144880 5652 144886 5704
rect 145484 5701 145512 5732
rect 147122 5720 147128 5732
rect 147180 5720 147186 5772
rect 148502 5720 148508 5772
rect 148560 5720 148566 5772
rect 151262 5760 151268 5772
rect 149532 5732 151268 5760
rect 145469 5695 145527 5701
rect 145469 5661 145481 5695
rect 145515 5661 145527 5695
rect 146481 5695 146539 5701
rect 146481 5692 146493 5695
rect 145469 5655 145527 5661
rect 145852 5664 146493 5692
rect 144089 5627 144147 5633
rect 144089 5624 144101 5627
rect 140608 5596 142384 5624
rect 142540 5596 144101 5624
rect 133288 5584 133294 5596
rect 120307 5528 120672 5556
rect 120813 5559 120871 5565
rect 120307 5525 120319 5528
rect 120261 5519 120319 5525
rect 120813 5525 120825 5559
rect 120859 5556 120871 5559
rect 121178 5556 121184 5568
rect 120859 5528 121184 5556
rect 120859 5525 120871 5528
rect 120813 5519 120871 5525
rect 121178 5516 121184 5528
rect 121236 5516 121242 5568
rect 135898 5516 135904 5568
rect 135956 5556 135962 5568
rect 136269 5559 136327 5565
rect 136269 5556 136281 5559
rect 135956 5528 136281 5556
rect 135956 5516 135962 5528
rect 136269 5525 136281 5528
rect 136315 5525 136327 5559
rect 136269 5519 136327 5525
rect 140314 5516 140320 5568
rect 140372 5556 140378 5568
rect 142540 5556 142568 5596
rect 144089 5593 144101 5596
rect 144135 5593 144147 5627
rect 144089 5587 144147 5593
rect 140372 5528 142568 5556
rect 143077 5559 143135 5565
rect 140372 5516 140378 5528
rect 143077 5525 143089 5559
rect 143123 5556 143135 5559
rect 143350 5556 143356 5568
rect 143123 5528 143356 5556
rect 143123 5525 143135 5528
rect 143077 5519 143135 5525
rect 143350 5516 143356 5528
rect 143408 5516 143414 5568
rect 144104 5556 144132 5587
rect 145558 5584 145564 5636
rect 145616 5624 145622 5636
rect 145745 5627 145803 5633
rect 145745 5624 145757 5627
rect 145616 5596 145757 5624
rect 145616 5584 145622 5596
rect 145745 5593 145757 5596
rect 145791 5593 145803 5627
rect 145745 5587 145803 5593
rect 145852 5556 145880 5664
rect 146481 5661 146493 5664
rect 146527 5661 146539 5695
rect 146481 5655 146539 5661
rect 146757 5695 146815 5701
rect 146757 5661 146769 5695
rect 146803 5692 146815 5695
rect 147950 5692 147956 5704
rect 146803 5664 147956 5692
rect 146803 5661 146815 5664
rect 146757 5655 146815 5661
rect 147950 5652 147956 5664
rect 148008 5652 148014 5704
rect 148134 5652 148140 5704
rect 148192 5692 148198 5704
rect 149532 5701 149560 5732
rect 151262 5720 151268 5732
rect 151320 5720 151326 5772
rect 151354 5720 151360 5772
rect 151412 5760 151418 5772
rect 151630 5760 151636 5772
rect 151412 5732 151636 5760
rect 151412 5720 151418 5732
rect 151630 5720 151636 5732
rect 151688 5720 151694 5772
rect 151740 5760 151768 5800
rect 153212 5800 154488 5828
rect 153212 5760 153240 5800
rect 154482 5788 154488 5800
rect 154540 5788 154546 5840
rect 188798 5788 188804 5840
rect 188856 5788 188862 5840
rect 190089 5831 190147 5837
rect 190089 5797 190101 5831
rect 190135 5828 190147 5831
rect 190454 5828 190460 5840
rect 190135 5800 190460 5828
rect 190135 5797 190147 5800
rect 190089 5791 190147 5797
rect 190454 5788 190460 5800
rect 190512 5788 190518 5840
rect 195946 5828 195974 5868
rect 210418 5856 210424 5908
rect 210476 5896 210482 5908
rect 216674 5896 216680 5908
rect 210476 5868 216680 5896
rect 210476 5856 210482 5868
rect 216674 5856 216680 5868
rect 216732 5856 216738 5908
rect 217413 5899 217471 5905
rect 217413 5865 217425 5899
rect 217459 5896 217471 5899
rect 217962 5896 217968 5908
rect 217459 5868 217968 5896
rect 217459 5865 217471 5868
rect 217413 5859 217471 5865
rect 217962 5856 217968 5868
rect 218020 5856 218026 5908
rect 218422 5856 218428 5908
rect 218480 5896 218486 5908
rect 218790 5896 218796 5908
rect 218480 5868 218796 5896
rect 218480 5856 218486 5868
rect 218790 5856 218796 5868
rect 218848 5856 218854 5908
rect 218974 5856 218980 5908
rect 219032 5896 219038 5908
rect 222654 5896 222660 5908
rect 219032 5868 222660 5896
rect 219032 5856 219038 5868
rect 222654 5856 222660 5868
rect 222712 5856 222718 5908
rect 222746 5856 222752 5908
rect 222804 5896 222810 5908
rect 224957 5899 225015 5905
rect 224957 5896 224969 5899
rect 222804 5868 224969 5896
rect 222804 5856 222810 5868
rect 224957 5865 224969 5868
rect 225003 5865 225015 5899
rect 224957 5859 225015 5865
rect 225046 5856 225052 5908
rect 225104 5896 225110 5908
rect 225693 5899 225751 5905
rect 225693 5896 225705 5899
rect 225104 5868 225705 5896
rect 225104 5856 225110 5868
rect 225693 5865 225705 5868
rect 225739 5865 225751 5899
rect 225693 5859 225751 5865
rect 226886 5856 226892 5908
rect 226944 5896 226950 5908
rect 245562 5896 245568 5908
rect 226944 5868 245568 5896
rect 226944 5856 226950 5868
rect 245562 5856 245568 5868
rect 245620 5856 245626 5908
rect 248046 5856 248052 5908
rect 248104 5856 248110 5908
rect 248230 5856 248236 5908
rect 248288 5856 248294 5908
rect 248782 5856 248788 5908
rect 248840 5896 248846 5908
rect 248877 5899 248935 5905
rect 248877 5896 248889 5899
rect 248840 5868 248889 5896
rect 248840 5856 248846 5868
rect 248877 5865 248889 5868
rect 248923 5896 248935 5899
rect 249705 5899 249763 5905
rect 249705 5896 249717 5899
rect 248923 5868 249717 5896
rect 248923 5865 248935 5868
rect 248877 5859 248935 5865
rect 249705 5865 249717 5868
rect 249751 5896 249763 5899
rect 251726 5896 251732 5908
rect 249751 5868 251732 5896
rect 249751 5865 249763 5868
rect 249705 5859 249763 5865
rect 251726 5856 251732 5868
rect 251784 5856 251790 5908
rect 256326 5896 256332 5908
rect 253906 5868 256332 5896
rect 213362 5828 213368 5840
rect 195946 5800 213368 5828
rect 213362 5788 213368 5800
rect 213420 5788 213426 5840
rect 213454 5788 213460 5840
rect 213512 5828 213518 5840
rect 223206 5828 223212 5840
rect 213512 5800 223212 5828
rect 213512 5788 213518 5800
rect 223206 5788 223212 5800
rect 223264 5788 223270 5840
rect 223298 5788 223304 5840
rect 223356 5788 223362 5840
rect 224770 5788 224776 5840
rect 224828 5828 224834 5840
rect 224828 5800 226196 5828
rect 224828 5788 224834 5800
rect 151740 5732 153240 5760
rect 153286 5720 153292 5772
rect 153344 5760 153350 5772
rect 153749 5763 153807 5769
rect 153749 5760 153761 5763
rect 153344 5732 153761 5760
rect 153344 5720 153350 5732
rect 153749 5729 153761 5732
rect 153795 5729 153807 5763
rect 153749 5723 153807 5729
rect 153838 5720 153844 5772
rect 153896 5760 153902 5772
rect 154393 5763 154451 5769
rect 154393 5760 154405 5763
rect 153896 5732 154405 5760
rect 153896 5720 153902 5732
rect 154393 5729 154405 5732
rect 154439 5729 154451 5763
rect 154393 5723 154451 5729
rect 154666 5720 154672 5772
rect 154724 5720 154730 5772
rect 154807 5763 154865 5769
rect 154807 5729 154819 5763
rect 154853 5760 154865 5763
rect 155862 5760 155868 5772
rect 154853 5732 155868 5760
rect 154853 5729 154865 5732
rect 154807 5723 154865 5729
rect 155862 5720 155868 5732
rect 155920 5720 155926 5772
rect 158806 5760 158812 5772
rect 157458 5732 158812 5760
rect 158806 5720 158812 5732
rect 158864 5720 158870 5772
rect 169662 5760 169668 5772
rect 166966 5732 169668 5760
rect 148229 5695 148287 5701
rect 148229 5692 148241 5695
rect 148192 5664 148241 5692
rect 148192 5652 148198 5664
rect 148229 5661 148241 5664
rect 148275 5661 148287 5695
rect 148229 5655 148287 5661
rect 149517 5695 149575 5701
rect 149517 5661 149529 5695
rect 149563 5661 149575 5695
rect 149977 5695 150035 5701
rect 149977 5692 149989 5695
rect 149517 5655 149575 5661
rect 149716 5664 149989 5692
rect 147968 5624 147996 5652
rect 149716 5636 149744 5664
rect 149977 5661 149989 5664
rect 150023 5661 150035 5695
rect 149977 5655 150035 5661
rect 150250 5652 150256 5704
rect 150308 5652 150314 5704
rect 150342 5652 150348 5704
rect 150400 5692 150406 5704
rect 150989 5695 151047 5701
rect 150989 5692 151001 5695
rect 150400 5664 151001 5692
rect 150400 5652 150406 5664
rect 150989 5661 151001 5664
rect 151035 5661 151047 5695
rect 150989 5655 151047 5661
rect 151170 5652 151176 5704
rect 151228 5652 151234 5704
rect 151906 5652 151912 5704
rect 151964 5652 151970 5704
rect 152090 5701 152096 5704
rect 152047 5695 152096 5701
rect 152047 5661 152059 5695
rect 152093 5661 152096 5695
rect 152047 5655 152096 5661
rect 152090 5652 152096 5655
rect 152148 5652 152154 5704
rect 152182 5652 152188 5704
rect 152240 5652 152246 5704
rect 153933 5695 153991 5701
rect 153933 5661 153945 5695
rect 153979 5661 153991 5695
rect 153933 5655 153991 5661
rect 149698 5624 149704 5636
rect 147968 5596 149704 5624
rect 149698 5584 149704 5596
rect 149756 5584 149762 5636
rect 149790 5584 149796 5636
rect 149848 5624 149854 5636
rect 150894 5624 150900 5636
rect 149848 5596 150900 5624
rect 149848 5584 149854 5596
rect 150894 5584 150900 5596
rect 150952 5584 150958 5636
rect 144104 5528 145880 5556
rect 149333 5559 149391 5565
rect 149333 5525 149345 5559
rect 149379 5556 149391 5559
rect 152642 5556 152648 5568
rect 149379 5528 152648 5556
rect 149379 5525 149391 5528
rect 149333 5519 149391 5525
rect 152642 5516 152648 5528
rect 152700 5516 152706 5568
rect 152826 5516 152832 5568
rect 152884 5516 152890 5568
rect 153948 5556 153976 5655
rect 154942 5652 154948 5704
rect 155000 5652 155006 5704
rect 156693 5695 156751 5701
rect 156693 5692 156705 5695
rect 156616 5664 156705 5692
rect 155589 5627 155647 5633
rect 155589 5593 155601 5627
rect 155635 5624 155647 5627
rect 155954 5624 155960 5636
rect 155635 5596 155960 5624
rect 155635 5593 155647 5596
rect 155589 5587 155647 5593
rect 155954 5584 155960 5596
rect 156012 5584 156018 5636
rect 156230 5584 156236 5636
rect 156288 5624 156294 5636
rect 156371 5627 156429 5633
rect 156371 5624 156383 5627
rect 156288 5596 156383 5624
rect 156288 5584 156294 5596
rect 156371 5593 156383 5596
rect 156417 5593 156429 5627
rect 156371 5587 156429 5593
rect 154850 5556 154856 5568
rect 153948 5528 154856 5556
rect 154850 5516 154856 5528
rect 154908 5516 154914 5568
rect 156616 5556 156644 5664
rect 156693 5661 156705 5664
rect 156739 5661 156751 5695
rect 159726 5692 159732 5704
rect 156693 5655 156751 5661
rect 156785 5661 156843 5667
rect 156785 5627 156797 5661
rect 156831 5658 156843 5661
rect 156874 5658 156880 5670
rect 156831 5630 156880 5658
rect 156831 5627 156843 5630
rect 156785 5621 156843 5627
rect 156874 5618 156880 5630
rect 156932 5658 156938 5670
rect 156984 5664 159732 5692
rect 156984 5658 157012 5664
rect 156932 5630 157012 5658
rect 159726 5652 159732 5664
rect 159784 5652 159790 5704
rect 159818 5652 159824 5704
rect 159876 5692 159882 5704
rect 166966 5692 166994 5732
rect 169662 5720 169668 5732
rect 169720 5720 169726 5772
rect 185486 5720 185492 5772
rect 185544 5760 185550 5772
rect 189813 5763 189871 5769
rect 189813 5760 189825 5763
rect 185544 5732 189825 5760
rect 185544 5720 185550 5732
rect 189813 5729 189825 5732
rect 189859 5760 189871 5763
rect 190365 5763 190423 5769
rect 190365 5760 190377 5763
rect 189859 5732 190377 5760
rect 189859 5729 189871 5732
rect 189813 5723 189871 5729
rect 190365 5729 190377 5732
rect 190411 5760 190423 5763
rect 215846 5760 215852 5772
rect 190411 5732 215852 5760
rect 190411 5729 190423 5732
rect 190365 5723 190423 5729
rect 215846 5720 215852 5732
rect 215904 5760 215910 5772
rect 216401 5763 216459 5769
rect 216401 5760 216413 5763
rect 215904 5732 216413 5760
rect 215904 5720 215910 5732
rect 216401 5729 216413 5732
rect 216447 5760 216459 5763
rect 216769 5763 216827 5769
rect 216769 5760 216781 5763
rect 216447 5732 216781 5760
rect 216447 5729 216459 5732
rect 216401 5723 216459 5729
rect 216769 5729 216781 5732
rect 216815 5729 216827 5763
rect 216769 5723 216827 5729
rect 217042 5720 217048 5772
rect 217100 5720 217106 5772
rect 220541 5763 220599 5769
rect 220541 5760 220553 5763
rect 217152 5732 220553 5760
rect 159876 5664 166994 5692
rect 168009 5695 168067 5701
rect 159876 5652 159882 5664
rect 168009 5661 168021 5695
rect 168055 5692 168067 5695
rect 168282 5692 168288 5704
rect 168055 5664 168288 5692
rect 168055 5661 168067 5664
rect 168009 5655 168067 5661
rect 168282 5652 168288 5664
rect 168340 5652 168346 5704
rect 168834 5652 168840 5704
rect 168892 5652 168898 5704
rect 169202 5652 169208 5704
rect 169260 5652 169266 5704
rect 169846 5652 169852 5704
rect 169904 5652 169910 5704
rect 188798 5652 188804 5704
rect 188856 5692 188862 5704
rect 189445 5695 189503 5701
rect 189445 5692 189457 5695
rect 188856 5664 189457 5692
rect 188856 5652 188862 5664
rect 189445 5661 189457 5664
rect 189491 5661 189503 5695
rect 189445 5655 189503 5661
rect 207290 5652 207296 5704
rect 207348 5652 207354 5704
rect 212810 5652 212816 5704
rect 212868 5652 212874 5704
rect 213273 5695 213331 5701
rect 213273 5661 213285 5695
rect 213319 5661 213331 5695
rect 213273 5655 213331 5661
rect 156932 5618 156938 5630
rect 157153 5627 157211 5633
rect 157153 5593 157165 5627
rect 157199 5624 157211 5627
rect 157242 5624 157248 5636
rect 157199 5596 157248 5624
rect 157199 5593 157211 5596
rect 157153 5587 157211 5593
rect 157242 5584 157248 5596
rect 157300 5584 157306 5636
rect 157521 5627 157579 5633
rect 157521 5593 157533 5627
rect 157567 5624 157579 5627
rect 158622 5624 158628 5636
rect 157567 5596 158628 5624
rect 157567 5593 157579 5596
rect 157521 5587 157579 5593
rect 158622 5584 158628 5596
rect 158680 5584 158686 5636
rect 168650 5584 168656 5636
rect 168708 5624 168714 5636
rect 169941 5627 169999 5633
rect 169941 5624 169953 5627
rect 168708 5596 169953 5624
rect 168708 5584 168714 5596
rect 169941 5593 169953 5596
rect 169987 5624 169999 5627
rect 189534 5624 189540 5636
rect 169987 5596 189540 5624
rect 169987 5593 169999 5596
rect 169941 5587 169999 5593
rect 189534 5584 189540 5596
rect 189592 5624 189598 5636
rect 189930 5627 189988 5633
rect 189930 5624 189942 5627
rect 189592 5596 189942 5624
rect 189592 5584 189598 5596
rect 189930 5593 189942 5596
rect 189976 5593 189988 5627
rect 189930 5587 189988 5593
rect 206738 5584 206744 5636
rect 206796 5624 206802 5636
rect 207106 5624 207112 5636
rect 206796 5596 207112 5624
rect 206796 5584 206802 5596
rect 207106 5584 207112 5596
rect 207164 5584 207170 5636
rect 207474 5584 207480 5636
rect 207532 5584 207538 5636
rect 209130 5584 209136 5636
rect 209188 5624 209194 5636
rect 213288 5624 213316 5655
rect 213362 5652 213368 5704
rect 213420 5652 213426 5704
rect 213638 5652 213644 5704
rect 213696 5652 213702 5704
rect 215202 5652 215208 5704
rect 215260 5692 215266 5704
rect 215389 5695 215447 5701
rect 215389 5692 215401 5695
rect 215260 5664 215401 5692
rect 215260 5652 215266 5664
rect 215389 5661 215401 5664
rect 215435 5661 215447 5695
rect 215389 5655 215447 5661
rect 216490 5652 216496 5704
rect 216548 5692 216554 5704
rect 217152 5692 217180 5732
rect 220541 5729 220553 5732
rect 220587 5729 220599 5763
rect 220541 5723 220599 5729
rect 220814 5720 220820 5772
rect 220872 5720 220878 5772
rect 222930 5720 222936 5772
rect 222988 5760 222994 5772
rect 223117 5763 223175 5769
rect 223117 5760 223129 5763
rect 222988 5732 223129 5760
rect 222988 5720 222994 5732
rect 223117 5729 223129 5732
rect 223163 5729 223175 5763
rect 223316 5760 223344 5788
rect 223117 5723 223175 5729
rect 223224 5732 223344 5760
rect 223224 5704 223252 5732
rect 223482 5720 223488 5772
rect 223540 5760 223546 5772
rect 223761 5763 223819 5769
rect 223761 5760 223773 5763
rect 223540 5732 223773 5760
rect 223540 5720 223546 5732
rect 223761 5729 223773 5732
rect 223807 5729 223819 5763
rect 223761 5723 223819 5729
rect 224034 5720 224040 5772
rect 224092 5720 224098 5772
rect 224175 5763 224233 5769
rect 224175 5729 224187 5763
rect 224221 5760 224233 5763
rect 226058 5760 226064 5772
rect 224221 5732 226064 5760
rect 224221 5729 224233 5732
rect 224175 5723 224233 5729
rect 226058 5720 226064 5732
rect 226116 5720 226122 5772
rect 226168 5760 226196 5800
rect 226426 5788 226432 5840
rect 226484 5828 226490 5840
rect 226610 5828 226616 5840
rect 226484 5800 226616 5828
rect 226484 5788 226490 5800
rect 226610 5788 226616 5800
rect 226668 5788 226674 5840
rect 227622 5788 227628 5840
rect 227680 5828 227686 5840
rect 236454 5828 236460 5840
rect 227680 5800 236460 5828
rect 227680 5788 227686 5800
rect 236454 5788 236460 5800
rect 236512 5788 236518 5840
rect 247678 5788 247684 5840
rect 247736 5828 247742 5840
rect 248414 5828 248420 5840
rect 247736 5800 248420 5828
rect 247736 5788 247742 5800
rect 248414 5788 248420 5800
rect 248472 5788 248478 5840
rect 248506 5788 248512 5840
rect 248564 5828 248570 5840
rect 249153 5831 249211 5837
rect 249153 5828 249165 5831
rect 248564 5800 249165 5828
rect 248564 5788 248570 5800
rect 249153 5797 249165 5800
rect 249199 5797 249211 5831
rect 249153 5791 249211 5797
rect 249426 5788 249432 5840
rect 249484 5828 249490 5840
rect 250533 5831 250591 5837
rect 250533 5828 250545 5831
rect 249484 5800 250545 5828
rect 249484 5788 249490 5800
rect 250533 5797 250545 5800
rect 250579 5797 250591 5831
rect 250533 5791 250591 5797
rect 250622 5788 250628 5840
rect 250680 5828 250686 5840
rect 250990 5828 250996 5840
rect 250680 5800 250996 5828
rect 250680 5788 250686 5800
rect 250990 5788 250996 5800
rect 251048 5828 251054 5840
rect 253906 5828 253934 5868
rect 256326 5856 256332 5868
rect 256384 5856 256390 5908
rect 259365 5899 259423 5905
rect 259365 5865 259377 5899
rect 259411 5896 259423 5899
rect 260834 5896 260840 5908
rect 259411 5868 260840 5896
rect 259411 5865 259423 5868
rect 259365 5859 259423 5865
rect 260834 5856 260840 5868
rect 260892 5856 260898 5908
rect 263134 5856 263140 5908
rect 263192 5856 263198 5908
rect 264882 5896 264888 5908
rect 263566 5868 264888 5896
rect 251048 5800 253934 5828
rect 251048 5788 251054 5800
rect 254578 5788 254584 5840
rect 254636 5788 254642 5840
rect 254670 5788 254676 5840
rect 254728 5828 254734 5840
rect 256786 5828 256792 5840
rect 254728 5800 256792 5828
rect 254728 5788 254734 5800
rect 256786 5788 256792 5800
rect 256844 5788 256850 5840
rect 259546 5828 259552 5840
rect 259380 5800 259552 5828
rect 239030 5760 239036 5772
rect 226168 5732 239036 5760
rect 239030 5720 239036 5732
rect 239088 5720 239094 5772
rect 245562 5720 245568 5772
rect 245620 5760 245626 5772
rect 247034 5760 247040 5772
rect 245620 5732 247040 5760
rect 245620 5720 245626 5732
rect 247034 5720 247040 5732
rect 247092 5720 247098 5772
rect 247865 5763 247923 5769
rect 247865 5760 247877 5763
rect 247144 5732 247877 5760
rect 216548 5664 217180 5692
rect 216548 5652 216554 5664
rect 217870 5652 217876 5704
rect 217928 5692 217934 5704
rect 218241 5695 218299 5701
rect 218241 5692 218253 5695
rect 217928 5664 218253 5692
rect 217928 5652 217934 5664
rect 216030 5624 216036 5636
rect 209188 5596 211200 5624
rect 213288 5596 216036 5624
rect 209188 5584 209194 5596
rect 156782 5556 156788 5568
rect 156616 5528 156788 5556
rect 156782 5516 156788 5528
rect 156840 5516 156846 5568
rect 167454 5516 167460 5568
rect 167512 5556 167518 5568
rect 168193 5559 168251 5565
rect 168193 5556 168205 5559
rect 167512 5528 168205 5556
rect 167512 5516 167518 5528
rect 168193 5525 168205 5528
rect 168239 5525 168251 5559
rect 168193 5519 168251 5525
rect 169386 5516 169392 5568
rect 169444 5516 169450 5568
rect 171042 5516 171048 5568
rect 171100 5556 171106 5568
rect 172606 5556 172612 5568
rect 171100 5528 172612 5556
rect 171100 5516 171106 5528
rect 172606 5516 172612 5528
rect 172664 5516 172670 5568
rect 189350 5516 189356 5568
rect 189408 5556 189414 5568
rect 189721 5559 189779 5565
rect 189721 5556 189733 5559
rect 189408 5528 189733 5556
rect 189408 5516 189414 5528
rect 189721 5525 189733 5528
rect 189767 5525 189779 5559
rect 189721 5519 189779 5525
rect 200758 5516 200764 5568
rect 200816 5556 200822 5568
rect 210418 5556 210424 5568
rect 200816 5528 210424 5556
rect 200816 5516 200822 5528
rect 210418 5516 210424 5528
rect 210476 5516 210482 5568
rect 211172 5556 211200 5596
rect 216030 5584 216036 5596
rect 216088 5584 216094 5636
rect 216125 5627 216183 5633
rect 216125 5593 216137 5627
rect 216171 5624 216183 5627
rect 216674 5624 216680 5636
rect 216171 5596 216680 5624
rect 216171 5593 216183 5596
rect 216125 5587 216183 5593
rect 216674 5584 216680 5596
rect 216732 5624 216738 5636
rect 217226 5624 217232 5636
rect 217284 5633 217290 5636
rect 217284 5627 217312 5633
rect 216732 5596 217232 5624
rect 216732 5584 216738 5596
rect 217226 5584 217232 5596
rect 217300 5593 217312 5627
rect 217284 5587 217312 5593
rect 217284 5584 217290 5587
rect 215110 5556 215116 5568
rect 211172 5528 215116 5556
rect 215110 5516 215116 5528
rect 215168 5516 215174 5568
rect 215205 5559 215263 5565
rect 215205 5525 215217 5559
rect 215251 5556 215263 5559
rect 216214 5556 216220 5568
rect 215251 5528 216220 5556
rect 215251 5525 215263 5528
rect 215205 5519 215263 5525
rect 216214 5516 216220 5528
rect 216272 5516 216278 5568
rect 217134 5516 217140 5568
rect 217192 5516 217198 5568
rect 217980 5556 218008 5664
rect 218241 5661 218253 5664
rect 218287 5661 218299 5695
rect 218241 5655 218299 5661
rect 218330 5652 218336 5704
rect 218388 5652 218394 5704
rect 218517 5695 218575 5701
rect 218517 5661 218529 5695
rect 218563 5661 218575 5695
rect 218517 5655 218575 5661
rect 218054 5584 218060 5636
rect 218112 5624 218118 5636
rect 218532 5624 218560 5655
rect 218790 5652 218796 5704
rect 218848 5692 218854 5704
rect 219526 5692 219532 5704
rect 218848 5664 219532 5692
rect 218848 5652 218854 5664
rect 219526 5652 219532 5664
rect 219584 5652 219590 5704
rect 220357 5695 220415 5701
rect 220357 5692 220369 5695
rect 220280 5664 220369 5692
rect 218112 5596 218560 5624
rect 218885 5627 218943 5633
rect 218112 5584 218118 5596
rect 218885 5593 218897 5627
rect 218931 5624 218943 5627
rect 220078 5624 220084 5636
rect 218931 5596 220084 5624
rect 218931 5593 218943 5596
rect 218885 5587 218943 5593
rect 220078 5584 220084 5596
rect 220136 5584 220142 5636
rect 220280 5595 220308 5664
rect 220357 5661 220369 5664
rect 220403 5661 220415 5695
rect 220357 5655 220415 5661
rect 223206 5652 223212 5704
rect 223264 5652 223270 5704
rect 223298 5652 223304 5704
rect 223356 5652 223362 5704
rect 224310 5652 224316 5704
rect 224368 5652 224374 5704
rect 224954 5652 224960 5704
rect 225012 5692 225018 5704
rect 225509 5695 225567 5701
rect 225509 5692 225521 5695
rect 225012 5664 225521 5692
rect 225012 5652 225018 5664
rect 225509 5661 225521 5664
rect 225555 5692 225567 5695
rect 225690 5692 225696 5704
rect 225555 5664 225696 5692
rect 225555 5661 225567 5664
rect 225509 5655 225567 5661
rect 225690 5652 225696 5664
rect 225748 5652 225754 5704
rect 246850 5652 246856 5704
rect 246908 5692 246914 5704
rect 247144 5692 247172 5732
rect 247865 5729 247877 5732
rect 247911 5729 247923 5763
rect 247865 5723 247923 5729
rect 247954 5720 247960 5772
rect 248012 5760 248018 5772
rect 248322 5760 248328 5772
rect 248012 5732 248328 5760
rect 248012 5720 248018 5732
rect 248322 5720 248328 5732
rect 248380 5760 248386 5772
rect 248877 5763 248935 5769
rect 248877 5760 248889 5763
rect 248380 5732 248889 5760
rect 248380 5720 248386 5732
rect 248877 5729 248889 5732
rect 248923 5760 248935 5763
rect 249794 5760 249800 5772
rect 248923 5732 249800 5760
rect 248923 5729 248935 5732
rect 248877 5723 248935 5729
rect 249794 5720 249800 5732
rect 249852 5720 249858 5772
rect 249978 5720 249984 5772
rect 250036 5760 250042 5772
rect 253290 5760 253296 5772
rect 250036 5732 253296 5760
rect 250036 5720 250042 5732
rect 253290 5720 253296 5732
rect 253348 5720 253354 5772
rect 259380 5769 259408 5800
rect 259546 5788 259552 5800
rect 259604 5788 259610 5840
rect 263566 5828 263594 5868
rect 264882 5856 264888 5868
rect 264940 5856 264946 5908
rect 265250 5856 265256 5908
rect 265308 5856 265314 5908
rect 265434 5856 265440 5908
rect 265492 5896 265498 5908
rect 265894 5896 265900 5908
rect 265492 5868 265900 5896
rect 265492 5856 265498 5868
rect 265894 5856 265900 5868
rect 265952 5856 265958 5908
rect 266170 5856 266176 5908
rect 266228 5896 266234 5908
rect 269022 5896 269028 5908
rect 266228 5868 269028 5896
rect 266228 5856 266234 5868
rect 269022 5856 269028 5868
rect 269080 5856 269086 5908
rect 268378 5828 268384 5840
rect 261036 5800 263594 5828
rect 263796 5800 268384 5828
rect 255041 5763 255099 5769
rect 255041 5760 255053 5763
rect 253400 5732 255053 5760
rect 246908 5664 247172 5692
rect 247313 5695 247371 5701
rect 246908 5652 246914 5664
rect 247313 5661 247325 5695
rect 247359 5692 247371 5695
rect 248049 5695 248107 5701
rect 247359 5664 248000 5692
rect 247359 5661 247371 5664
rect 247313 5655 247371 5661
rect 227070 5624 227076 5636
rect 224788 5596 227076 5624
rect 219710 5556 219716 5568
rect 217980 5528 219716 5556
rect 219710 5516 219716 5528
rect 219768 5516 219774 5568
rect 220280 5567 220400 5595
rect 220372 5556 220400 5567
rect 224788 5556 224816 5596
rect 227070 5584 227076 5596
rect 227128 5584 227134 5636
rect 227714 5584 227720 5636
rect 227772 5624 227778 5636
rect 243078 5624 243084 5636
rect 227772 5596 243084 5624
rect 227772 5584 227778 5596
rect 243078 5584 243084 5596
rect 243136 5584 243142 5636
rect 247034 5584 247040 5636
rect 247092 5624 247098 5636
rect 247770 5624 247776 5636
rect 247092 5596 247776 5624
rect 247092 5584 247098 5596
rect 247770 5584 247776 5596
rect 247828 5584 247834 5636
rect 247972 5624 248000 5664
rect 248049 5661 248061 5695
rect 248095 5692 248107 5695
rect 248230 5692 248236 5704
rect 248095 5664 248236 5692
rect 248095 5661 248107 5664
rect 248049 5655 248107 5661
rect 248230 5652 248236 5664
rect 248288 5652 248294 5704
rect 248414 5652 248420 5704
rect 248472 5692 248478 5704
rect 248969 5695 249027 5701
rect 248472 5664 248736 5692
rect 248472 5652 248478 5664
rect 248708 5633 248736 5664
rect 248969 5661 248981 5695
rect 249015 5692 249027 5695
rect 249150 5692 249156 5704
rect 249015 5664 249156 5692
rect 249015 5661 249027 5664
rect 248969 5655 249027 5661
rect 249150 5652 249156 5664
rect 249208 5692 249214 5704
rect 249889 5695 249947 5701
rect 249889 5692 249901 5695
rect 249208 5664 249901 5692
rect 249208 5652 249214 5664
rect 249889 5661 249901 5664
rect 249935 5692 249947 5695
rect 250530 5692 250536 5704
rect 249935 5664 250536 5692
rect 249935 5661 249947 5664
rect 249889 5655 249947 5661
rect 250530 5652 250536 5664
rect 250588 5652 250594 5704
rect 250714 5652 250720 5704
rect 250772 5652 250778 5704
rect 253400 5692 253428 5732
rect 255041 5729 255053 5732
rect 255087 5760 255099 5763
rect 259365 5763 259423 5769
rect 255087 5732 259316 5760
rect 255087 5729 255099 5732
rect 255041 5723 255099 5729
rect 251146 5664 253428 5692
rect 248693 5627 248751 5633
rect 247972 5596 248644 5624
rect 220372 5528 224816 5556
rect 238754 5516 238760 5568
rect 238812 5556 238818 5568
rect 242986 5556 242992 5568
rect 238812 5528 242992 5556
rect 238812 5516 238818 5528
rect 242986 5516 242992 5528
rect 243044 5516 243050 5568
rect 247129 5559 247187 5565
rect 247129 5525 247141 5559
rect 247175 5556 247187 5559
rect 248506 5556 248512 5568
rect 247175 5528 248512 5556
rect 247175 5525 247187 5528
rect 247129 5519 247187 5525
rect 248506 5516 248512 5528
rect 248564 5516 248570 5568
rect 248616 5556 248644 5596
rect 248693 5593 248705 5627
rect 248739 5624 248751 5627
rect 249334 5624 249340 5636
rect 248739 5596 249340 5624
rect 248739 5593 248751 5596
rect 248693 5587 248751 5593
rect 249334 5584 249340 5596
rect 249392 5624 249398 5636
rect 249613 5627 249671 5633
rect 249613 5624 249625 5627
rect 249392 5596 249625 5624
rect 249392 5584 249398 5596
rect 249613 5593 249625 5596
rect 249659 5624 249671 5627
rect 249659 5596 250576 5624
rect 249659 5593 249671 5596
rect 249613 5587 249671 5593
rect 249978 5556 249984 5568
rect 248616 5528 249984 5556
rect 249978 5516 249984 5528
rect 250036 5516 250042 5568
rect 250073 5559 250131 5565
rect 250073 5525 250085 5559
rect 250119 5556 250131 5559
rect 250438 5556 250444 5568
rect 250119 5528 250444 5556
rect 250119 5525 250131 5528
rect 250073 5519 250131 5525
rect 250438 5516 250444 5528
rect 250496 5516 250502 5568
rect 250548 5556 250576 5596
rect 251146 5556 251174 5664
rect 253842 5652 253848 5704
rect 253900 5652 253906 5704
rect 255317 5695 255375 5701
rect 255317 5661 255329 5695
rect 255363 5692 255375 5695
rect 255406 5692 255412 5704
rect 255363 5664 255412 5692
rect 255363 5661 255375 5664
rect 255317 5655 255375 5661
rect 255406 5652 255412 5664
rect 255464 5652 255470 5704
rect 256326 5652 256332 5704
rect 256384 5692 256390 5704
rect 256421 5695 256479 5701
rect 256421 5692 256433 5695
rect 256384 5664 256433 5692
rect 256384 5652 256390 5664
rect 256421 5661 256433 5664
rect 256467 5661 256479 5695
rect 256421 5655 256479 5661
rect 256697 5695 256755 5701
rect 256697 5661 256709 5695
rect 256743 5692 256755 5695
rect 256786 5692 256792 5704
rect 256743 5664 256792 5692
rect 256743 5661 256755 5664
rect 256697 5655 256755 5661
rect 256786 5652 256792 5664
rect 256844 5692 256850 5704
rect 257614 5692 257620 5704
rect 256844 5664 257620 5692
rect 256844 5652 256850 5664
rect 257614 5652 257620 5664
rect 257672 5652 257678 5704
rect 257893 5695 257951 5701
rect 257893 5661 257905 5695
rect 257939 5692 257951 5695
rect 259178 5692 259184 5704
rect 257939 5664 259184 5692
rect 257939 5661 257951 5664
rect 257893 5655 257951 5661
rect 259178 5652 259184 5664
rect 259236 5652 259242 5704
rect 259288 5701 259316 5732
rect 259365 5729 259377 5763
rect 259411 5729 259423 5763
rect 260926 5760 260932 5772
rect 259365 5723 259423 5729
rect 259472 5732 260932 5760
rect 259273 5695 259331 5701
rect 259273 5661 259285 5695
rect 259319 5692 259331 5695
rect 259472 5692 259500 5732
rect 260926 5720 260932 5732
rect 260984 5720 260990 5772
rect 259319 5664 259500 5692
rect 259549 5695 259607 5701
rect 259319 5661 259331 5664
rect 259273 5655 259331 5661
rect 259549 5661 259561 5695
rect 259595 5692 259607 5695
rect 259638 5692 259644 5704
rect 259595 5664 259644 5692
rect 259595 5661 259607 5664
rect 259549 5655 259607 5661
rect 259638 5652 259644 5664
rect 259696 5652 259702 5704
rect 260374 5652 260380 5704
rect 260432 5652 260438 5704
rect 261036 5692 261064 5800
rect 261570 5720 261576 5772
rect 261628 5760 261634 5772
rect 261628 5732 262996 5760
rect 261628 5720 261634 5732
rect 260484 5664 261064 5692
rect 251266 5584 251272 5636
rect 251324 5624 251330 5636
rect 254302 5624 254308 5636
rect 251324 5596 254308 5624
rect 251324 5584 251330 5596
rect 254302 5584 254308 5596
rect 254360 5584 254366 5636
rect 254394 5584 254400 5636
rect 254452 5624 254458 5636
rect 259454 5624 259460 5636
rect 254452 5596 259460 5624
rect 254452 5584 254458 5596
rect 259454 5584 259460 5596
rect 259512 5584 259518 5636
rect 260484 5624 260512 5664
rect 261662 5652 261668 5704
rect 261720 5652 261726 5704
rect 259564 5596 260512 5624
rect 250548 5528 251174 5556
rect 253661 5559 253719 5565
rect 253661 5525 253673 5559
rect 253707 5556 253719 5559
rect 254210 5556 254216 5568
rect 253707 5528 254216 5556
rect 253707 5525 253719 5528
rect 253661 5519 253719 5525
rect 254210 5516 254216 5528
rect 254268 5516 254274 5568
rect 255682 5516 255688 5568
rect 255740 5556 255746 5568
rect 257709 5559 257767 5565
rect 257709 5556 257721 5559
rect 255740 5528 257721 5556
rect 255740 5516 255746 5528
rect 257709 5525 257721 5528
rect 257755 5525 257767 5559
rect 257709 5519 257767 5525
rect 257798 5516 257804 5568
rect 257856 5556 257862 5568
rect 259564 5556 259592 5596
rect 260742 5584 260748 5636
rect 260800 5584 260806 5636
rect 261018 5584 261024 5636
rect 261076 5624 261082 5636
rect 262033 5627 262091 5633
rect 262033 5624 262045 5627
rect 261076 5596 262045 5624
rect 261076 5584 261082 5596
rect 262033 5593 262045 5596
rect 262079 5593 262091 5627
rect 262033 5587 262091 5593
rect 257856 5528 259592 5556
rect 259733 5559 259791 5565
rect 257856 5516 257862 5528
rect 259733 5525 259745 5559
rect 259779 5556 259791 5559
rect 259822 5556 259828 5568
rect 259779 5528 259828 5556
rect 259779 5525 259791 5528
rect 259733 5519 259791 5525
rect 259822 5516 259828 5528
rect 259880 5516 259886 5568
rect 262784 5556 262812 5732
rect 262968 5701 262996 5732
rect 263796 5701 263824 5800
rect 268378 5788 268384 5800
rect 268436 5788 268442 5840
rect 268930 5788 268936 5840
rect 268988 5828 268994 5840
rect 270497 5831 270555 5837
rect 270497 5828 270509 5831
rect 268988 5800 270509 5828
rect 268988 5788 268994 5800
rect 270497 5797 270509 5800
rect 270543 5797 270555 5831
rect 270497 5791 270555 5797
rect 264974 5760 264980 5772
rect 264624 5732 264980 5760
rect 262861 5695 262919 5701
rect 262861 5661 262873 5695
rect 262907 5661 262919 5695
rect 262861 5655 262919 5661
rect 262953 5695 263011 5701
rect 262953 5661 262965 5695
rect 262999 5661 263011 5695
rect 262953 5655 263011 5661
rect 263781 5695 263839 5701
rect 263781 5661 263793 5695
rect 263827 5661 263839 5695
rect 263781 5655 263839 5661
rect 264333 5695 264391 5701
rect 264333 5661 264345 5695
rect 264379 5692 264391 5695
rect 264422 5692 264428 5704
rect 264379 5664 264428 5692
rect 264379 5661 264391 5664
rect 264333 5655 264391 5661
rect 262876 5624 262904 5655
rect 264422 5652 264428 5664
rect 264480 5652 264486 5704
rect 264624 5624 264652 5732
rect 264974 5720 264980 5732
rect 265032 5720 265038 5772
rect 265250 5720 265256 5772
rect 265308 5760 265314 5772
rect 268286 5760 268292 5772
rect 265308 5732 268292 5760
rect 265308 5720 265314 5732
rect 268286 5720 268292 5732
rect 268344 5720 268350 5772
rect 269853 5763 269911 5769
rect 269853 5760 269865 5763
rect 268396 5732 269865 5760
rect 264882 5652 264888 5704
rect 264940 5652 264946 5704
rect 265069 5695 265127 5701
rect 265069 5661 265081 5695
rect 265115 5692 265127 5695
rect 265710 5692 265716 5704
rect 265115 5664 265716 5692
rect 265115 5661 265127 5664
rect 265069 5655 265127 5661
rect 265710 5652 265716 5664
rect 265768 5652 265774 5704
rect 265897 5695 265955 5701
rect 265897 5661 265909 5695
rect 265943 5661 265955 5695
rect 265897 5655 265955 5661
rect 265912 5624 265940 5655
rect 266906 5652 266912 5704
rect 266964 5652 266970 5704
rect 268396 5701 268424 5732
rect 269853 5729 269865 5732
rect 269899 5729 269911 5763
rect 269853 5723 269911 5729
rect 268381 5695 268439 5701
rect 268381 5661 268393 5695
rect 268427 5661 268439 5695
rect 268381 5655 268439 5661
rect 269574 5652 269580 5704
rect 269632 5652 269638 5704
rect 269669 5695 269727 5701
rect 269669 5661 269681 5695
rect 269715 5661 269727 5695
rect 269669 5655 269727 5661
rect 262876 5596 264652 5624
rect 265084 5596 265940 5624
rect 265084 5556 265112 5596
rect 266354 5584 266360 5636
rect 266412 5624 266418 5636
rect 267277 5627 267335 5633
rect 267277 5624 267289 5627
rect 266412 5596 267289 5624
rect 266412 5584 266418 5596
rect 267277 5593 267289 5596
rect 267323 5593 267335 5627
rect 267277 5587 267335 5593
rect 268010 5584 268016 5636
rect 268068 5624 268074 5636
rect 268749 5627 268807 5633
rect 268749 5624 268761 5627
rect 268068 5596 268761 5624
rect 268068 5584 268074 5596
rect 268749 5593 268761 5596
rect 268795 5593 268807 5627
rect 269684 5624 269712 5655
rect 269942 5652 269948 5704
rect 270000 5692 270006 5704
rect 270313 5695 270371 5701
rect 270313 5692 270325 5695
rect 270000 5664 270325 5692
rect 270000 5652 270006 5664
rect 270313 5661 270325 5664
rect 270359 5661 270371 5695
rect 270313 5655 270371 5661
rect 269850 5624 269856 5636
rect 269684 5596 269856 5624
rect 268749 5587 268807 5593
rect 269850 5584 269856 5596
rect 269908 5584 269914 5636
rect 271230 5624 271236 5636
rect 271064 5596 271236 5624
rect 262784 5528 265112 5556
rect 265710 5516 265716 5568
rect 265768 5556 265774 5568
rect 265986 5556 265992 5568
rect 265768 5528 265992 5556
rect 265768 5516 265774 5528
rect 265986 5516 265992 5528
rect 266044 5516 266050 5568
rect 267090 5516 267096 5568
rect 267148 5556 267154 5568
rect 271064 5556 271092 5596
rect 271230 5584 271236 5596
rect 271288 5584 271294 5636
rect 267148 5528 271092 5556
rect 267148 5516 267154 5528
rect 271138 5516 271144 5568
rect 271196 5556 271202 5568
rect 271782 5556 271788 5568
rect 271196 5528 271788 5556
rect 271196 5516 271202 5528
rect 271782 5516 271788 5528
rect 271840 5516 271846 5568
rect 1104 5466 271651 5488
rect 1104 5414 68546 5466
rect 68598 5414 68610 5466
rect 68662 5414 68674 5466
rect 68726 5414 68738 5466
rect 68790 5414 68802 5466
rect 68854 5414 136143 5466
rect 136195 5414 136207 5466
rect 136259 5414 136271 5466
rect 136323 5414 136335 5466
rect 136387 5414 136399 5466
rect 136451 5414 203740 5466
rect 203792 5414 203804 5466
rect 203856 5414 203868 5466
rect 203920 5414 203932 5466
rect 203984 5414 203996 5466
rect 204048 5414 271337 5466
rect 271389 5414 271401 5466
rect 271453 5414 271465 5466
rect 271517 5414 271529 5466
rect 271581 5414 271593 5466
rect 271645 5414 271651 5466
rect 1104 5392 271651 5414
rect 35529 5355 35587 5361
rect 35529 5321 35541 5355
rect 35575 5352 35587 5355
rect 36078 5352 36084 5364
rect 35575 5324 36084 5352
rect 35575 5321 35587 5324
rect 35529 5315 35587 5321
rect 36078 5312 36084 5324
rect 36136 5312 36142 5364
rect 36998 5312 37004 5364
rect 37056 5352 37062 5364
rect 37056 5324 94360 5352
rect 37056 5312 37062 5324
rect 35802 5244 35808 5296
rect 35860 5244 35866 5296
rect 36262 5244 36268 5296
rect 36320 5244 36326 5296
rect 36633 5287 36691 5293
rect 36633 5253 36645 5287
rect 36679 5253 36691 5287
rect 36633 5247 36691 5253
rect 35894 5176 35900 5228
rect 35952 5176 35958 5228
rect 35986 5176 35992 5228
rect 36044 5216 36050 5228
rect 36648 5216 36676 5247
rect 45830 5244 45836 5296
rect 45888 5244 45894 5296
rect 46014 5244 46020 5296
rect 46072 5284 46078 5296
rect 46109 5287 46167 5293
rect 46109 5284 46121 5287
rect 46072 5256 46121 5284
rect 46072 5244 46078 5256
rect 46109 5253 46121 5256
rect 46155 5253 46167 5287
rect 46109 5247 46167 5253
rect 46658 5244 46664 5296
rect 46716 5284 46722 5296
rect 46937 5287 46995 5293
rect 46937 5284 46949 5287
rect 46716 5256 46949 5284
rect 46716 5244 46722 5256
rect 46937 5253 46949 5256
rect 46983 5253 46995 5287
rect 46937 5247 46995 5253
rect 50448 5256 50936 5284
rect 36044 5188 36676 5216
rect 36044 5176 36050 5188
rect 36722 5176 36728 5228
rect 36780 5216 36786 5228
rect 44082 5216 44088 5228
rect 36780 5188 44088 5216
rect 36780 5176 36786 5188
rect 44082 5176 44088 5188
rect 44140 5176 44146 5228
rect 46198 5176 46204 5228
rect 46256 5176 46262 5228
rect 46566 5176 46572 5228
rect 46624 5176 46630 5228
rect 46750 5176 46756 5228
rect 46808 5216 46814 5228
rect 50448 5225 50476 5256
rect 50433 5219 50491 5225
rect 50433 5216 50445 5219
rect 46808 5188 50445 5216
rect 46808 5176 46814 5188
rect 50433 5185 50445 5188
rect 50479 5185 50491 5219
rect 50908 5216 50936 5256
rect 50982 5244 50988 5296
rect 51040 5244 51046 5296
rect 52089 5287 52147 5293
rect 52089 5284 52101 5287
rect 51184 5256 52101 5284
rect 51184 5216 51212 5256
rect 52089 5253 52101 5256
rect 52135 5253 52147 5287
rect 52089 5247 52147 5253
rect 50908 5188 51212 5216
rect 50433 5179 50491 5185
rect 51258 5176 51264 5228
rect 51316 5176 51322 5228
rect 51350 5176 51356 5228
rect 51408 5176 51414 5228
rect 51718 5176 51724 5228
rect 51776 5176 51782 5228
rect 52917 5219 52975 5225
rect 52917 5185 52929 5219
rect 52963 5216 52975 5219
rect 53561 5219 53619 5225
rect 53561 5216 53573 5219
rect 52963 5188 53573 5216
rect 52963 5185 52975 5188
rect 52917 5179 52975 5185
rect 53561 5185 53573 5188
rect 53607 5216 53619 5219
rect 92382 5216 92388 5228
rect 53607 5188 92388 5216
rect 53607 5185 53619 5188
rect 53561 5179 53619 5185
rect 92382 5176 92388 5188
rect 92440 5176 92446 5228
rect 94332 5225 94360 5324
rect 95142 5312 95148 5364
rect 95200 5352 95206 5364
rect 96062 5352 96068 5364
rect 95200 5324 96068 5352
rect 95200 5312 95206 5324
rect 96062 5312 96068 5324
rect 96120 5312 96126 5364
rect 96154 5312 96160 5364
rect 96212 5352 96218 5364
rect 96430 5352 96436 5364
rect 96212 5324 96436 5352
rect 96212 5312 96218 5324
rect 96430 5312 96436 5324
rect 96488 5312 96494 5364
rect 96614 5312 96620 5364
rect 96672 5352 96678 5364
rect 96982 5352 96988 5364
rect 96672 5324 96988 5352
rect 96672 5312 96678 5324
rect 96982 5312 96988 5324
rect 97040 5352 97046 5364
rect 97994 5352 98000 5364
rect 97040 5324 98000 5352
rect 97040 5312 97046 5324
rect 97994 5312 98000 5324
rect 98052 5312 98058 5364
rect 98086 5312 98092 5364
rect 98144 5352 98150 5364
rect 99837 5355 99895 5361
rect 99837 5352 99849 5355
rect 98144 5324 99849 5352
rect 98144 5312 98150 5324
rect 99837 5321 99849 5324
rect 99883 5321 99895 5355
rect 99837 5315 99895 5321
rect 100018 5312 100024 5364
rect 100076 5352 100082 5364
rect 100849 5355 100907 5361
rect 100849 5352 100861 5355
rect 100076 5324 100861 5352
rect 100076 5312 100082 5324
rect 100849 5321 100861 5324
rect 100895 5321 100907 5355
rect 100849 5315 100907 5321
rect 101398 5312 101404 5364
rect 101456 5352 101462 5364
rect 101861 5355 101919 5361
rect 101861 5352 101873 5355
rect 101456 5324 101873 5352
rect 101456 5312 101462 5324
rect 101861 5321 101873 5324
rect 101907 5321 101919 5355
rect 101861 5315 101919 5321
rect 102689 5355 102747 5361
rect 102689 5321 102701 5355
rect 102735 5321 102747 5355
rect 102689 5315 102747 5321
rect 95234 5244 95240 5296
rect 95292 5284 95298 5296
rect 95292 5256 99512 5284
rect 95292 5244 95298 5256
rect 93581 5219 93639 5225
rect 93581 5185 93593 5219
rect 93627 5185 93639 5219
rect 93581 5179 93639 5185
rect 94317 5219 94375 5225
rect 94317 5185 94329 5219
rect 94363 5185 94375 5219
rect 94317 5179 94375 5185
rect 37090 5148 37096 5160
rect 36570 5120 37096 5148
rect 37090 5108 37096 5120
rect 37148 5108 37154 5160
rect 46474 5108 46480 5160
rect 46532 5108 46538 5160
rect 52086 5148 52092 5160
rect 52026 5120 52092 5148
rect 52086 5108 52092 5120
rect 52144 5148 52150 5160
rect 53006 5148 53012 5160
rect 52144 5120 53012 5148
rect 52144 5108 52150 5120
rect 53006 5108 53012 5120
rect 53064 5108 53070 5160
rect 93596 5148 93624 5179
rect 98454 5176 98460 5228
rect 98512 5176 98518 5228
rect 99285 5219 99343 5225
rect 99285 5185 99297 5219
rect 99331 5216 99343 5219
rect 99374 5216 99380 5228
rect 99331 5188 99380 5216
rect 99331 5185 99343 5188
rect 99285 5179 99343 5185
rect 99374 5176 99380 5188
rect 99432 5176 99438 5228
rect 99484 5216 99512 5256
rect 99558 5244 99564 5296
rect 99616 5284 99622 5296
rect 100386 5284 100392 5296
rect 99616 5256 100392 5284
rect 99616 5244 99622 5256
rect 100386 5244 100392 5256
rect 100444 5244 100450 5296
rect 101232 5256 102640 5284
rect 99484 5188 99972 5216
rect 94501 5151 94559 5157
rect 93596 5120 94452 5148
rect 38746 5040 38752 5092
rect 38804 5080 38810 5092
rect 40954 5080 40960 5092
rect 38804 5052 40960 5080
rect 38804 5040 38810 5052
rect 40954 5040 40960 5052
rect 41012 5080 41018 5092
rect 42242 5080 42248 5092
rect 41012 5052 42248 5080
rect 41012 5040 41018 5052
rect 42242 5040 42248 5052
rect 42300 5040 42306 5092
rect 47118 5040 47124 5092
rect 47176 5040 47182 5092
rect 52178 5040 52184 5092
rect 52236 5080 52242 5092
rect 52273 5083 52331 5089
rect 52273 5080 52285 5083
rect 52236 5052 52285 5080
rect 52236 5040 52242 5052
rect 52273 5049 52285 5052
rect 52319 5049 52331 5083
rect 52273 5043 52331 5049
rect 52362 5040 52368 5092
rect 52420 5080 52426 5092
rect 53101 5083 53159 5089
rect 53101 5080 53113 5083
rect 52420 5052 53113 5080
rect 52420 5040 52426 5052
rect 53101 5049 53113 5052
rect 53147 5049 53159 5083
rect 53101 5043 53159 5049
rect 55858 5040 55864 5092
rect 55916 5080 55922 5092
rect 94314 5080 94320 5092
rect 55916 5052 94320 5080
rect 55916 5040 55922 5052
rect 94314 5040 94320 5052
rect 94372 5040 94378 5092
rect 94424 5080 94452 5120
rect 94501 5117 94513 5151
rect 94547 5148 94559 5151
rect 95970 5148 95976 5160
rect 94547 5120 95976 5148
rect 94547 5117 94559 5120
rect 94501 5111 94559 5117
rect 95970 5108 95976 5120
rect 96028 5108 96034 5160
rect 96157 5151 96215 5157
rect 96157 5117 96169 5151
rect 96203 5117 96215 5151
rect 96157 5111 96215 5117
rect 95326 5080 95332 5092
rect 94424 5052 95332 5080
rect 95326 5040 95332 5052
rect 95384 5040 95390 5092
rect 96172 5080 96200 5111
rect 96614 5108 96620 5160
rect 96672 5108 96678 5160
rect 96801 5151 96859 5157
rect 96801 5117 96813 5151
rect 96847 5148 96859 5151
rect 97442 5148 97448 5160
rect 96847 5120 97448 5148
rect 96847 5117 96859 5120
rect 96801 5111 96859 5117
rect 97442 5108 97448 5120
rect 97500 5108 97506 5160
rect 97718 5108 97724 5160
rect 97776 5148 97782 5160
rect 98822 5148 98828 5160
rect 97776 5120 98828 5148
rect 97776 5108 97782 5120
rect 98822 5108 98828 5120
rect 98880 5108 98886 5160
rect 99558 5108 99564 5160
rect 99616 5108 99622 5160
rect 99944 5148 99972 5188
rect 100294 5176 100300 5228
rect 100352 5176 100358 5228
rect 101232 5216 101260 5256
rect 100496 5188 101260 5216
rect 100496 5148 100524 5188
rect 101306 5176 101312 5228
rect 101364 5176 101370 5228
rect 101674 5176 101680 5228
rect 101732 5176 101738 5228
rect 101858 5176 101864 5228
rect 101916 5216 101922 5228
rect 102318 5216 102324 5228
rect 101916 5188 102324 5216
rect 101916 5176 101922 5188
rect 102318 5176 102324 5188
rect 102376 5176 102382 5228
rect 99944 5120 100524 5148
rect 100570 5108 100576 5160
rect 100628 5148 100634 5160
rect 101692 5148 101720 5176
rect 100628 5120 101720 5148
rect 100628 5108 100634 5120
rect 102410 5108 102416 5160
rect 102468 5108 102474 5160
rect 102612 5148 102640 5256
rect 102704 5216 102732 5315
rect 108850 5312 108856 5364
rect 108908 5352 108914 5364
rect 108945 5355 109003 5361
rect 108945 5352 108957 5355
rect 108908 5324 108957 5352
rect 108908 5312 108914 5324
rect 108945 5321 108957 5324
rect 108991 5321 109003 5355
rect 108945 5315 109003 5321
rect 113177 5355 113235 5361
rect 113177 5321 113189 5355
rect 113223 5352 113235 5355
rect 115198 5352 115204 5364
rect 113223 5324 115204 5352
rect 113223 5321 113235 5324
rect 113177 5315 113235 5321
rect 115198 5312 115204 5324
rect 115256 5312 115262 5364
rect 116029 5355 116087 5361
rect 116029 5321 116041 5355
rect 116075 5321 116087 5355
rect 117314 5352 117320 5364
rect 116029 5315 116087 5321
rect 116136 5324 117320 5352
rect 108022 5284 108028 5296
rect 105004 5256 108028 5284
rect 105004 5225 105032 5256
rect 108022 5244 108028 5256
rect 108080 5244 108086 5296
rect 110966 5244 110972 5296
rect 111024 5244 111030 5296
rect 112625 5287 112683 5293
rect 112625 5253 112637 5287
rect 112671 5284 112683 5287
rect 113542 5284 113548 5296
rect 112671 5256 113548 5284
rect 112671 5253 112683 5256
rect 112625 5247 112683 5253
rect 113542 5244 113548 5256
rect 113600 5244 113606 5296
rect 113726 5244 113732 5296
rect 113784 5284 113790 5296
rect 114278 5284 114284 5296
rect 113784 5256 114284 5284
rect 113784 5244 113790 5256
rect 114278 5244 114284 5256
rect 114336 5284 114342 5296
rect 114336 5256 114876 5284
rect 114336 5244 114342 5256
rect 103333 5219 103391 5225
rect 103333 5216 103345 5219
rect 102704 5188 103345 5216
rect 103333 5185 103345 5188
rect 103379 5185 103391 5219
rect 103333 5179 103391 5185
rect 104989 5219 105047 5225
rect 104989 5185 105001 5219
rect 105035 5185 105047 5219
rect 104989 5179 105047 5185
rect 105725 5219 105783 5225
rect 105725 5185 105737 5219
rect 105771 5185 105783 5219
rect 105725 5179 105783 5185
rect 105265 5151 105323 5157
rect 105265 5148 105277 5151
rect 102612 5120 105277 5148
rect 105265 5117 105277 5120
rect 105311 5148 105323 5151
rect 105740 5148 105768 5179
rect 107010 5176 107016 5228
rect 107068 5216 107074 5228
rect 107654 5216 107660 5228
rect 107068 5188 107660 5216
rect 107068 5176 107074 5188
rect 107654 5176 107660 5188
rect 107712 5176 107718 5228
rect 108574 5176 108580 5228
rect 108632 5176 108638 5228
rect 108666 5176 108672 5228
rect 108724 5176 108730 5228
rect 109773 5219 109831 5225
rect 109773 5185 109785 5219
rect 109819 5185 109831 5219
rect 109773 5179 109831 5185
rect 110141 5219 110199 5225
rect 110141 5185 110153 5219
rect 110187 5216 110199 5219
rect 110506 5216 110512 5228
rect 110187 5188 110512 5216
rect 110187 5185 110199 5188
rect 110141 5179 110199 5185
rect 105814 5148 105820 5160
rect 105311 5120 105820 5148
rect 105311 5117 105323 5120
rect 105265 5111 105323 5117
rect 105814 5108 105820 5120
rect 105872 5108 105878 5160
rect 107194 5108 107200 5160
rect 107252 5148 107258 5160
rect 107289 5151 107347 5157
rect 107289 5148 107301 5151
rect 107252 5120 107301 5148
rect 107252 5108 107258 5120
rect 107289 5117 107301 5120
rect 107335 5117 107347 5151
rect 109788 5148 109816 5179
rect 110506 5176 110512 5188
rect 110564 5176 110570 5228
rect 110782 5176 110788 5228
rect 110840 5176 110846 5228
rect 113361 5220 113419 5225
rect 113361 5219 113496 5220
rect 113361 5185 113373 5219
rect 113407 5192 113496 5219
rect 113407 5185 113419 5192
rect 113361 5179 113419 5185
rect 110230 5148 110236 5160
rect 109788 5120 110236 5148
rect 107289 5111 107347 5117
rect 110230 5108 110236 5120
rect 110288 5108 110294 5160
rect 96890 5080 96896 5092
rect 96172 5052 96896 5080
rect 96890 5040 96896 5052
rect 96948 5080 96954 5092
rect 99834 5080 99840 5092
rect 96948 5052 99840 5080
rect 96948 5040 96954 5052
rect 99834 5040 99840 5052
rect 99892 5040 99898 5092
rect 100018 5040 100024 5092
rect 100076 5080 100082 5092
rect 111426 5080 111432 5092
rect 100076 5052 111432 5080
rect 100076 5040 100082 5052
rect 111426 5040 111432 5052
rect 111484 5040 111490 5092
rect 113468 5080 113496 5192
rect 113821 5219 113879 5225
rect 113821 5185 113833 5219
rect 113867 5216 113879 5219
rect 114186 5216 114192 5228
rect 113867 5188 114192 5216
rect 113867 5185 113879 5188
rect 113821 5179 113879 5185
rect 114186 5176 114192 5188
rect 114244 5216 114250 5228
rect 114848 5225 114876 5256
rect 114922 5244 114928 5296
rect 114980 5284 114986 5296
rect 116044 5284 116072 5315
rect 114980 5256 116072 5284
rect 114980 5244 114986 5256
rect 114741 5219 114799 5225
rect 114741 5216 114753 5219
rect 114244 5188 114753 5216
rect 114244 5176 114250 5188
rect 114741 5185 114753 5188
rect 114787 5185 114799 5219
rect 114741 5179 114799 5185
rect 114833 5219 114891 5225
rect 114833 5185 114845 5219
rect 114879 5185 114891 5219
rect 114833 5179 114891 5185
rect 115845 5219 115903 5225
rect 115845 5185 115857 5219
rect 115891 5216 115903 5219
rect 116136 5216 116164 5324
rect 117314 5312 117320 5324
rect 117372 5312 117378 5364
rect 122466 5312 122472 5364
rect 122524 5352 122530 5364
rect 143721 5355 143779 5361
rect 122524 5324 143580 5352
rect 122524 5312 122530 5324
rect 117498 5284 117504 5296
rect 116228 5256 116440 5284
rect 116228 5228 116256 5256
rect 115891 5188 116164 5216
rect 115891 5185 115903 5188
rect 115845 5179 115903 5185
rect 113726 5108 113732 5160
rect 113784 5148 113790 5160
rect 113913 5151 113971 5157
rect 113913 5148 113925 5151
rect 113784 5120 113925 5148
rect 113784 5108 113790 5120
rect 113913 5117 113925 5120
rect 113959 5117 113971 5151
rect 114756 5148 114784 5179
rect 116210 5176 116216 5228
rect 116268 5176 116274 5228
rect 116026 5148 116032 5160
rect 114756 5120 116032 5148
rect 113913 5111 113971 5117
rect 116026 5108 116032 5120
rect 116084 5108 116090 5160
rect 116412 5148 116440 5256
rect 116504 5256 117504 5284
rect 116504 5225 116532 5256
rect 117498 5244 117504 5256
rect 117556 5244 117562 5296
rect 117590 5244 117596 5296
rect 117648 5284 117654 5296
rect 143442 5284 143448 5296
rect 117648 5256 143448 5284
rect 117648 5244 117654 5256
rect 143442 5244 143448 5256
rect 143500 5244 143506 5296
rect 116489 5219 116547 5225
rect 116489 5185 116501 5219
rect 116535 5185 116547 5219
rect 116489 5179 116547 5185
rect 116946 5176 116952 5228
rect 117004 5176 117010 5228
rect 118789 5219 118847 5225
rect 118789 5185 118801 5219
rect 118835 5216 118847 5219
rect 119246 5216 119252 5228
rect 118835 5188 119252 5216
rect 118835 5185 118847 5188
rect 118789 5179 118847 5185
rect 119246 5176 119252 5188
rect 119304 5176 119310 5228
rect 119893 5219 119951 5225
rect 119893 5185 119905 5219
rect 119939 5216 119951 5219
rect 119982 5216 119988 5228
rect 119939 5188 119988 5216
rect 119939 5185 119951 5188
rect 119893 5179 119951 5185
rect 119982 5176 119988 5188
rect 120040 5176 120046 5228
rect 120629 5219 120687 5225
rect 120629 5185 120641 5219
rect 120675 5185 120687 5219
rect 120629 5179 120687 5185
rect 116670 5148 116676 5160
rect 116412 5120 116676 5148
rect 116670 5108 116676 5120
rect 116728 5108 116734 5160
rect 117133 5151 117191 5157
rect 117133 5117 117145 5151
rect 117179 5148 117191 5151
rect 117406 5148 117412 5160
rect 117179 5120 117412 5148
rect 117179 5117 117191 5120
rect 117133 5111 117191 5117
rect 117406 5108 117412 5120
rect 117464 5108 117470 5160
rect 120644 5148 120672 5179
rect 120994 5176 121000 5228
rect 121052 5176 121058 5228
rect 121822 5176 121828 5228
rect 121880 5176 121886 5228
rect 121914 5176 121920 5228
rect 121972 5216 121978 5228
rect 122469 5219 122527 5225
rect 122469 5216 122481 5219
rect 121972 5188 122481 5216
rect 121972 5176 121978 5188
rect 122469 5185 122481 5188
rect 122515 5185 122527 5219
rect 122469 5179 122527 5185
rect 137462 5176 137468 5228
rect 137520 5176 137526 5228
rect 138750 5176 138756 5228
rect 138808 5176 138814 5228
rect 139394 5176 139400 5228
rect 139452 5216 139458 5228
rect 139452 5188 140268 5216
rect 139452 5176 139458 5188
rect 121270 5148 121276 5160
rect 120644 5120 121276 5148
rect 121270 5108 121276 5120
rect 121328 5108 121334 5160
rect 122742 5108 122748 5160
rect 122800 5148 122806 5160
rect 137741 5151 137799 5157
rect 122800 5120 137692 5148
rect 122800 5108 122806 5120
rect 114462 5080 114468 5092
rect 113468 5052 114468 5080
rect 114462 5040 114468 5052
rect 114520 5040 114526 5092
rect 115106 5040 115112 5092
rect 115164 5040 115170 5092
rect 120166 5040 120172 5092
rect 120224 5080 120230 5092
rect 121181 5083 121239 5089
rect 121181 5080 121193 5083
rect 120224 5052 121193 5080
rect 120224 5040 120230 5052
rect 121181 5049 121193 5052
rect 121227 5049 121239 5083
rect 121181 5043 121239 5049
rect 122374 5040 122380 5092
rect 122432 5080 122438 5092
rect 137278 5080 137284 5092
rect 122432 5052 137284 5080
rect 122432 5040 122438 5052
rect 137278 5040 137284 5052
rect 137336 5040 137342 5092
rect 12066 4972 12072 5024
rect 12124 5012 12130 5024
rect 35526 5012 35532 5024
rect 12124 4984 35532 5012
rect 12124 4972 12130 4984
rect 35526 4972 35532 4984
rect 35584 4972 35590 5024
rect 36814 4972 36820 5024
rect 36872 4972 36878 5024
rect 36906 4972 36912 5024
rect 36964 5012 36970 5024
rect 42610 5012 42616 5024
rect 36964 4984 42616 5012
rect 36964 4972 36970 4984
rect 42610 4972 42616 4984
rect 42668 4972 42674 5024
rect 92290 4972 92296 5024
rect 92348 5012 92354 5024
rect 93302 5012 93308 5024
rect 92348 4984 93308 5012
rect 92348 4972 92354 4984
rect 93302 4972 93308 4984
rect 93360 4972 93366 5024
rect 93397 5015 93455 5021
rect 93397 4981 93409 5015
rect 93443 5012 93455 5015
rect 94498 5012 94504 5024
rect 93443 4984 94504 5012
rect 93443 4981 93455 4984
rect 93397 4975 93455 4981
rect 94498 4972 94504 4984
rect 94556 4972 94562 5024
rect 94682 4972 94688 5024
rect 94740 5012 94746 5024
rect 99190 5012 99196 5024
rect 94740 4984 99196 5012
rect 94740 4972 94746 4984
rect 99190 4972 99196 4984
rect 99248 4972 99254 5024
rect 99653 5015 99711 5021
rect 99653 4981 99665 5015
rect 99699 5012 99711 5015
rect 100110 5012 100116 5024
rect 99699 4984 100116 5012
rect 99699 4981 99711 4984
rect 99653 4975 99711 4981
rect 100110 4972 100116 4984
rect 100168 4972 100174 5024
rect 100386 4972 100392 5024
rect 100444 5012 100450 5024
rect 101398 5012 101404 5024
rect 100444 4984 101404 5012
rect 100444 4972 100450 4984
rect 101398 4972 101404 4984
rect 101456 4972 101462 5024
rect 101766 4972 101772 5024
rect 101824 5012 101830 5024
rect 102321 5015 102379 5021
rect 102321 5012 102333 5015
rect 101824 4984 102333 5012
rect 101824 4972 101830 4984
rect 102321 4981 102333 4984
rect 102367 4981 102379 5015
rect 102321 4975 102379 4981
rect 103146 4972 103152 5024
rect 103204 4972 103210 5024
rect 103238 4972 103244 5024
rect 103296 5012 103302 5024
rect 104805 5015 104863 5021
rect 104805 5012 104817 5015
rect 103296 4984 104817 5012
rect 103296 4972 103302 4984
rect 104805 4981 104817 4984
rect 104851 4981 104863 5015
rect 104805 4975 104863 4981
rect 105722 4972 105728 5024
rect 105780 5012 105786 5024
rect 105817 5015 105875 5021
rect 105817 5012 105829 5015
rect 105780 4984 105829 5012
rect 105780 4972 105786 4984
rect 105817 4981 105829 4984
rect 105863 4981 105875 5015
rect 105817 4975 105875 4981
rect 105998 4972 106004 5024
rect 106056 5012 106062 5024
rect 106918 5012 106924 5024
rect 106056 4984 106924 5012
rect 106056 4972 106062 4984
rect 106918 4972 106924 4984
rect 106976 4972 106982 5024
rect 108758 4972 108764 5024
rect 108816 4972 108822 5024
rect 109770 4972 109776 5024
rect 109828 5012 109834 5024
rect 109865 5015 109923 5021
rect 109865 5012 109877 5015
rect 109828 4984 109877 5012
rect 109828 4972 109834 4984
rect 109865 4981 109877 4984
rect 109911 4981 109923 5015
rect 109865 4975 109923 4981
rect 109954 4972 109960 5024
rect 110012 5012 110018 5024
rect 110325 5015 110383 5021
rect 110325 5012 110337 5015
rect 110012 4984 110337 5012
rect 110012 4972 110018 4984
rect 110325 4981 110337 4984
rect 110371 4981 110383 5015
rect 110325 4975 110383 4981
rect 113358 4972 113364 5024
rect 113416 5012 113422 5024
rect 113821 5015 113879 5021
rect 113821 5012 113833 5015
rect 113416 4984 113833 5012
rect 113416 4972 113422 4984
rect 113821 4981 113833 4984
rect 113867 5012 113879 5015
rect 114002 5012 114008 5024
rect 113867 4984 114008 5012
rect 113867 4981 113879 4984
rect 113821 4975 113879 4981
rect 114002 4972 114008 4984
rect 114060 4972 114066 5024
rect 114186 4972 114192 5024
rect 114244 4972 114250 5024
rect 114370 4972 114376 5024
rect 114428 5012 114434 5024
rect 114741 5015 114799 5021
rect 114741 5012 114753 5015
rect 114428 4984 114753 5012
rect 114428 4972 114434 4984
rect 114741 4981 114753 4984
rect 114787 5012 114799 5015
rect 116026 5012 116032 5024
rect 114787 4984 116032 5012
rect 114787 4981 114799 4984
rect 114741 4975 114799 4981
rect 116026 4972 116032 4984
rect 116084 4972 116090 5024
rect 116302 4972 116308 5024
rect 116360 4972 116366 5024
rect 117130 4972 117136 5024
rect 117188 5012 117194 5024
rect 118142 5012 118148 5024
rect 117188 4984 118148 5012
rect 117188 4972 117194 4984
rect 118142 4972 118148 4984
rect 118200 4972 118206 5024
rect 120077 5015 120135 5021
rect 120077 4981 120089 5015
rect 120123 5012 120135 5015
rect 120902 5012 120908 5024
rect 120123 4984 120908 5012
rect 120123 4981 120135 4984
rect 120077 4975 120135 4981
rect 120902 4972 120908 4984
rect 120960 4972 120966 5024
rect 121638 4972 121644 5024
rect 121696 4972 121702 5024
rect 122282 4972 122288 5024
rect 122340 4972 122346 5024
rect 135898 4972 135904 5024
rect 135956 5012 135962 5024
rect 137557 5015 137615 5021
rect 137557 5012 137569 5015
rect 135956 4984 137569 5012
rect 135956 4972 135962 4984
rect 137557 4981 137569 4984
rect 137603 4981 137615 5015
rect 137664 5012 137692 5120
rect 137741 5117 137753 5151
rect 137787 5148 137799 5151
rect 139578 5148 139584 5160
rect 137787 5120 138612 5148
rect 137787 5117 137799 5120
rect 137741 5111 137799 5117
rect 138017 5083 138075 5089
rect 138017 5049 138029 5083
rect 138063 5080 138075 5083
rect 138106 5080 138112 5092
rect 138063 5052 138112 5080
rect 138063 5049 138075 5052
rect 138017 5043 138075 5049
rect 138106 5040 138112 5052
rect 138164 5040 138170 5092
rect 138584 5080 138612 5120
rect 139320 5120 139584 5148
rect 138937 5083 138995 5089
rect 138937 5080 138949 5083
rect 138584 5052 138949 5080
rect 138937 5049 138949 5052
rect 138983 5080 138995 5083
rect 139026 5080 139032 5092
rect 138983 5052 139032 5080
rect 138983 5049 138995 5052
rect 138937 5043 138995 5049
rect 139026 5040 139032 5052
rect 139084 5040 139090 5092
rect 139320 5012 139348 5120
rect 139578 5108 139584 5120
rect 139636 5108 139642 5160
rect 139673 5151 139731 5157
rect 139673 5117 139685 5151
rect 139719 5148 139731 5151
rect 139762 5148 139768 5160
rect 139719 5120 139768 5148
rect 139719 5117 139731 5120
rect 139673 5111 139731 5117
rect 139762 5108 139768 5120
rect 139820 5148 139826 5160
rect 140240 5148 140268 5188
rect 140314 5176 140320 5228
rect 140372 5216 140378 5228
rect 140501 5219 140559 5225
rect 140501 5216 140513 5219
rect 140372 5188 140513 5216
rect 140372 5176 140378 5188
rect 140501 5185 140513 5188
rect 140547 5185 140559 5219
rect 141878 5216 141884 5228
rect 140501 5179 140559 5185
rect 140792 5188 141884 5216
rect 140792 5157 140820 5188
rect 141878 5176 141884 5188
rect 141936 5216 141942 5228
rect 142157 5219 142215 5225
rect 142157 5216 142169 5219
rect 141936 5188 142169 5216
rect 141936 5176 141942 5188
rect 142157 5185 142169 5188
rect 142203 5216 142215 5219
rect 143169 5219 143227 5225
rect 143169 5216 143181 5219
rect 142203 5188 143181 5216
rect 142203 5185 142215 5188
rect 142157 5179 142215 5185
rect 143169 5185 143181 5188
rect 143215 5185 143227 5219
rect 143169 5179 143227 5185
rect 140777 5151 140835 5157
rect 140777 5148 140789 5151
rect 139820 5120 140176 5148
rect 140240 5120 140789 5148
rect 139820 5108 139826 5120
rect 139949 5083 140007 5089
rect 139949 5049 139961 5083
rect 139995 5080 140007 5083
rect 140038 5080 140044 5092
rect 139995 5052 140044 5080
rect 139995 5049 140007 5052
rect 139949 5043 140007 5049
rect 140038 5040 140044 5052
rect 140096 5040 140102 5092
rect 140148 5080 140176 5120
rect 140777 5117 140789 5120
rect 140823 5117 140835 5151
rect 140777 5111 140835 5117
rect 142433 5151 142491 5157
rect 142433 5117 142445 5151
rect 142479 5148 142491 5151
rect 143445 5151 143503 5157
rect 143445 5148 143457 5151
rect 142479 5120 143457 5148
rect 142479 5117 142491 5120
rect 142433 5111 142491 5117
rect 143445 5117 143457 5120
rect 143491 5117 143503 5151
rect 143552 5148 143580 5324
rect 143721 5321 143733 5355
rect 143767 5321 143779 5355
rect 143721 5315 143779 5321
rect 143736 5284 143764 5315
rect 145558 5312 145564 5364
rect 145616 5352 145622 5364
rect 165614 5352 165620 5364
rect 145616 5324 165620 5352
rect 145616 5312 145622 5324
rect 165614 5312 165620 5324
rect 165672 5312 165678 5364
rect 166966 5324 167868 5352
rect 147490 5284 147496 5296
rect 143736 5256 145052 5284
rect 143626 5176 143632 5228
rect 143684 5216 143690 5228
rect 145024 5225 145052 5256
rect 145668 5256 147496 5284
rect 145668 5225 145696 5256
rect 147490 5244 147496 5256
rect 147548 5244 147554 5296
rect 150618 5284 150624 5296
rect 150452 5256 150624 5284
rect 144365 5219 144423 5225
rect 144365 5216 144377 5219
rect 143684 5188 144377 5216
rect 143684 5176 143690 5188
rect 144365 5185 144377 5188
rect 144411 5185 144423 5219
rect 144365 5179 144423 5185
rect 145009 5219 145067 5225
rect 145009 5185 145021 5219
rect 145055 5185 145067 5219
rect 145009 5179 145067 5185
rect 145653 5219 145711 5225
rect 145653 5185 145665 5219
rect 145699 5185 145711 5219
rect 145653 5179 145711 5185
rect 148134 5176 148140 5228
rect 148192 5216 148198 5228
rect 148229 5219 148287 5225
rect 148229 5216 148241 5219
rect 148192 5188 148241 5216
rect 148192 5176 148198 5188
rect 148229 5185 148241 5188
rect 148275 5185 148287 5219
rect 148229 5179 148287 5185
rect 148502 5176 148508 5228
rect 148560 5176 148566 5228
rect 149698 5176 149704 5228
rect 149756 5225 149762 5228
rect 149756 5216 149764 5225
rect 150452 5216 150480 5256
rect 150618 5244 150624 5256
rect 150676 5244 150682 5296
rect 152642 5244 152648 5296
rect 152700 5284 152706 5296
rect 153289 5287 153347 5293
rect 153289 5284 153301 5287
rect 152700 5256 153301 5284
rect 152700 5244 152706 5256
rect 153289 5253 153301 5256
rect 153335 5253 153347 5287
rect 153289 5247 153347 5253
rect 153378 5244 153384 5296
rect 153436 5284 153442 5296
rect 156141 5287 156199 5293
rect 156141 5284 156153 5287
rect 153436 5256 156153 5284
rect 153436 5244 153442 5256
rect 156141 5253 156153 5256
rect 156187 5253 156199 5287
rect 156141 5247 156199 5253
rect 156414 5244 156420 5296
rect 156472 5284 156478 5296
rect 166966 5284 166994 5324
rect 156472 5256 166994 5284
rect 156472 5244 156478 5256
rect 149756 5188 150480 5216
rect 149756 5179 149764 5188
rect 149756 5176 149762 5179
rect 150526 5176 150532 5228
rect 150584 5216 150590 5228
rect 150805 5219 150863 5225
rect 150805 5216 150817 5219
rect 150584 5188 150817 5216
rect 150584 5176 150590 5188
rect 150805 5185 150817 5188
rect 150851 5185 150863 5219
rect 150805 5179 150863 5185
rect 145558 5148 145564 5160
rect 143552 5120 145564 5148
rect 143445 5111 143503 5117
rect 142448 5080 142476 5111
rect 145558 5108 145564 5120
rect 145616 5108 145622 5160
rect 145837 5151 145895 5157
rect 145837 5117 145849 5151
rect 145883 5117 145895 5151
rect 145837 5111 145895 5117
rect 142522 5080 142528 5092
rect 140148 5052 142528 5080
rect 142522 5040 142528 5052
rect 142580 5040 142586 5092
rect 144181 5083 144239 5089
rect 144181 5049 144193 5083
rect 144227 5080 144239 5083
rect 145852 5080 145880 5111
rect 146386 5108 146392 5160
rect 146444 5108 146450 5160
rect 148520 5148 148548 5176
rect 151722 5174 151728 5226
rect 151780 5214 151786 5226
rect 152734 5216 152740 5228
rect 151780 5186 151823 5214
rect 152568 5188 152740 5216
rect 151780 5174 151786 5186
rect 149977 5151 150035 5157
rect 149977 5148 149989 5151
rect 148520 5120 149989 5148
rect 149977 5117 149989 5120
rect 150023 5117 150035 5151
rect 149977 5111 150035 5117
rect 150986 5108 150992 5160
rect 151044 5108 151050 5160
rect 151906 5157 151912 5160
rect 151863 5151 151912 5157
rect 151863 5117 151875 5151
rect 151909 5117 151912 5151
rect 151863 5111 151912 5117
rect 151906 5108 151912 5111
rect 151964 5108 151970 5160
rect 152001 5151 152059 5157
rect 152001 5117 152013 5151
rect 152047 5148 152059 5151
rect 152568 5148 152596 5188
rect 152734 5176 152740 5188
rect 152792 5176 152798 5228
rect 155954 5176 155960 5228
rect 156012 5176 156018 5228
rect 159726 5176 159732 5228
rect 159784 5216 159790 5228
rect 167454 5216 167460 5228
rect 159784 5188 167460 5216
rect 159784 5176 159790 5188
rect 167454 5176 167460 5188
rect 167512 5176 167518 5228
rect 167840 5216 167868 5324
rect 167914 5312 167920 5364
rect 167972 5352 167978 5364
rect 171042 5352 171048 5364
rect 167972 5324 171048 5352
rect 167972 5312 167978 5324
rect 171042 5312 171048 5324
rect 171100 5312 171106 5364
rect 206738 5352 206744 5364
rect 195946 5324 206744 5352
rect 195946 5284 195974 5324
rect 206738 5312 206744 5324
rect 206796 5312 206802 5364
rect 206925 5355 206983 5361
rect 206925 5321 206937 5355
rect 206971 5352 206983 5355
rect 207474 5352 207480 5364
rect 206971 5324 207480 5352
rect 206971 5321 206983 5324
rect 206925 5315 206983 5321
rect 207474 5312 207480 5324
rect 207532 5312 207538 5364
rect 207584 5324 209912 5352
rect 207584 5284 207612 5324
rect 168116 5256 195974 5284
rect 206756 5256 207612 5284
rect 168116 5216 168144 5256
rect 167840 5188 168144 5216
rect 169570 5176 169576 5228
rect 169628 5216 169634 5228
rect 169941 5219 169999 5225
rect 169941 5216 169953 5219
rect 169628 5188 169953 5216
rect 169628 5176 169634 5188
rect 169941 5185 169953 5188
rect 169987 5185 169999 5219
rect 169941 5179 169999 5185
rect 205634 5176 205640 5228
rect 205692 5216 205698 5228
rect 206557 5219 206615 5225
rect 206557 5216 206569 5219
rect 205692 5188 206569 5216
rect 205692 5176 205698 5188
rect 206557 5185 206569 5188
rect 206603 5185 206615 5219
rect 206557 5179 206615 5185
rect 206646 5176 206652 5228
rect 206704 5176 206710 5228
rect 206756 5225 206784 5256
rect 206741 5219 206799 5225
rect 206741 5185 206753 5219
rect 206787 5185 206799 5219
rect 206741 5179 206799 5185
rect 153105 5151 153163 5157
rect 153105 5148 153117 5151
rect 152047 5120 152596 5148
rect 152844 5120 153117 5148
rect 152047 5117 152059 5120
rect 152001 5111 152059 5117
rect 144227 5052 145880 5080
rect 144227 5049 144239 5052
rect 144181 5043 144239 5049
rect 148134 5040 148140 5092
rect 148192 5080 148198 5092
rect 148192 5052 148456 5080
rect 148192 5040 148198 5052
rect 137664 4984 139348 5012
rect 137557 4975 137615 4981
rect 139486 4972 139492 5024
rect 139544 4972 139550 5024
rect 142246 4972 142252 5024
rect 142304 4972 142310 5024
rect 142706 4972 142712 5024
rect 142764 4972 142770 5024
rect 143442 4972 143448 5024
rect 143500 4972 143506 5024
rect 144825 5015 144883 5021
rect 144825 4981 144837 5015
rect 144871 5012 144883 5015
rect 145650 5012 145656 5024
rect 144871 4984 145656 5012
rect 144871 4981 144883 4984
rect 144825 4975 144883 4981
rect 145650 4972 145656 4984
rect 145708 4972 145714 5024
rect 148318 4972 148324 5024
rect 148376 4972 148382 5024
rect 148428 5012 148456 5052
rect 148778 5040 148784 5092
rect 148836 5040 148842 5092
rect 150253 5083 150311 5089
rect 148888 5052 149928 5080
rect 148888 5012 148916 5052
rect 148428 4984 148916 5012
rect 149238 4972 149244 5024
rect 149296 5012 149302 5024
rect 149790 5012 149796 5024
rect 149296 4984 149796 5012
rect 149296 4972 149302 4984
rect 149790 4972 149796 4984
rect 149848 4972 149854 5024
rect 149900 5012 149928 5052
rect 150253 5049 150265 5083
rect 150299 5080 150311 5083
rect 150434 5080 150440 5092
rect 150299 5052 150440 5080
rect 150299 5049 150311 5052
rect 150253 5043 150311 5049
rect 150434 5040 150440 5052
rect 150492 5040 150498 5092
rect 150618 5040 150624 5092
rect 150676 5080 150682 5092
rect 151262 5080 151268 5092
rect 150676 5052 151268 5080
rect 150676 5040 150682 5052
rect 151262 5040 151268 5052
rect 151320 5040 151326 5092
rect 151446 5040 151452 5092
rect 151504 5040 151510 5092
rect 150342 5012 150348 5024
rect 149900 4984 150348 5012
rect 150342 4972 150348 4984
rect 150400 5012 150406 5024
rect 152384 5012 152412 5120
rect 152844 5080 152872 5120
rect 153105 5117 153117 5120
rect 153151 5117 153163 5151
rect 153105 5111 153163 5117
rect 154758 5108 154764 5160
rect 154816 5108 154822 5160
rect 154942 5108 154948 5160
rect 155000 5148 155006 5160
rect 156874 5148 156880 5160
rect 155000 5120 156880 5148
rect 155000 5108 155006 5120
rect 156874 5108 156880 5120
rect 156932 5108 156938 5160
rect 157794 5108 157800 5160
rect 157852 5148 157858 5160
rect 167914 5148 167920 5160
rect 157852 5120 167920 5148
rect 157852 5108 157858 5120
rect 167914 5108 167920 5120
rect 167972 5108 167978 5160
rect 168098 5108 168104 5160
rect 168156 5108 168162 5160
rect 168282 5108 168288 5160
rect 168340 5148 168346 5160
rect 169846 5148 169852 5160
rect 168340 5120 169852 5148
rect 168340 5108 168346 5120
rect 169846 5108 169852 5120
rect 169904 5108 169910 5160
rect 205818 5108 205824 5160
rect 205876 5148 205882 5160
rect 206756 5148 206784 5179
rect 206830 5176 206836 5228
rect 206888 5216 206894 5228
rect 209884 5225 209912 5324
rect 214098 5312 214104 5364
rect 214156 5352 214162 5364
rect 217134 5352 217140 5364
rect 214156 5324 217140 5352
rect 214156 5312 214162 5324
rect 217134 5312 217140 5324
rect 217192 5312 217198 5364
rect 219894 5352 219900 5364
rect 218072 5324 219900 5352
rect 216122 5284 216128 5296
rect 215220 5256 216128 5284
rect 207477 5219 207535 5225
rect 207477 5216 207489 5219
rect 206888 5188 207489 5216
rect 206888 5176 206894 5188
rect 207477 5185 207489 5188
rect 207523 5185 207535 5219
rect 207477 5179 207535 5185
rect 209869 5219 209927 5225
rect 209869 5185 209881 5219
rect 209915 5216 209927 5219
rect 210326 5216 210332 5228
rect 209915 5188 210332 5216
rect 209915 5185 209927 5188
rect 209869 5179 209927 5185
rect 210326 5176 210332 5188
rect 210384 5176 210390 5228
rect 213178 5176 213184 5228
rect 213236 5176 213242 5228
rect 213270 5176 213276 5228
rect 213328 5216 213334 5228
rect 213457 5219 213515 5225
rect 213457 5216 213469 5219
rect 213328 5188 213469 5216
rect 213328 5176 213334 5188
rect 213457 5185 213469 5188
rect 213503 5185 213515 5219
rect 213457 5179 213515 5185
rect 214374 5176 214380 5228
rect 214432 5176 214438 5228
rect 214466 5176 214472 5228
rect 214524 5225 214530 5228
rect 214524 5219 214552 5225
rect 214540 5185 214552 5219
rect 214524 5179 214552 5185
rect 214524 5176 214530 5179
rect 205876 5120 206784 5148
rect 205876 5108 205882 5120
rect 207106 5108 207112 5160
rect 207164 5148 207170 5160
rect 207661 5151 207719 5157
rect 207661 5148 207673 5151
rect 207164 5120 207673 5148
rect 207164 5108 207170 5120
rect 207661 5117 207673 5120
rect 207707 5117 207719 5151
rect 207661 5111 207719 5117
rect 208394 5108 208400 5160
rect 208452 5108 208458 5160
rect 208578 5157 208584 5160
rect 208535 5151 208584 5157
rect 208535 5117 208547 5151
rect 208581 5117 208584 5151
rect 208535 5111 208584 5117
rect 208578 5108 208584 5111
rect 208636 5108 208642 5160
rect 208673 5151 208731 5157
rect 208673 5117 208685 5151
rect 208719 5148 208731 5151
rect 209222 5148 209228 5160
rect 208719 5120 209228 5148
rect 208719 5117 208731 5120
rect 208673 5111 208731 5117
rect 209222 5108 209228 5120
rect 209280 5108 209286 5160
rect 213546 5108 213552 5160
rect 213604 5148 213610 5160
rect 213641 5151 213699 5157
rect 213641 5148 213653 5151
rect 213604 5120 213653 5148
rect 213604 5108 213610 5120
rect 213641 5117 213653 5120
rect 213687 5117 213699 5151
rect 213641 5111 213699 5117
rect 214098 5108 214104 5160
rect 214156 5108 214162 5160
rect 214653 5151 214711 5157
rect 214653 5148 214665 5151
rect 214208 5120 214665 5148
rect 152660 5052 152872 5080
rect 152660 5021 152688 5052
rect 152918 5040 152924 5092
rect 152976 5080 152982 5092
rect 207566 5080 207572 5092
rect 152976 5052 207572 5080
rect 152976 5040 152982 5052
rect 207566 5040 207572 5052
rect 207624 5040 207630 5092
rect 207750 5040 207756 5092
rect 207808 5080 207814 5092
rect 208121 5083 208179 5089
rect 208121 5080 208133 5083
rect 207808 5052 208133 5080
rect 207808 5040 207814 5052
rect 208121 5049 208133 5052
rect 208167 5049 208179 5083
rect 208121 5043 208179 5049
rect 213454 5040 213460 5092
rect 213512 5080 213518 5092
rect 214116 5080 214144 5108
rect 213512 5052 214144 5080
rect 213512 5040 213518 5052
rect 150400 4984 152412 5012
rect 152645 5015 152703 5021
rect 150400 4972 150406 4984
rect 152645 4981 152657 5015
rect 152691 4981 152703 5015
rect 152645 4975 152703 4981
rect 153286 4972 153292 5024
rect 153344 5012 153350 5024
rect 153930 5012 153936 5024
rect 153344 4984 153936 5012
rect 153344 4972 153350 4984
rect 153930 4972 153936 4984
rect 153988 4972 153994 5024
rect 154022 4972 154028 5024
rect 154080 5012 154086 5024
rect 155310 5012 155316 5024
rect 154080 4984 155316 5012
rect 154080 4972 154086 4984
rect 155310 4972 155316 4984
rect 155368 4972 155374 5024
rect 165614 4972 165620 5024
rect 165672 5012 165678 5024
rect 168282 5012 168288 5024
rect 165672 4984 168288 5012
rect 165672 4972 165678 4984
rect 168282 4972 168288 4984
rect 168340 4972 168346 5024
rect 172514 4972 172520 5024
rect 172572 5012 172578 5024
rect 184566 5012 184572 5024
rect 172572 4984 184572 5012
rect 172572 4972 172578 4984
rect 184566 4972 184572 4984
rect 184624 4972 184630 5024
rect 206462 4972 206468 5024
rect 206520 5012 206526 5024
rect 209317 5015 209375 5021
rect 209317 5012 209329 5015
rect 206520 4984 209329 5012
rect 206520 4972 206526 4984
rect 209317 4981 209329 4984
rect 209363 4981 209375 5015
rect 209317 4975 209375 4981
rect 209958 4972 209964 5024
rect 210016 4972 210022 5024
rect 214006 4972 214012 5024
rect 214064 5012 214070 5024
rect 214208 5012 214236 5120
rect 214653 5117 214665 5120
rect 214699 5148 214711 5151
rect 215220 5148 215248 5256
rect 216122 5244 216128 5256
rect 216180 5244 216186 5296
rect 216490 5244 216496 5296
rect 216548 5244 216554 5296
rect 215570 5176 215576 5228
rect 215628 5216 215634 5228
rect 215849 5219 215907 5225
rect 215849 5216 215861 5219
rect 215628 5188 215861 5216
rect 215628 5176 215634 5188
rect 215849 5185 215861 5188
rect 215895 5185 215907 5219
rect 215849 5179 215907 5185
rect 215938 5176 215944 5228
rect 215996 5176 216002 5228
rect 216306 5176 216312 5228
rect 216364 5176 216370 5228
rect 217134 5176 217140 5228
rect 217192 5176 217198 5228
rect 217778 5176 217784 5228
rect 217836 5216 217842 5228
rect 218072 5225 218100 5324
rect 219894 5312 219900 5324
rect 219952 5312 219958 5364
rect 221366 5352 221372 5364
rect 220004 5324 221372 5352
rect 219710 5244 219716 5296
rect 219768 5284 219774 5296
rect 220004 5284 220032 5324
rect 221366 5312 221372 5324
rect 221424 5312 221430 5364
rect 221476 5324 223252 5352
rect 219768 5256 220032 5284
rect 219768 5244 219774 5256
rect 220078 5244 220084 5296
rect 220136 5284 220142 5296
rect 220357 5287 220415 5293
rect 220357 5284 220369 5287
rect 220136 5256 220369 5284
rect 220136 5244 220142 5256
rect 220357 5253 220369 5256
rect 220403 5253 220415 5287
rect 220357 5247 220415 5253
rect 220630 5244 220636 5296
rect 220688 5284 220694 5296
rect 221476 5284 221504 5324
rect 220688 5256 221504 5284
rect 220688 5244 220694 5256
rect 223114 5244 223120 5296
rect 223172 5244 223178 5296
rect 223224 5284 223252 5324
rect 223758 5312 223764 5364
rect 223816 5352 223822 5364
rect 246206 5352 246212 5364
rect 223816 5324 246212 5352
rect 223816 5312 223822 5324
rect 246206 5312 246212 5324
rect 246264 5312 246270 5364
rect 247221 5355 247279 5361
rect 247221 5321 247233 5355
rect 247267 5352 247279 5355
rect 247267 5324 248092 5352
rect 247267 5321 247279 5324
rect 247221 5315 247279 5321
rect 224954 5284 224960 5296
rect 223224 5256 224960 5284
rect 224954 5244 224960 5256
rect 225012 5244 225018 5296
rect 225417 5287 225475 5293
rect 225417 5284 225429 5287
rect 225064 5256 225429 5284
rect 217873 5219 217931 5225
rect 217873 5216 217885 5219
rect 217836 5188 217885 5216
rect 217836 5176 217842 5188
rect 217873 5185 217885 5188
rect 217919 5185 217931 5219
rect 217873 5179 217931 5185
rect 218057 5219 218115 5225
rect 218057 5185 218069 5219
rect 218103 5185 218115 5219
rect 218057 5179 218115 5185
rect 218790 5176 218796 5228
rect 218848 5176 218854 5228
rect 219069 5219 219127 5225
rect 219069 5185 219081 5219
rect 219115 5185 219127 5219
rect 219069 5179 219127 5185
rect 214699 5120 215248 5148
rect 214699 5117 214711 5120
rect 214653 5111 214711 5117
rect 215386 5108 215392 5160
rect 215444 5148 215450 5160
rect 218422 5148 218428 5160
rect 215444 5120 218428 5148
rect 215444 5108 215450 5120
rect 218422 5108 218428 5120
rect 218480 5108 218486 5160
rect 218517 5151 218575 5157
rect 218517 5117 218529 5151
rect 218563 5148 218575 5151
rect 218606 5148 218612 5160
rect 218563 5120 218612 5148
rect 218563 5117 218575 5120
rect 218517 5111 218575 5117
rect 218606 5108 218612 5120
rect 218664 5108 218670 5160
rect 218974 5157 218980 5160
rect 218931 5151 218980 5157
rect 218931 5117 218943 5151
rect 218977 5117 218980 5151
rect 218931 5111 218980 5117
rect 218974 5108 218980 5111
rect 219032 5108 219038 5160
rect 219084 5148 219112 5179
rect 220170 5176 220176 5228
rect 220228 5176 220234 5228
rect 224402 5176 224408 5228
rect 224460 5216 224466 5228
rect 225064 5216 225092 5256
rect 225417 5253 225429 5256
rect 225463 5253 225475 5287
rect 225417 5247 225475 5253
rect 242986 5244 242992 5296
rect 243044 5284 243050 5296
rect 245010 5284 245016 5296
rect 243044 5256 245016 5284
rect 243044 5244 243050 5256
rect 245010 5244 245016 5256
rect 245068 5244 245074 5296
rect 246574 5244 246580 5296
rect 246632 5284 246638 5296
rect 246761 5287 246819 5293
rect 246761 5284 246773 5287
rect 246632 5256 246773 5284
rect 246632 5244 246638 5256
rect 246761 5253 246773 5256
rect 246807 5284 246819 5287
rect 246942 5284 246948 5296
rect 246807 5256 246948 5284
rect 246807 5253 246819 5256
rect 246761 5247 246819 5253
rect 246942 5244 246948 5256
rect 247000 5244 247006 5296
rect 247678 5244 247684 5296
rect 247736 5244 247742 5296
rect 248064 5284 248092 5324
rect 248138 5312 248144 5364
rect 248196 5312 248202 5364
rect 248800 5324 251956 5352
rect 248800 5284 248828 5324
rect 248064 5256 248828 5284
rect 248874 5244 248880 5296
rect 248932 5244 248938 5296
rect 251085 5287 251143 5293
rect 251085 5253 251097 5287
rect 251131 5284 251143 5287
rect 251726 5284 251732 5296
rect 251131 5256 251732 5284
rect 251131 5253 251143 5256
rect 251085 5247 251143 5253
rect 251726 5244 251732 5256
rect 251784 5244 251790 5296
rect 228634 5216 228640 5228
rect 224460 5188 225092 5216
rect 226628 5188 228640 5216
rect 224460 5176 224466 5188
rect 220722 5148 220728 5160
rect 219084 5120 220728 5148
rect 220722 5108 220728 5120
rect 220780 5108 220786 5160
rect 220814 5108 220820 5160
rect 220872 5108 220878 5160
rect 221734 5108 221740 5160
rect 221792 5148 221798 5160
rect 221792 5120 222884 5148
rect 221792 5108 221798 5120
rect 215110 5040 215116 5092
rect 215168 5080 215174 5092
rect 216306 5080 216312 5092
rect 215168 5052 216312 5080
rect 215168 5040 215174 5052
rect 216306 5040 216312 5052
rect 216364 5040 216370 5092
rect 219526 5040 219532 5092
rect 219584 5080 219590 5092
rect 219584 5052 220124 5080
rect 219584 5040 219590 5052
rect 214064 4984 214236 5012
rect 214064 4972 214070 4984
rect 215294 4972 215300 5024
rect 215352 4972 215358 5024
rect 216950 4972 216956 5024
rect 217008 4972 217014 5024
rect 217962 4972 217968 5024
rect 218020 5012 218026 5024
rect 220096 5021 220124 5052
rect 220906 5040 220912 5092
rect 220964 5080 220970 5092
rect 222378 5080 222384 5092
rect 220964 5052 222384 5080
rect 220964 5040 220970 5052
rect 222378 5040 222384 5052
rect 222436 5040 222442 5092
rect 222856 5080 222884 5120
rect 222930 5108 222936 5160
rect 222988 5108 222994 5160
rect 223758 5108 223764 5160
rect 223816 5148 223822 5160
rect 225138 5148 225144 5160
rect 223816 5120 225144 5148
rect 223816 5108 223822 5120
rect 225138 5108 225144 5120
rect 225196 5108 225202 5160
rect 225230 5108 225236 5160
rect 225288 5108 225294 5160
rect 226628 5148 226656 5188
rect 228634 5176 228640 5188
rect 228692 5176 228698 5228
rect 246117 5219 246175 5225
rect 246117 5185 246129 5219
rect 246163 5216 246175 5219
rect 246666 5216 246672 5228
rect 246163 5188 246672 5216
rect 246163 5185 246175 5188
rect 246117 5179 246175 5185
rect 246666 5176 246672 5188
rect 246724 5176 246730 5228
rect 247034 5176 247040 5228
rect 247092 5176 247098 5228
rect 247218 5176 247224 5228
rect 247276 5216 247282 5228
rect 247862 5216 247868 5228
rect 247276 5188 247868 5216
rect 247276 5176 247282 5188
rect 247862 5176 247868 5188
rect 247920 5176 247926 5228
rect 247957 5219 248015 5225
rect 247957 5185 247969 5219
rect 248003 5185 248015 5219
rect 247957 5179 248015 5185
rect 225984 5120 226656 5148
rect 227073 5151 227131 5157
rect 223482 5080 223488 5092
rect 222856 5052 223488 5080
rect 223482 5040 223488 5052
rect 223540 5040 223546 5092
rect 223574 5040 223580 5092
rect 223632 5080 223638 5092
rect 225984 5080 226012 5120
rect 227073 5117 227085 5151
rect 227119 5148 227131 5151
rect 227438 5148 227444 5160
rect 227119 5120 227444 5148
rect 227119 5117 227131 5120
rect 227073 5111 227131 5117
rect 227438 5108 227444 5120
rect 227496 5108 227502 5160
rect 227622 5108 227628 5160
rect 227680 5148 227686 5160
rect 237282 5148 237288 5160
rect 227680 5120 237288 5148
rect 227680 5108 227686 5120
rect 237282 5108 237288 5120
rect 237340 5108 237346 5160
rect 246850 5108 246856 5160
rect 246908 5108 246914 5160
rect 247972 5148 248000 5179
rect 248690 5176 248696 5228
rect 248748 5176 248754 5228
rect 251928 5225 251956 5324
rect 254486 5312 254492 5364
rect 254544 5352 254550 5364
rect 256418 5352 256424 5364
rect 254544 5324 256424 5352
rect 254544 5312 254550 5324
rect 256418 5312 256424 5324
rect 256476 5312 256482 5364
rect 261570 5312 261576 5364
rect 261628 5352 261634 5364
rect 262306 5352 262312 5364
rect 261628 5324 262312 5352
rect 261628 5312 261634 5324
rect 262306 5312 262312 5324
rect 262364 5312 262370 5364
rect 262490 5312 262496 5364
rect 262548 5312 262554 5364
rect 263413 5355 263471 5361
rect 263413 5321 263425 5355
rect 263459 5352 263471 5355
rect 263686 5352 263692 5364
rect 263459 5324 263692 5352
rect 263459 5321 263471 5324
rect 263413 5315 263471 5321
rect 263686 5312 263692 5324
rect 263744 5312 263750 5364
rect 264974 5312 264980 5364
rect 265032 5352 265038 5364
rect 265069 5355 265127 5361
rect 265069 5352 265081 5355
rect 265032 5324 265081 5352
rect 265032 5312 265038 5324
rect 265069 5321 265081 5324
rect 265115 5321 265127 5355
rect 265069 5315 265127 5321
rect 266538 5312 266544 5364
rect 266596 5352 266602 5364
rect 266817 5355 266875 5361
rect 266817 5352 266829 5355
rect 266596 5324 266829 5352
rect 266596 5312 266602 5324
rect 266817 5321 266829 5324
rect 266863 5321 266875 5355
rect 266817 5315 266875 5321
rect 267734 5312 267740 5364
rect 267792 5312 267798 5364
rect 268378 5312 268384 5364
rect 268436 5352 268442 5364
rect 268565 5355 268623 5361
rect 268565 5352 268577 5355
rect 268436 5324 268577 5352
rect 268436 5312 268442 5324
rect 268565 5321 268577 5324
rect 268611 5321 268623 5355
rect 268565 5315 268623 5321
rect 269390 5312 269396 5364
rect 269448 5352 269454 5364
rect 269669 5355 269727 5361
rect 269669 5352 269681 5355
rect 269448 5324 269681 5352
rect 269448 5312 269454 5324
rect 269669 5321 269681 5324
rect 269715 5321 269727 5355
rect 269669 5315 269727 5321
rect 254118 5244 254124 5296
rect 254176 5284 254182 5296
rect 254213 5287 254271 5293
rect 254213 5284 254225 5287
rect 254176 5256 254225 5284
rect 254176 5244 254182 5256
rect 254213 5253 254225 5256
rect 254259 5284 254271 5287
rect 254259 5256 255084 5284
rect 254259 5253 254271 5256
rect 254213 5247 254271 5253
rect 251913 5219 251971 5225
rect 251913 5185 251925 5219
rect 251959 5185 251971 5219
rect 251913 5179 251971 5185
rect 253293 5219 253351 5225
rect 253293 5185 253305 5219
rect 253339 5185 253351 5219
rect 254489 5219 254547 5225
rect 254489 5216 254501 5219
rect 253293 5179 253351 5185
rect 253906 5188 254501 5216
rect 249150 5148 249156 5160
rect 247972 5120 249156 5148
rect 249150 5108 249156 5120
rect 249208 5108 249214 5160
rect 250533 5151 250591 5157
rect 250533 5117 250545 5151
rect 250579 5148 250591 5151
rect 252646 5148 252652 5160
rect 250579 5120 252652 5148
rect 250579 5117 250591 5120
rect 250533 5111 250591 5117
rect 252646 5108 252652 5120
rect 252704 5108 252710 5160
rect 223632 5052 226012 5080
rect 223632 5040 223638 5052
rect 226058 5040 226064 5092
rect 226116 5080 226122 5092
rect 247034 5080 247040 5092
rect 226116 5052 247040 5080
rect 226116 5040 226122 5052
rect 247034 5040 247040 5052
rect 247092 5040 247098 5092
rect 248322 5040 248328 5092
rect 248380 5080 248386 5092
rect 251266 5080 251272 5092
rect 248380 5052 251272 5080
rect 248380 5040 248386 5052
rect 251266 5040 251272 5052
rect 251324 5040 251330 5092
rect 253308 5080 253336 5179
rect 253906 5160 253934 5188
rect 254489 5185 254501 5188
rect 254535 5216 254547 5219
rect 254670 5216 254676 5228
rect 254535 5188 254676 5216
rect 254535 5185 254547 5188
rect 254489 5179 254547 5185
rect 254670 5176 254676 5188
rect 254728 5176 254734 5228
rect 253842 5108 253848 5160
rect 253900 5120 253934 5160
rect 254397 5151 254455 5157
rect 253900 5108 253906 5120
rect 254397 5117 254409 5151
rect 254443 5148 254455 5151
rect 254578 5148 254584 5160
rect 254443 5120 254584 5148
rect 254443 5117 254455 5120
rect 254397 5111 254455 5117
rect 254578 5108 254584 5120
rect 254636 5108 254642 5160
rect 255056 5148 255084 5256
rect 255314 5244 255320 5296
rect 255372 5244 255378 5296
rect 255406 5244 255412 5296
rect 255464 5284 255470 5296
rect 256973 5287 257031 5293
rect 255464 5256 256556 5284
rect 255464 5244 255470 5256
rect 255130 5176 255136 5228
rect 255188 5176 255194 5228
rect 256528 5216 256556 5256
rect 256973 5253 256985 5287
rect 257019 5284 257031 5287
rect 260282 5284 260288 5296
rect 257019 5256 260288 5284
rect 257019 5253 257031 5256
rect 256973 5247 257031 5253
rect 260282 5244 260288 5256
rect 260340 5244 260346 5296
rect 265805 5287 265863 5293
rect 260944 5256 265388 5284
rect 257338 5216 257344 5228
rect 256528 5188 257344 5216
rect 257338 5176 257344 5188
rect 257396 5216 257402 5228
rect 257433 5219 257491 5225
rect 257433 5216 257445 5219
rect 257396 5188 257445 5216
rect 257396 5176 257402 5188
rect 257433 5185 257445 5188
rect 257479 5185 257491 5219
rect 257433 5179 257491 5185
rect 257614 5176 257620 5228
rect 257672 5216 257678 5228
rect 257709 5219 257767 5225
rect 257709 5216 257721 5219
rect 257672 5188 257721 5216
rect 257672 5176 257678 5188
rect 257709 5185 257721 5188
rect 257755 5216 257767 5219
rect 259362 5216 259368 5228
rect 257755 5188 259368 5216
rect 257755 5185 257767 5188
rect 257709 5179 257767 5185
rect 259362 5176 259368 5188
rect 259420 5176 259426 5228
rect 259825 5219 259883 5225
rect 259825 5185 259837 5219
rect 259871 5216 259883 5219
rect 260944 5216 260972 5256
rect 259871 5188 260972 5216
rect 259871 5185 259883 5188
rect 259825 5179 259883 5185
rect 261018 5176 261024 5228
rect 261076 5176 261082 5228
rect 262306 5176 262312 5228
rect 262364 5176 262370 5228
rect 263594 5176 263600 5228
rect 263652 5176 263658 5228
rect 264606 5176 264612 5228
rect 264664 5176 264670 5228
rect 265250 5176 265256 5228
rect 265308 5176 265314 5228
rect 265360 5216 265388 5256
rect 265805 5253 265817 5287
rect 265851 5284 265863 5287
rect 265986 5284 265992 5296
rect 265851 5256 265992 5284
rect 265851 5253 265863 5256
rect 265805 5247 265863 5253
rect 265986 5244 265992 5256
rect 266044 5284 266050 5296
rect 266044 5256 266676 5284
rect 266044 5244 266050 5256
rect 266446 5216 266452 5228
rect 265360 5188 266452 5216
rect 266446 5176 266452 5188
rect 266504 5176 266510 5228
rect 266538 5176 266544 5228
rect 266596 5176 266602 5228
rect 266648 5225 266676 5256
rect 266906 5244 266912 5296
rect 266964 5284 266970 5296
rect 270497 5287 270555 5293
rect 270497 5284 270509 5287
rect 266964 5256 270509 5284
rect 266964 5244 266970 5256
rect 270497 5253 270509 5256
rect 270543 5253 270555 5287
rect 270497 5247 270555 5253
rect 266633 5219 266691 5225
rect 266633 5185 266645 5219
rect 266679 5216 266691 5219
rect 267274 5216 267280 5228
rect 266679 5188 267280 5216
rect 266679 5185 266691 5188
rect 266633 5179 266691 5185
rect 267274 5176 267280 5188
rect 267332 5176 267338 5228
rect 267461 5219 267519 5225
rect 267461 5185 267473 5219
rect 267507 5185 267519 5219
rect 267461 5179 267519 5185
rect 255406 5148 255412 5160
rect 255056 5120 255412 5148
rect 255406 5108 255412 5120
rect 255464 5108 255470 5160
rect 256694 5108 256700 5160
rect 256752 5148 256758 5160
rect 257522 5148 257528 5160
rect 256752 5120 257528 5148
rect 256752 5108 256758 5120
rect 257522 5108 257528 5120
rect 257580 5148 257586 5160
rect 258718 5148 258724 5160
rect 257580 5120 258724 5148
rect 257580 5108 257586 5120
rect 258718 5108 258724 5120
rect 258776 5108 258782 5160
rect 260098 5108 260104 5160
rect 260156 5108 260162 5160
rect 261386 5108 261392 5160
rect 261444 5108 261450 5160
rect 262125 5151 262183 5157
rect 262125 5117 262137 5151
rect 262171 5148 262183 5151
rect 262582 5148 262588 5160
rect 262171 5120 262588 5148
rect 262171 5117 262183 5120
rect 262125 5111 262183 5117
rect 262582 5108 262588 5120
rect 262640 5108 262646 5160
rect 267476 5148 267504 5179
rect 267550 5176 267556 5228
rect 267608 5216 267614 5228
rect 268286 5216 268292 5228
rect 267608 5188 268292 5216
rect 267608 5176 267614 5188
rect 268286 5176 268292 5188
rect 268344 5216 268350 5228
rect 268381 5219 268439 5225
rect 268381 5216 268393 5219
rect 268344 5188 268393 5216
rect 268344 5176 268350 5188
rect 268381 5185 268393 5188
rect 268427 5185 268439 5219
rect 268381 5179 268439 5185
rect 267826 5148 267832 5160
rect 267476 5120 267832 5148
rect 267826 5108 267832 5120
rect 267884 5108 267890 5160
rect 268194 5108 268200 5160
rect 268252 5108 268258 5160
rect 268396 5148 268424 5179
rect 268470 5176 268476 5228
rect 268528 5216 268534 5228
rect 269301 5219 269359 5225
rect 269301 5216 269313 5219
rect 268528 5188 269313 5216
rect 268528 5176 268534 5188
rect 269301 5185 269313 5188
rect 269347 5185 269359 5219
rect 269301 5179 269359 5185
rect 269485 5219 269543 5225
rect 269485 5185 269497 5219
rect 269531 5185 269543 5219
rect 270313 5219 270371 5225
rect 270313 5216 270325 5219
rect 269485 5179 269543 5185
rect 269868 5188 270325 5216
rect 269500 5148 269528 5179
rect 269868 5160 269896 5188
rect 270313 5185 270325 5188
rect 270359 5185 270371 5219
rect 270313 5179 270371 5185
rect 269850 5148 269856 5160
rect 268396 5120 269856 5148
rect 269850 5108 269856 5120
rect 269908 5108 269914 5160
rect 270129 5151 270187 5157
rect 270129 5117 270141 5151
rect 270175 5117 270187 5151
rect 270129 5111 270187 5117
rect 257893 5083 257951 5089
rect 257893 5080 257905 5083
rect 253308 5052 257905 5080
rect 257893 5049 257905 5052
rect 257939 5049 257951 5083
rect 258626 5080 258632 5092
rect 257893 5043 257951 5049
rect 258000 5052 258632 5080
rect 219713 5015 219771 5021
rect 219713 5012 219725 5015
rect 218020 4984 219725 5012
rect 218020 4972 218026 4984
rect 219713 4981 219725 4984
rect 219759 4981 219771 5015
rect 219713 4975 219771 4981
rect 220081 5015 220139 5021
rect 220081 4981 220093 5015
rect 220127 5012 220139 5015
rect 244918 5012 244924 5024
rect 220127 4984 244924 5012
rect 220127 4981 220139 4984
rect 220081 4975 220139 4981
rect 244918 4972 244924 4984
rect 244976 4972 244982 5024
rect 245102 4972 245108 5024
rect 245160 5012 245166 5024
rect 245933 5015 245991 5021
rect 245933 5012 245945 5015
rect 245160 4984 245945 5012
rect 245160 4972 245166 4984
rect 245933 4981 245945 4984
rect 245979 4981 245991 5015
rect 245933 4975 245991 4981
rect 246942 4972 246948 5024
rect 247000 4972 247006 5024
rect 247957 5015 248015 5021
rect 247957 4981 247969 5015
rect 248003 5012 248015 5015
rect 248782 5012 248788 5024
rect 248003 4984 248788 5012
rect 248003 4981 248015 4984
rect 247957 4975 248015 4981
rect 248782 4972 248788 4984
rect 248840 4972 248846 5024
rect 251174 4972 251180 5024
rect 251232 4972 251238 5024
rect 251726 4972 251732 5024
rect 251784 4972 251790 5024
rect 253109 5015 253167 5021
rect 253109 4981 253121 5015
rect 253155 5012 253167 5015
rect 253934 5012 253940 5024
rect 253155 4984 253940 5012
rect 253155 4981 253167 4984
rect 253109 4975 253167 4981
rect 253934 4972 253940 4984
rect 253992 4972 253998 5024
rect 254486 4972 254492 5024
rect 254544 4972 254550 5024
rect 254673 5015 254731 5021
rect 254673 4981 254685 5015
rect 254719 5012 254731 5015
rect 255866 5012 255872 5024
rect 254719 4984 255872 5012
rect 254719 4981 254731 4984
rect 254673 4975 254731 4981
rect 255866 4972 255872 4984
rect 255924 4972 255930 5024
rect 256418 4972 256424 5024
rect 256476 5012 256482 5024
rect 257709 5015 257767 5021
rect 257709 5012 257721 5015
rect 256476 4984 257721 5012
rect 256476 4972 256482 4984
rect 257709 4981 257721 4984
rect 257755 5012 257767 5015
rect 258000 5012 258028 5052
rect 258626 5040 258632 5052
rect 258684 5040 258690 5092
rect 264425 5083 264483 5089
rect 264425 5080 264437 5083
rect 262784 5052 264437 5080
rect 257755 4984 258028 5012
rect 257755 4981 257767 4984
rect 257709 4975 257767 4981
rect 258810 4972 258816 5024
rect 258868 5012 258874 5024
rect 262784 5012 262812 5052
rect 264425 5049 264437 5052
rect 264471 5049 264483 5083
rect 264425 5043 264483 5049
rect 265342 5040 265348 5092
rect 265400 5080 265406 5092
rect 270144 5080 270172 5111
rect 265400 5052 270172 5080
rect 265400 5040 265406 5052
rect 258868 4984 262812 5012
rect 258868 4972 258874 4984
rect 264974 4972 264980 5024
rect 265032 5012 265038 5024
rect 265710 5012 265716 5024
rect 265032 4984 265716 5012
rect 265032 4972 265038 4984
rect 265710 4972 265716 4984
rect 265768 4972 265774 5024
rect 265897 5015 265955 5021
rect 265897 4981 265909 5015
rect 265943 5012 265955 5015
rect 267090 5012 267096 5024
rect 265943 4984 267096 5012
rect 265943 4981 265955 4984
rect 265897 4975 265955 4981
rect 267090 4972 267096 4984
rect 267148 5012 267154 5024
rect 267550 5012 267556 5024
rect 267148 4984 267556 5012
rect 267148 4972 267154 4984
rect 267550 4972 267556 4984
rect 267608 4972 267614 5024
rect 1104 4922 271492 4944
rect 1104 4870 34748 4922
rect 34800 4870 34812 4922
rect 34864 4870 34876 4922
rect 34928 4870 34940 4922
rect 34992 4870 35004 4922
rect 35056 4870 102345 4922
rect 102397 4870 102409 4922
rect 102461 4870 102473 4922
rect 102525 4870 102537 4922
rect 102589 4870 102601 4922
rect 102653 4870 169942 4922
rect 169994 4870 170006 4922
rect 170058 4870 170070 4922
rect 170122 4870 170134 4922
rect 170186 4870 170198 4922
rect 170250 4870 237539 4922
rect 237591 4870 237603 4922
rect 237655 4870 237667 4922
rect 237719 4870 237731 4922
rect 237783 4870 237795 4922
rect 237847 4870 271492 4922
rect 1104 4848 271492 4870
rect 3326 4768 3332 4820
rect 3384 4808 3390 4820
rect 28994 4808 29000 4820
rect 3384 4780 29000 4808
rect 3384 4768 3390 4780
rect 28994 4768 29000 4780
rect 29052 4768 29058 4820
rect 36998 4768 37004 4820
rect 37056 4768 37062 4820
rect 40954 4768 40960 4820
rect 41012 4768 41018 4820
rect 42794 4768 42800 4820
rect 42852 4768 42858 4820
rect 44082 4768 44088 4820
rect 44140 4808 44146 4820
rect 46750 4808 46756 4820
rect 44140 4780 46756 4808
rect 44140 4768 44146 4780
rect 46750 4768 46756 4780
rect 46808 4768 46814 4820
rect 48038 4768 48044 4820
rect 48096 4768 48102 4820
rect 48130 4768 48136 4820
rect 48188 4808 48194 4820
rect 55858 4808 55864 4820
rect 48188 4780 55864 4808
rect 48188 4768 48194 4780
rect 55858 4768 55864 4780
rect 55916 4768 55922 4820
rect 86954 4768 86960 4820
rect 87012 4808 87018 4820
rect 99466 4808 99472 4820
rect 87012 4780 99472 4808
rect 87012 4768 87018 4780
rect 99466 4768 99472 4780
rect 99524 4768 99530 4820
rect 100110 4768 100116 4820
rect 100168 4768 100174 4820
rect 100386 4768 100392 4820
rect 100444 4808 100450 4820
rect 100849 4811 100907 4817
rect 100849 4808 100861 4811
rect 100444 4780 100861 4808
rect 100444 4768 100450 4780
rect 100849 4777 100861 4780
rect 100895 4777 100907 4811
rect 100849 4771 100907 4777
rect 101214 4768 101220 4820
rect 101272 4808 101278 4820
rect 101309 4811 101367 4817
rect 101309 4808 101321 4811
rect 101272 4780 101321 4808
rect 101272 4768 101278 4780
rect 101309 4777 101321 4780
rect 101355 4777 101367 4811
rect 101309 4771 101367 4777
rect 102778 4768 102784 4820
rect 102836 4808 102842 4820
rect 103974 4808 103980 4820
rect 102836 4780 103980 4808
rect 102836 4768 102842 4780
rect 103974 4768 103980 4780
rect 104032 4768 104038 4820
rect 105998 4768 106004 4820
rect 106056 4768 106062 4820
rect 106090 4768 106096 4820
rect 106148 4808 106154 4820
rect 106148 4780 106596 4808
rect 106148 4768 106154 4780
rect 45462 4700 45468 4752
rect 45520 4740 45526 4752
rect 46382 4740 46388 4752
rect 45520 4712 46388 4740
rect 45520 4700 45526 4712
rect 46382 4700 46388 4712
rect 46440 4740 46446 4752
rect 46440 4712 46612 4740
rect 46440 4700 46446 4712
rect 42524 4684 42576 4690
rect 36814 4672 36820 4684
rect 36754 4644 36820 4672
rect 36814 4632 36820 4644
rect 36872 4672 36878 4684
rect 37090 4672 37096 4684
rect 36872 4644 37096 4672
rect 36872 4632 36878 4644
rect 37090 4632 37096 4644
rect 37148 4632 37154 4684
rect 42702 4632 42708 4684
rect 42760 4672 42766 4684
rect 46474 4672 46480 4684
rect 42760 4644 46480 4672
rect 42760 4632 42766 4644
rect 46474 4632 46480 4644
rect 46532 4632 46538 4684
rect 46584 4658 46612 4712
rect 50890 4700 50896 4752
rect 50948 4740 50954 4752
rect 51350 4740 51356 4752
rect 50948 4712 51356 4740
rect 50948 4700 50954 4712
rect 51350 4700 51356 4712
rect 51408 4740 51414 4752
rect 52362 4740 52368 4752
rect 51408 4712 52368 4740
rect 51408 4700 51414 4712
rect 52362 4700 52368 4712
rect 52420 4700 52426 4752
rect 92198 4700 92204 4752
rect 92256 4700 92262 4752
rect 103790 4740 103796 4752
rect 94424 4712 99788 4740
rect 50982 4632 50988 4684
rect 51040 4672 51046 4684
rect 51902 4672 51908 4684
rect 51040 4644 51908 4672
rect 51040 4632 51046 4644
rect 51902 4632 51908 4644
rect 51960 4632 51966 4684
rect 88334 4632 88340 4684
rect 88392 4672 88398 4684
rect 91557 4675 91615 4681
rect 91557 4672 91569 4675
rect 88392 4644 91569 4672
rect 88392 4632 88398 4644
rect 91557 4641 91569 4644
rect 91603 4641 91615 4675
rect 91557 4635 91615 4641
rect 92290 4632 92296 4684
rect 92348 4672 92354 4684
rect 92477 4675 92535 4681
rect 92477 4672 92489 4675
rect 92348 4644 92489 4672
rect 92348 4632 92354 4644
rect 92477 4641 92489 4644
rect 92523 4641 92535 4675
rect 92477 4635 92535 4641
rect 92615 4675 92673 4681
rect 92615 4641 92627 4675
rect 92661 4672 92673 4675
rect 94424 4672 94452 4712
rect 92661 4644 94452 4672
rect 92661 4641 92673 4644
rect 92615 4635 92673 4641
rect 94498 4632 94504 4684
rect 94556 4632 94562 4684
rect 94590 4632 94596 4684
rect 94648 4672 94654 4684
rect 97445 4675 97503 4681
rect 97445 4672 97457 4675
rect 94648 4644 97457 4672
rect 94648 4632 94654 4644
rect 97445 4641 97457 4644
rect 97491 4641 97503 4675
rect 97445 4635 97503 4641
rect 97629 4675 97687 4681
rect 97629 4641 97641 4675
rect 97675 4672 97687 4675
rect 98362 4672 98368 4684
rect 97675 4644 98368 4672
rect 97675 4641 97687 4644
rect 97629 4635 97687 4641
rect 98362 4632 98368 4644
rect 98420 4632 98426 4684
rect 98638 4632 98644 4684
rect 98696 4632 98702 4684
rect 99760 4672 99788 4712
rect 99944 4712 103796 4740
rect 99944 4672 99972 4712
rect 103790 4700 103796 4712
rect 103848 4700 103854 4752
rect 105170 4700 105176 4752
rect 105228 4740 105234 4752
rect 105228 4712 106228 4740
rect 105228 4700 105234 4712
rect 99760 4644 99972 4672
rect 100846 4632 100852 4684
rect 100904 4672 100910 4684
rect 102321 4675 102379 4681
rect 102321 4672 102333 4675
rect 100904 4644 102333 4672
rect 100904 4632 100910 4644
rect 102321 4641 102333 4644
rect 102367 4641 102379 4675
rect 102321 4635 102379 4641
rect 102505 4675 102563 4681
rect 102505 4641 102517 4675
rect 102551 4672 102563 4675
rect 103146 4672 103152 4684
rect 102551 4644 103152 4672
rect 102551 4641 102563 4644
rect 102505 4635 102563 4641
rect 103146 4632 103152 4644
rect 103204 4632 103210 4684
rect 106090 4672 106096 4684
rect 105464 4644 106096 4672
rect 42524 4626 42576 4632
rect 35618 4564 35624 4616
rect 35676 4604 35682 4616
rect 35989 4607 36047 4613
rect 35989 4604 36001 4607
rect 35676 4576 36001 4604
rect 35676 4564 35682 4576
rect 35989 4573 36001 4576
rect 36035 4573 36047 4607
rect 37274 4604 37280 4616
rect 35989 4567 36047 4573
rect 36096 4576 37280 4604
rect 35176 4508 35848 4536
rect 21266 4428 21272 4480
rect 21324 4468 21330 4480
rect 35176 4477 35204 4508
rect 35161 4471 35219 4477
rect 35161 4468 35173 4471
rect 21324 4440 35173 4468
rect 21324 4428 21330 4440
rect 35161 4437 35173 4440
rect 35207 4437 35219 4471
rect 35161 4431 35219 4437
rect 35434 4428 35440 4480
rect 35492 4468 35498 4480
rect 35713 4471 35771 4477
rect 35713 4468 35725 4471
rect 35492 4440 35725 4468
rect 35492 4428 35498 4440
rect 35713 4437 35725 4440
rect 35759 4437 35771 4471
rect 35820 4468 35848 4508
rect 35894 4496 35900 4548
rect 35952 4536 35958 4548
rect 36096 4545 36124 4576
rect 37274 4564 37280 4576
rect 37332 4604 37338 4616
rect 38010 4604 38016 4616
rect 37332 4576 38016 4604
rect 37332 4564 37338 4576
rect 38010 4564 38016 4576
rect 38068 4564 38074 4616
rect 41782 4564 41788 4616
rect 41840 4564 41846 4616
rect 42242 4564 42248 4616
rect 42300 4564 42306 4616
rect 44358 4564 44364 4616
rect 44416 4604 44422 4616
rect 46934 4604 46940 4616
rect 44416 4576 46940 4604
rect 44416 4564 44422 4576
rect 46934 4564 46940 4576
rect 46992 4564 46998 4616
rect 47026 4564 47032 4616
rect 47084 4564 47090 4616
rect 47486 4564 47492 4616
rect 47544 4564 47550 4616
rect 81434 4564 81440 4616
rect 81492 4604 81498 4616
rect 91741 4607 91799 4613
rect 91741 4604 91753 4607
rect 81492 4576 91753 4604
rect 81492 4564 81498 4576
rect 91741 4573 91753 4576
rect 91787 4573 91799 4607
rect 91741 4567 91799 4573
rect 92750 4564 92756 4616
rect 92808 4564 92814 4616
rect 94314 4564 94320 4616
rect 94372 4564 94378 4616
rect 96430 4564 96436 4616
rect 96488 4604 96494 4616
rect 96709 4607 96767 4613
rect 96709 4604 96721 4607
rect 96488 4576 96721 4604
rect 96488 4564 96494 4576
rect 96709 4573 96721 4576
rect 96755 4573 96767 4607
rect 96709 4567 96767 4573
rect 99374 4564 99380 4616
rect 99432 4604 99438 4616
rect 99745 4607 99803 4613
rect 99745 4604 99757 4607
rect 99432 4576 99757 4604
rect 99432 4564 99438 4576
rect 99745 4573 99757 4576
rect 99791 4573 99803 4607
rect 99745 4567 99803 4573
rect 100113 4607 100171 4613
rect 100113 4573 100125 4607
rect 100159 4573 100171 4607
rect 100113 4567 100171 4573
rect 36081 4539 36139 4545
rect 36081 4536 36093 4539
rect 35952 4508 36093 4536
rect 35952 4496 35958 4508
rect 36081 4505 36093 4508
rect 36127 4505 36139 4539
rect 36081 4499 36139 4505
rect 36446 4496 36452 4548
rect 36504 4496 36510 4548
rect 36538 4496 36544 4548
rect 36596 4536 36602 4548
rect 36596 4508 41828 4536
rect 36596 4496 36602 4508
rect 36817 4471 36875 4477
rect 36817 4468 36829 4471
rect 35820 4440 36829 4468
rect 35713 4431 35771 4437
rect 36817 4437 36829 4440
rect 36863 4437 36875 4471
rect 36817 4431 36875 4437
rect 41509 4471 41567 4477
rect 41509 4437 41521 4471
rect 41555 4468 41567 4471
rect 41598 4468 41604 4480
rect 41555 4440 41604 4468
rect 41555 4437 41567 4440
rect 41509 4431 41567 4437
rect 41598 4428 41604 4440
rect 41656 4428 41662 4480
rect 41800 4468 41828 4508
rect 41874 4496 41880 4548
rect 41932 4496 41938 4548
rect 45738 4496 45744 4548
rect 45796 4536 45802 4548
rect 46198 4536 46204 4548
rect 45796 4508 46204 4536
rect 45796 4496 45802 4508
rect 46198 4496 46204 4508
rect 46256 4536 46262 4548
rect 47121 4539 47179 4545
rect 47121 4536 47133 4539
rect 46256 4508 47133 4536
rect 46256 4496 46262 4508
rect 47121 4505 47133 4508
rect 47167 4536 47179 4539
rect 48314 4536 48320 4548
rect 47167 4508 48320 4536
rect 47167 4505 47179 4508
rect 47121 4499 47179 4505
rect 48314 4496 48320 4508
rect 48372 4536 48378 4548
rect 48498 4536 48504 4548
rect 48372 4508 48504 4536
rect 48372 4496 48378 4508
rect 48498 4496 48504 4508
rect 48556 4496 48562 4548
rect 49786 4496 49792 4548
rect 49844 4536 49850 4548
rect 55858 4536 55864 4548
rect 49844 4508 55864 4536
rect 49844 4496 49850 4508
rect 55858 4496 55864 4508
rect 55916 4496 55922 4548
rect 93486 4496 93492 4548
rect 93544 4536 93550 4548
rect 94682 4536 94688 4548
rect 93544 4508 94688 4536
rect 93544 4496 93550 4508
rect 94682 4496 94688 4508
rect 94740 4496 94746 4548
rect 96154 4496 96160 4548
rect 96212 4496 96218 4548
rect 97166 4496 97172 4548
rect 97224 4536 97230 4548
rect 97224 4508 98500 4536
rect 97224 4496 97230 4508
rect 42613 4471 42671 4477
rect 42613 4468 42625 4471
rect 41800 4440 42625 4468
rect 42613 4437 42625 4440
rect 42659 4437 42671 4471
rect 42613 4431 42671 4437
rect 44450 4428 44456 4480
rect 44508 4468 44514 4480
rect 45278 4468 45284 4480
rect 44508 4440 45284 4468
rect 44508 4428 44514 4440
rect 45278 4428 45284 4440
rect 45336 4428 45342 4480
rect 46753 4471 46811 4477
rect 46753 4437 46765 4471
rect 46799 4468 46811 4471
rect 47026 4468 47032 4480
rect 46799 4440 47032 4468
rect 46799 4437 46811 4440
rect 46753 4431 46811 4437
rect 47026 4428 47032 4440
rect 47084 4428 47090 4480
rect 47854 4428 47860 4480
rect 47912 4428 47918 4480
rect 47946 4428 47952 4480
rect 48004 4468 48010 4480
rect 48682 4468 48688 4480
rect 48004 4440 48688 4468
rect 48004 4428 48010 4440
rect 48682 4428 48688 4440
rect 48740 4468 48746 4480
rect 49050 4468 49056 4480
rect 48740 4440 49056 4468
rect 48740 4428 48746 4440
rect 49050 4428 49056 4440
rect 49108 4428 49114 4480
rect 92382 4428 92388 4480
rect 92440 4468 92446 4480
rect 93026 4468 93032 4480
rect 92440 4440 93032 4468
rect 92440 4428 92446 4440
rect 93026 4428 93032 4440
rect 93084 4428 93090 4480
rect 93397 4471 93455 4477
rect 93397 4437 93409 4471
rect 93443 4468 93455 4471
rect 94590 4468 94596 4480
rect 93443 4440 94596 4468
rect 93443 4437 93455 4440
rect 93397 4431 93455 4437
rect 94590 4428 94596 4440
rect 94648 4428 94654 4480
rect 95326 4428 95332 4480
rect 95384 4468 95390 4480
rect 95602 4468 95608 4480
rect 95384 4440 95608 4468
rect 95384 4428 95390 4440
rect 95602 4428 95608 4440
rect 95660 4428 95666 4480
rect 96893 4471 96951 4477
rect 96893 4437 96905 4471
rect 96939 4468 96951 4471
rect 97534 4468 97540 4480
rect 96939 4440 97540 4468
rect 96939 4437 96951 4440
rect 96893 4431 96951 4437
rect 97534 4428 97540 4440
rect 97592 4428 97598 4480
rect 98472 4468 98500 4508
rect 99558 4496 99564 4548
rect 99616 4536 99622 4548
rect 100128 4536 100156 4567
rect 100294 4564 100300 4616
rect 100352 4604 100358 4616
rect 100757 4607 100815 4613
rect 100757 4604 100769 4607
rect 100352 4576 100769 4604
rect 100352 4564 100358 4576
rect 100757 4573 100769 4576
rect 100803 4573 100815 4607
rect 100757 4567 100815 4573
rect 101033 4607 101091 4613
rect 101033 4573 101045 4607
rect 101079 4573 101091 4607
rect 101033 4567 101091 4573
rect 104805 4607 104863 4613
rect 104805 4573 104817 4607
rect 104851 4604 104863 4607
rect 104894 4604 104900 4616
rect 104851 4576 104900 4604
rect 104851 4573 104863 4576
rect 104805 4567 104863 4573
rect 100570 4536 100576 4548
rect 99616 4508 100576 4536
rect 99616 4496 99622 4508
rect 100570 4496 100576 4508
rect 100628 4536 100634 4548
rect 101048 4536 101076 4567
rect 104894 4564 104900 4576
rect 104952 4564 104958 4616
rect 105464 4613 105492 4644
rect 106090 4632 106096 4644
rect 106148 4632 106154 4684
rect 106200 4681 106228 4712
rect 106458 4700 106464 4752
rect 106516 4700 106522 4752
rect 106568 4740 106596 4780
rect 106918 4768 106924 4820
rect 106976 4808 106982 4820
rect 107105 4811 107163 4817
rect 107105 4808 107117 4811
rect 106976 4780 107117 4808
rect 106976 4768 106982 4780
rect 107105 4777 107117 4780
rect 107151 4808 107163 4811
rect 108117 4811 108175 4817
rect 108117 4808 108129 4811
rect 107151 4780 108129 4808
rect 107151 4777 107163 4780
rect 107105 4771 107163 4777
rect 108117 4777 108129 4780
rect 108163 4777 108175 4811
rect 108117 4771 108175 4777
rect 108206 4768 108212 4820
rect 108264 4808 108270 4820
rect 112165 4811 112223 4817
rect 108264 4780 108712 4808
rect 108264 4768 108270 4780
rect 108577 4743 108635 4749
rect 108577 4740 108589 4743
rect 106568 4712 108589 4740
rect 108577 4709 108589 4712
rect 108623 4709 108635 4743
rect 108577 4703 108635 4709
rect 106185 4675 106243 4681
rect 106185 4641 106197 4675
rect 106231 4641 106243 4675
rect 106185 4635 106243 4641
rect 107289 4675 107347 4681
rect 107289 4641 107301 4675
rect 107335 4672 107347 4675
rect 107378 4672 107384 4684
rect 107335 4644 107384 4672
rect 107335 4641 107347 4644
rect 107289 4635 107347 4641
rect 107378 4632 107384 4644
rect 107436 4672 107442 4684
rect 108684 4672 108712 4780
rect 112165 4777 112177 4811
rect 112211 4808 112223 4811
rect 113818 4808 113824 4820
rect 112211 4780 113824 4808
rect 112211 4777 112223 4780
rect 112165 4771 112223 4777
rect 113818 4768 113824 4780
rect 113876 4768 113882 4820
rect 114002 4768 114008 4820
rect 114060 4808 114066 4820
rect 114097 4811 114155 4817
rect 114097 4808 114109 4811
rect 114060 4780 114109 4808
rect 114060 4768 114066 4780
rect 114097 4777 114109 4780
rect 114143 4808 114155 4811
rect 114370 4808 114376 4820
rect 114143 4780 114376 4808
rect 114143 4777 114155 4780
rect 114097 4771 114155 4777
rect 114370 4768 114376 4780
rect 114428 4768 114434 4820
rect 114462 4768 114468 4820
rect 114520 4768 114526 4820
rect 117406 4768 117412 4820
rect 117464 4808 117470 4820
rect 117685 4811 117743 4817
rect 117685 4808 117697 4811
rect 117464 4780 117697 4808
rect 117464 4768 117470 4780
rect 117685 4777 117697 4780
rect 117731 4777 117743 4811
rect 118970 4808 118976 4820
rect 117685 4771 117743 4777
rect 117792 4780 118976 4808
rect 112809 4743 112867 4749
rect 112809 4709 112821 4743
rect 112855 4740 112867 4743
rect 113358 4740 113364 4752
rect 112855 4712 113364 4740
rect 112855 4709 112867 4712
rect 112809 4703 112867 4709
rect 113358 4700 113364 4712
rect 113416 4700 113422 4752
rect 113453 4743 113511 4749
rect 113453 4709 113465 4743
rect 113499 4740 113511 4743
rect 114830 4740 114836 4752
rect 113499 4712 114836 4740
rect 113499 4709 113511 4712
rect 113453 4703 113511 4709
rect 114830 4700 114836 4712
rect 114888 4700 114894 4752
rect 116302 4700 116308 4752
rect 116360 4740 116366 4752
rect 117792 4749 117820 4780
rect 118970 4768 118976 4780
rect 119028 4768 119034 4820
rect 120629 4811 120687 4817
rect 120629 4777 120641 4811
rect 120675 4808 120687 4811
rect 120902 4808 120908 4820
rect 120675 4780 120908 4808
rect 120675 4777 120687 4780
rect 120629 4771 120687 4777
rect 120902 4768 120908 4780
rect 120960 4808 120966 4820
rect 121641 4811 121699 4817
rect 121641 4808 121653 4811
rect 120960 4780 121653 4808
rect 120960 4768 120966 4780
rect 121641 4777 121653 4780
rect 121687 4777 121699 4811
rect 121641 4771 121699 4777
rect 117777 4743 117835 4749
rect 117777 4740 117789 4743
rect 116360 4712 117789 4740
rect 116360 4700 116366 4712
rect 117777 4709 117789 4712
rect 117823 4709 117835 4743
rect 117777 4703 117835 4709
rect 117961 4743 118019 4749
rect 117961 4709 117973 4743
rect 118007 4740 118019 4743
rect 118050 4740 118056 4752
rect 118007 4712 118056 4740
rect 118007 4709 118019 4712
rect 117961 4703 118019 4709
rect 118050 4700 118056 4712
rect 118108 4700 118114 4752
rect 118694 4700 118700 4752
rect 118752 4700 118758 4752
rect 119617 4743 119675 4749
rect 119617 4740 119629 4743
rect 118804 4712 119629 4740
rect 109313 4675 109371 4681
rect 109313 4672 109325 4675
rect 107436 4644 108436 4672
rect 108684 4644 109325 4672
rect 107436 4632 107442 4644
rect 105449 4607 105507 4613
rect 105449 4573 105461 4607
rect 105495 4573 105507 4607
rect 105449 4567 105507 4573
rect 105538 4564 105544 4616
rect 105596 4604 105602 4616
rect 105909 4607 105967 4613
rect 105909 4604 105921 4607
rect 105596 4576 105921 4604
rect 105596 4564 105602 4576
rect 105909 4573 105921 4576
rect 105955 4604 105967 4607
rect 107013 4607 107071 4613
rect 107013 4604 107025 4607
rect 105955 4600 106228 4604
rect 106384 4600 107025 4604
rect 105955 4576 107025 4600
rect 105955 4573 105967 4576
rect 105909 4567 105967 4573
rect 106200 4572 106412 4576
rect 107013 4573 107025 4576
rect 107059 4604 107071 4607
rect 107194 4604 107200 4616
rect 107059 4576 107200 4604
rect 107059 4573 107071 4576
rect 107013 4567 107071 4573
rect 107194 4564 107200 4576
rect 107252 4604 107258 4616
rect 108025 4607 108083 4613
rect 108025 4604 108037 4607
rect 107252 4576 108037 4604
rect 107252 4564 107258 4576
rect 108025 4573 108037 4576
rect 108071 4604 108083 4607
rect 108114 4604 108120 4616
rect 108071 4576 108120 4604
rect 108071 4573 108083 4576
rect 108025 4567 108083 4573
rect 108114 4564 108120 4576
rect 108172 4564 108178 4616
rect 108408 4613 108436 4644
rect 109313 4641 109325 4644
rect 109359 4641 109371 4675
rect 109313 4635 109371 4641
rect 110874 4632 110880 4684
rect 110932 4672 110938 4684
rect 111978 4672 111984 4684
rect 110932 4644 111984 4672
rect 110932 4632 110938 4644
rect 111978 4632 111984 4644
rect 112036 4632 112042 4684
rect 113542 4672 113548 4684
rect 112364 4644 113548 4672
rect 108393 4607 108451 4613
rect 108393 4573 108405 4607
rect 108439 4604 108451 4607
rect 108758 4604 108764 4616
rect 108439 4576 108764 4604
rect 108439 4573 108451 4576
rect 108393 4567 108451 4573
rect 108758 4564 108764 4576
rect 108816 4564 108822 4616
rect 109126 4564 109132 4616
rect 109184 4564 109190 4616
rect 111610 4564 111616 4616
rect 111668 4564 111674 4616
rect 112364 4613 112392 4644
rect 113542 4632 113548 4644
rect 113600 4632 113606 4684
rect 115106 4672 115112 4684
rect 113652 4644 115112 4672
rect 112349 4607 112407 4613
rect 112349 4573 112361 4607
rect 112395 4573 112407 4607
rect 112349 4567 112407 4573
rect 112993 4607 113051 4613
rect 112993 4573 113005 4607
rect 113039 4604 113051 4607
rect 113082 4604 113088 4616
rect 113039 4576 113088 4604
rect 113039 4573 113051 4576
rect 112993 4567 113051 4573
rect 113082 4564 113088 4576
rect 113140 4564 113146 4616
rect 113652 4613 113680 4644
rect 115106 4632 115112 4644
rect 115164 4632 115170 4684
rect 117866 4632 117872 4684
rect 117924 4672 117930 4684
rect 118418 4672 118424 4684
rect 117924 4644 118424 4672
rect 117924 4632 117930 4644
rect 118418 4632 118424 4644
rect 118476 4672 118482 4684
rect 118804 4672 118832 4712
rect 119617 4709 119629 4712
rect 119663 4709 119675 4743
rect 119617 4703 119675 4709
rect 120813 4743 120871 4749
rect 120813 4709 120825 4743
rect 120859 4709 120871 4743
rect 121656 4740 121684 4771
rect 121822 4768 121828 4820
rect 121880 4768 121886 4820
rect 122745 4811 122803 4817
rect 122745 4777 122757 4811
rect 122791 4808 122803 4811
rect 137462 4808 137468 4820
rect 122791 4780 137468 4808
rect 122791 4777 122803 4780
rect 122745 4771 122803 4777
rect 122760 4740 122788 4771
rect 137462 4768 137468 4780
rect 137520 4768 137526 4820
rect 138842 4768 138848 4820
rect 138900 4808 138906 4820
rect 138900 4780 138980 4808
rect 138900 4768 138906 4780
rect 121656 4712 122788 4740
rect 120813 4703 120871 4709
rect 120828 4672 120856 4703
rect 118476 4644 118832 4672
rect 118896 4644 120856 4672
rect 118476 4632 118482 4644
rect 113637 4607 113695 4613
rect 113637 4573 113649 4607
rect 113683 4573 113695 4607
rect 113637 4567 113695 4573
rect 114094 4564 114100 4616
rect 114152 4564 114158 4616
rect 114278 4564 114284 4616
rect 114336 4564 114342 4616
rect 114922 4564 114928 4616
rect 114980 4564 114986 4616
rect 117314 4564 117320 4616
rect 117372 4604 117378 4616
rect 118510 4604 118516 4616
rect 117372 4576 118516 4604
rect 117372 4564 117378 4576
rect 118510 4564 118516 4576
rect 118568 4564 118574 4616
rect 118896 4613 118924 4644
rect 120994 4632 121000 4684
rect 121052 4672 121058 4684
rect 121549 4675 121607 4681
rect 121549 4672 121561 4675
rect 121052 4644 121561 4672
rect 121052 4632 121058 4644
rect 121549 4641 121561 4644
rect 121595 4672 121607 4675
rect 122742 4672 122748 4684
rect 121595 4644 122748 4672
rect 121595 4641 121607 4644
rect 121549 4635 121607 4641
rect 122742 4632 122748 4644
rect 122800 4632 122806 4684
rect 138201 4675 138259 4681
rect 138201 4641 138213 4675
rect 138247 4672 138259 4675
rect 138566 4672 138572 4684
rect 138247 4644 138572 4672
rect 138247 4641 138259 4644
rect 138201 4635 138259 4641
rect 138566 4632 138572 4644
rect 138624 4632 138630 4684
rect 138842 4632 138848 4684
rect 138900 4632 138906 4684
rect 138952 4672 138980 4780
rect 139118 4768 139124 4820
rect 139176 4808 139182 4820
rect 140038 4808 140044 4820
rect 139176 4780 140044 4808
rect 139176 4768 139182 4780
rect 140038 4768 140044 4780
rect 140096 4768 140102 4820
rect 141160 4780 142108 4808
rect 141160 4752 141188 4780
rect 139854 4700 139860 4752
rect 139912 4740 139918 4752
rect 139912 4712 140728 4740
rect 139912 4700 139918 4712
rect 138952 4644 139164 4672
rect 118881 4607 118939 4613
rect 118881 4573 118893 4607
rect 118927 4573 118939 4607
rect 118881 4567 118939 4573
rect 119430 4564 119436 4616
rect 119488 4564 119494 4616
rect 120261 4607 120319 4613
rect 120261 4573 120273 4607
rect 120307 4573 120319 4607
rect 120261 4567 120319 4573
rect 120629 4607 120687 4613
rect 120629 4573 120641 4607
rect 120675 4604 120687 4607
rect 121012 4604 121040 4632
rect 120675 4576 121040 4604
rect 120675 4573 120687 4576
rect 120629 4567 120687 4573
rect 100628 4508 101076 4536
rect 104161 4539 104219 4545
rect 100628 4496 100634 4508
rect 104161 4505 104173 4539
rect 104207 4536 104219 4539
rect 106550 4536 106556 4548
rect 104207 4508 106556 4536
rect 104207 4505 104219 4508
rect 104161 4499 104219 4505
rect 106550 4496 106556 4508
rect 106608 4496 106614 4548
rect 110969 4539 111027 4545
rect 110969 4505 110981 4539
rect 111015 4536 111027 4539
rect 111015 4508 113312 4536
rect 111015 4505 111027 4508
rect 110969 4499 111027 4505
rect 100297 4471 100355 4477
rect 100297 4468 100309 4471
rect 98472 4440 100309 4468
rect 100297 4437 100309 4440
rect 100343 4437 100355 4471
rect 100297 4431 100355 4437
rect 101398 4428 101404 4480
rect 101456 4468 101462 4480
rect 104342 4468 104348 4480
rect 101456 4440 104348 4468
rect 101456 4428 101462 4440
rect 104342 4428 104348 4440
rect 104400 4428 104406 4480
rect 104621 4471 104679 4477
rect 104621 4437 104633 4471
rect 104667 4468 104679 4471
rect 104710 4468 104716 4480
rect 104667 4440 104716 4468
rect 104667 4437 104679 4440
rect 104621 4431 104679 4437
rect 104710 4428 104716 4440
rect 104768 4428 104774 4480
rect 105265 4471 105323 4477
rect 105265 4437 105277 4471
rect 105311 4468 105323 4471
rect 106228 4468 106234 4480
rect 105311 4440 106234 4468
rect 105311 4437 105323 4440
rect 105265 4431 105323 4437
rect 106228 4428 106234 4440
rect 106286 4428 106292 4480
rect 107470 4428 107476 4480
rect 107528 4468 107534 4480
rect 107565 4471 107623 4477
rect 107565 4468 107577 4471
rect 107528 4440 107577 4468
rect 107528 4428 107534 4440
rect 107565 4437 107577 4440
rect 107611 4437 107623 4471
rect 107565 4431 107623 4437
rect 111429 4471 111487 4477
rect 111429 4437 111441 4471
rect 111475 4468 111487 4471
rect 111794 4468 111800 4480
rect 111475 4440 111800 4468
rect 111475 4437 111487 4440
rect 111429 4431 111487 4437
rect 111794 4428 111800 4440
rect 111852 4428 111858 4480
rect 113284 4468 113312 4508
rect 113358 4496 113364 4548
rect 113416 4536 113422 4548
rect 115109 4539 115167 4545
rect 115109 4536 115121 4539
rect 113416 4508 115121 4536
rect 113416 4496 113422 4508
rect 115109 4505 115121 4508
rect 115155 4505 115167 4539
rect 115109 4499 115167 4505
rect 116765 4539 116823 4545
rect 116765 4505 116777 4539
rect 116811 4536 116823 4539
rect 120074 4536 120080 4548
rect 116811 4508 120080 4536
rect 116811 4505 116823 4508
rect 116765 4499 116823 4505
rect 120074 4496 120080 4508
rect 120132 4496 120138 4548
rect 120276 4536 120304 4567
rect 121270 4564 121276 4616
rect 121328 4604 121334 4616
rect 122466 4604 122472 4616
rect 121328 4576 122472 4604
rect 121328 4564 121334 4576
rect 122466 4564 122472 4576
rect 122524 4564 122530 4616
rect 138382 4564 138388 4616
rect 138440 4564 138446 4616
rect 139136 4613 139164 4644
rect 139210 4632 139216 4684
rect 139268 4681 139274 4684
rect 139268 4675 139296 4681
rect 139284 4641 139296 4675
rect 139268 4635 139296 4641
rect 139397 4675 139455 4681
rect 139397 4641 139409 4675
rect 139443 4672 139455 4675
rect 139946 4672 139952 4684
rect 139443 4644 139952 4672
rect 139443 4641 139455 4644
rect 139397 4635 139455 4641
rect 139268 4632 139274 4635
rect 139946 4632 139952 4644
rect 140004 4672 140010 4684
rect 140004 4644 140360 4672
rect 140004 4632 140010 4644
rect 139121 4607 139179 4613
rect 139121 4573 139133 4607
rect 139167 4573 139179 4607
rect 140332 4604 140360 4644
rect 140406 4632 140412 4684
rect 140464 4672 140470 4684
rect 140700 4681 140728 4712
rect 141142 4700 141148 4752
rect 141200 4700 141206 4752
rect 142080 4740 142108 4780
rect 142246 4768 142252 4820
rect 142304 4808 142310 4820
rect 143169 4811 143227 4817
rect 143169 4808 143181 4811
rect 142304 4780 143181 4808
rect 142304 4768 142310 4780
rect 143169 4777 143181 4780
rect 143215 4808 143227 4811
rect 143442 4808 143448 4820
rect 143215 4780 143448 4808
rect 143215 4777 143227 4780
rect 143169 4771 143227 4777
rect 143442 4768 143448 4780
rect 143500 4768 143506 4820
rect 143626 4768 143632 4820
rect 143684 4768 143690 4820
rect 143736 4780 147674 4808
rect 143736 4740 143764 4780
rect 142080 4712 143764 4740
rect 147646 4740 147674 4780
rect 149164 4780 150756 4808
rect 147646 4712 148548 4740
rect 140501 4675 140559 4681
rect 140501 4672 140513 4675
rect 140464 4644 140513 4672
rect 140464 4632 140470 4644
rect 140501 4641 140513 4644
rect 140547 4641 140559 4675
rect 140501 4635 140559 4641
rect 140685 4675 140743 4681
rect 140685 4641 140697 4675
rect 140731 4641 140743 4675
rect 140685 4635 140743 4641
rect 141418 4632 141424 4684
rect 141476 4632 141482 4684
rect 141694 4632 141700 4684
rect 141752 4672 141758 4684
rect 141752 4644 142476 4672
rect 141752 4632 141758 4644
rect 141602 4613 141608 4616
rect 141559 4607 141608 4613
rect 140332 4576 140728 4604
rect 139121 4567 139179 4573
rect 120442 4536 120448 4548
rect 120276 4508 120448 4536
rect 120442 4496 120448 4508
rect 120500 4536 120506 4548
rect 121288 4536 121316 4564
rect 120500 4508 121316 4536
rect 120500 4496 120506 4508
rect 121362 4496 121368 4548
rect 121420 4536 121426 4548
rect 121420 4508 132494 4536
rect 121420 4496 121426 4508
rect 113726 4468 113732 4480
rect 113284 4440 113732 4468
rect 113726 4428 113732 4440
rect 113784 4428 113790 4480
rect 118234 4428 118240 4480
rect 118292 4468 118298 4480
rect 119982 4468 119988 4480
rect 118292 4440 119988 4468
rect 118292 4428 118298 4440
rect 119982 4428 119988 4440
rect 120040 4468 120046 4480
rect 122374 4468 122380 4480
rect 120040 4440 122380 4468
rect 120040 4428 120046 4440
rect 122374 4428 122380 4440
rect 122432 4428 122438 4480
rect 123018 4428 123024 4480
rect 123076 4428 123082 4480
rect 132466 4468 132494 4508
rect 135898 4468 135904 4480
rect 132466 4440 135904 4468
rect 135898 4428 135904 4440
rect 135956 4428 135962 4480
rect 139670 4428 139676 4480
rect 139728 4468 139734 4480
rect 140041 4471 140099 4477
rect 140041 4468 140053 4471
rect 139728 4440 140053 4468
rect 139728 4428 139734 4440
rect 140041 4437 140053 4440
rect 140087 4437 140099 4471
rect 140700 4468 140728 4576
rect 141559 4573 141571 4607
rect 141605 4573 141608 4607
rect 141559 4567 141608 4573
rect 141602 4564 141608 4567
rect 141660 4564 141666 4616
rect 141694 4468 141700 4480
rect 140700 4440 141700 4468
rect 140041 4431 140099 4437
rect 141694 4428 141700 4440
rect 141752 4428 141758 4480
rect 142154 4428 142160 4480
rect 142212 4468 142218 4480
rect 142341 4471 142399 4477
rect 142341 4468 142353 4471
rect 142212 4440 142353 4468
rect 142212 4428 142218 4440
rect 142341 4437 142353 4440
rect 142387 4437 142399 4471
rect 142448 4468 142476 4644
rect 143166 4632 143172 4684
rect 143224 4672 143230 4684
rect 143353 4675 143411 4681
rect 143353 4672 143365 4675
rect 143224 4644 143365 4672
rect 143224 4632 143230 4644
rect 143353 4641 143365 4644
rect 143399 4641 143411 4675
rect 143353 4635 143411 4641
rect 144362 4632 144368 4684
rect 144420 4672 144426 4684
rect 144457 4675 144515 4681
rect 144457 4672 144469 4675
rect 144420 4644 144469 4672
rect 144420 4632 144426 4644
rect 144457 4641 144469 4644
rect 144503 4641 144515 4675
rect 144457 4635 144515 4641
rect 144641 4675 144699 4681
rect 144641 4641 144653 4675
rect 144687 4672 144699 4675
rect 145006 4672 145012 4684
rect 144687 4644 145012 4672
rect 144687 4641 144699 4644
rect 144641 4635 144699 4641
rect 145006 4632 145012 4644
rect 145064 4632 145070 4684
rect 145098 4632 145104 4684
rect 145156 4632 145162 4684
rect 145374 4632 145380 4684
rect 145432 4632 145438 4684
rect 145653 4675 145711 4681
rect 145653 4641 145665 4675
rect 145699 4672 145711 4675
rect 146846 4672 146852 4684
rect 145699 4644 146852 4672
rect 145699 4641 145711 4644
rect 145653 4635 145711 4641
rect 146846 4632 146852 4644
rect 146904 4632 146910 4684
rect 142982 4564 142988 4616
rect 143040 4604 143046 4616
rect 145558 4613 145564 4616
rect 143077 4607 143135 4613
rect 143077 4604 143089 4607
rect 143040 4576 143089 4604
rect 143040 4564 143046 4576
rect 143077 4573 143089 4576
rect 143123 4573 143135 4607
rect 143077 4567 143135 4573
rect 145515 4607 145564 4613
rect 145515 4573 145527 4607
rect 145561 4573 145564 4607
rect 145515 4567 145564 4573
rect 145558 4564 145564 4567
rect 145616 4564 145622 4616
rect 147122 4564 147128 4616
rect 147180 4564 147186 4616
rect 148134 4604 148140 4616
rect 147232 4576 148140 4604
rect 147232 4536 147260 4576
rect 148134 4564 148140 4576
rect 148192 4564 148198 4616
rect 148410 4564 148416 4616
rect 148468 4564 148474 4616
rect 148520 4604 148548 4712
rect 148870 4632 148876 4684
rect 148928 4672 148934 4684
rect 149164 4681 149192 4780
rect 148965 4675 149023 4681
rect 148965 4672 148977 4675
rect 148928 4644 148977 4672
rect 148928 4632 148934 4644
rect 148965 4641 148977 4644
rect 149011 4641 149023 4675
rect 148965 4635 149023 4641
rect 149149 4675 149207 4681
rect 149149 4641 149161 4675
rect 149195 4641 149207 4675
rect 149609 4675 149667 4681
rect 149609 4672 149621 4675
rect 149149 4635 149207 4641
rect 149256 4644 149621 4672
rect 149256 4604 149284 4644
rect 149609 4641 149621 4644
rect 149655 4641 149667 4675
rect 149609 4635 149667 4641
rect 149882 4632 149888 4684
rect 149940 4632 149946 4684
rect 150158 4632 150164 4684
rect 150216 4672 150222 4684
rect 150342 4672 150348 4684
rect 150216 4644 150348 4672
rect 150216 4632 150222 4644
rect 150342 4632 150348 4644
rect 150400 4632 150406 4684
rect 150728 4672 150756 4780
rect 150894 4768 150900 4820
rect 150952 4808 150958 4820
rect 151357 4811 151415 4817
rect 151357 4808 151369 4811
rect 150952 4780 151369 4808
rect 150952 4768 150958 4780
rect 151357 4777 151369 4780
rect 151403 4808 151415 4811
rect 152369 4811 152427 4817
rect 151403 4780 151860 4808
rect 151403 4777 151415 4780
rect 151357 4771 151415 4777
rect 151832 4740 151860 4780
rect 152369 4777 152381 4811
rect 152415 4777 152427 4811
rect 152369 4771 152427 4777
rect 152384 4740 152412 4771
rect 153102 4768 153108 4820
rect 153160 4808 153166 4820
rect 154758 4808 154764 4820
rect 153160 4780 154764 4808
rect 153160 4768 153166 4780
rect 154758 4768 154764 4780
rect 154816 4768 154822 4820
rect 155862 4768 155868 4820
rect 155920 4808 155926 4820
rect 161382 4808 161388 4820
rect 155920 4780 161388 4808
rect 155920 4768 155926 4780
rect 161382 4768 161388 4780
rect 161440 4768 161446 4820
rect 165617 4811 165675 4817
rect 165617 4777 165629 4811
rect 165663 4808 165675 4811
rect 167178 4808 167184 4820
rect 165663 4780 167184 4808
rect 165663 4777 165675 4780
rect 165617 4771 165675 4777
rect 167178 4768 167184 4780
rect 167236 4808 167242 4820
rect 167236 4780 167868 4808
rect 167236 4768 167242 4780
rect 151832 4712 152412 4740
rect 153746 4700 153752 4752
rect 153804 4740 153810 4752
rect 153804 4712 155908 4740
rect 153804 4700 153810 4712
rect 151354 4672 151360 4684
rect 150728 4644 151360 4672
rect 151354 4632 151360 4644
rect 151412 4632 151418 4684
rect 152550 4632 152556 4684
rect 152608 4632 152614 4684
rect 152826 4632 152832 4684
rect 152884 4672 152890 4684
rect 153381 4675 153439 4681
rect 153381 4672 153393 4675
rect 152884 4644 153393 4672
rect 152884 4632 152890 4644
rect 153381 4641 153393 4644
rect 153427 4641 153439 4675
rect 153381 4635 153439 4641
rect 153562 4632 153568 4684
rect 153620 4632 153626 4684
rect 154574 4632 154580 4684
rect 154632 4632 154638 4684
rect 155880 4681 155908 4712
rect 156322 4700 156328 4752
rect 156380 4740 156386 4752
rect 167840 4740 167868 4780
rect 168098 4768 168104 4820
rect 168156 4768 168162 4820
rect 186314 4808 186320 4820
rect 168208 4780 186320 4808
rect 168208 4740 168236 4780
rect 186314 4768 186320 4780
rect 186372 4768 186378 4820
rect 208578 4768 208584 4820
rect 208636 4808 208642 4820
rect 216766 4808 216772 4820
rect 208636 4780 216772 4808
rect 208636 4768 208642 4780
rect 216766 4768 216772 4780
rect 216824 4768 216830 4820
rect 217226 4768 217232 4820
rect 217284 4808 217290 4820
rect 222838 4808 222844 4820
rect 217284 4780 222844 4808
rect 217284 4768 217290 4780
rect 222838 4768 222844 4780
rect 222896 4768 222902 4820
rect 222930 4768 222936 4820
rect 222988 4768 222994 4820
rect 223114 4768 223120 4820
rect 223172 4808 223178 4820
rect 223853 4811 223911 4817
rect 223853 4808 223865 4811
rect 223172 4780 223865 4808
rect 223172 4768 223178 4780
rect 223853 4777 223865 4780
rect 223899 4808 223911 4811
rect 224310 4808 224316 4820
rect 223899 4780 224316 4808
rect 223899 4777 223911 4780
rect 223853 4771 223911 4777
rect 224310 4768 224316 4780
rect 224368 4768 224374 4820
rect 224497 4811 224555 4817
rect 224497 4777 224509 4811
rect 224543 4808 224555 4811
rect 224543 4780 224908 4808
rect 224543 4777 224555 4780
rect 224497 4771 224555 4777
rect 156380 4712 158852 4740
rect 167840 4712 168236 4740
rect 169113 4743 169171 4749
rect 156380 4700 156386 4712
rect 158824 4684 158852 4712
rect 169113 4709 169125 4743
rect 169159 4740 169171 4743
rect 169846 4740 169852 4752
rect 169159 4712 169852 4740
rect 169159 4709 169171 4712
rect 169113 4703 169171 4709
rect 169846 4700 169852 4712
rect 169904 4700 169910 4752
rect 170858 4700 170864 4752
rect 170916 4740 170922 4752
rect 205634 4740 205640 4752
rect 170916 4712 205640 4740
rect 170916 4700 170922 4712
rect 205634 4700 205640 4712
rect 205692 4700 205698 4752
rect 206646 4740 206652 4752
rect 205928 4712 206652 4740
rect 155865 4675 155923 4681
rect 155865 4641 155877 4675
rect 155911 4641 155923 4675
rect 155865 4635 155923 4641
rect 156046 4632 156052 4684
rect 156104 4672 156110 4684
rect 156141 4675 156199 4681
rect 156141 4672 156153 4675
rect 156104 4644 156153 4672
rect 156104 4632 156110 4644
rect 156141 4641 156153 4644
rect 156187 4672 156199 4675
rect 156414 4672 156420 4684
rect 156187 4644 156420 4672
rect 156187 4641 156199 4644
rect 156141 4635 156199 4641
rect 156414 4632 156420 4644
rect 156472 4632 156478 4684
rect 156506 4632 156512 4684
rect 156564 4672 156570 4684
rect 158533 4675 158591 4681
rect 158533 4672 158545 4675
rect 156564 4644 158545 4672
rect 156564 4632 156570 4644
rect 158533 4641 158545 4644
rect 158579 4641 158591 4675
rect 158533 4635 158591 4641
rect 158806 4632 158812 4684
rect 158864 4672 158870 4684
rect 159177 4675 159235 4681
rect 159177 4672 159189 4675
rect 158864 4644 159189 4672
rect 158864 4632 158870 4644
rect 159177 4641 159189 4644
rect 159223 4672 159235 4675
rect 159223 4644 160324 4672
rect 159223 4641 159235 4644
rect 159177 4635 159235 4641
rect 150066 4613 150072 4616
rect 148520 4576 149284 4604
rect 150023 4607 150072 4613
rect 146128 4508 147260 4536
rect 146128 4468 146156 4508
rect 147306 4496 147312 4548
rect 147364 4496 147370 4548
rect 148318 4496 148324 4548
rect 148376 4536 148382 4548
rect 148520 4536 148548 4576
rect 150023 4573 150035 4607
rect 150069 4573 150072 4607
rect 150023 4567 150072 4573
rect 150066 4564 150072 4567
rect 150124 4564 150130 4616
rect 151262 4564 151268 4616
rect 151320 4564 151326 4616
rect 151538 4564 151544 4616
rect 151596 4564 151602 4616
rect 152277 4607 152335 4613
rect 152277 4573 152289 4607
rect 152323 4573 152335 4607
rect 152277 4567 152335 4573
rect 148376 4508 148548 4536
rect 151280 4536 151308 4564
rect 152297 4536 152325 4567
rect 155678 4564 155684 4616
rect 155736 4564 155742 4616
rect 158717 4607 158775 4613
rect 158717 4604 158729 4607
rect 157306 4576 158729 4604
rect 155862 4536 155868 4548
rect 151280 4508 152325 4536
rect 154960 4508 155868 4536
rect 148376 4496 148382 4508
rect 142448 4440 146156 4468
rect 142341 4431 142399 4437
rect 146294 4428 146300 4480
rect 146352 4428 146358 4480
rect 148229 4471 148287 4477
rect 148229 4437 148241 4471
rect 148275 4468 148287 4471
rect 148778 4468 148784 4480
rect 148275 4440 148784 4468
rect 148275 4437 148287 4440
rect 148229 4431 148287 4437
rect 148778 4428 148784 4440
rect 148836 4428 148842 4480
rect 150802 4428 150808 4480
rect 150860 4428 150866 4480
rect 151817 4471 151875 4477
rect 151817 4437 151829 4471
rect 151863 4468 151875 4471
rect 152550 4468 152556 4480
rect 151863 4440 152556 4468
rect 151863 4437 151875 4440
rect 151817 4431 151875 4437
rect 152550 4428 152556 4440
rect 152608 4428 152614 4480
rect 152826 4428 152832 4480
rect 152884 4428 152890 4480
rect 152918 4428 152924 4480
rect 152976 4468 152982 4480
rect 154960 4468 154988 4508
rect 155862 4496 155868 4508
rect 155920 4496 155926 4548
rect 152976 4440 154988 4468
rect 152976 4428 152982 4440
rect 155126 4428 155132 4480
rect 155184 4468 155190 4480
rect 157306 4468 157334 4576
rect 158717 4573 158729 4576
rect 158763 4573 158775 4607
rect 158717 4567 158775 4573
rect 159450 4564 159456 4616
rect 159508 4564 159514 4616
rect 159634 4613 159640 4616
rect 159591 4607 159640 4613
rect 159591 4573 159603 4607
rect 159637 4573 159640 4607
rect 159591 4567 159640 4573
rect 159634 4564 159640 4567
rect 159692 4564 159698 4616
rect 159726 4564 159732 4616
rect 159784 4564 159790 4616
rect 160296 4536 160324 4644
rect 164234 4632 164240 4684
rect 164292 4672 164298 4684
rect 166445 4675 166503 4681
rect 166445 4672 166457 4675
rect 164292 4644 166457 4672
rect 164292 4632 164298 4644
rect 166445 4641 166457 4644
rect 166491 4641 166503 4675
rect 166905 4675 166963 4681
rect 166905 4672 166917 4675
rect 166445 4635 166503 4641
rect 166552 4644 166917 4672
rect 164326 4564 164332 4616
rect 164384 4604 164390 4616
rect 166261 4607 166319 4613
rect 166261 4604 166273 4607
rect 164384 4576 166273 4604
rect 164384 4564 164390 4576
rect 166261 4573 166273 4576
rect 166307 4573 166319 4607
rect 166552 4604 166580 4644
rect 166905 4641 166917 4644
rect 166951 4641 166963 4675
rect 166905 4635 166963 4641
rect 167295 4632 167301 4684
rect 167353 4681 167359 4684
rect 167353 4675 167377 4681
rect 167365 4641 167377 4675
rect 167353 4635 167377 4641
rect 167353 4632 167359 4635
rect 168282 4632 168288 4684
rect 168340 4672 168346 4684
rect 168340 4644 176654 4672
rect 168340 4632 168346 4644
rect 166261 4567 166319 4573
rect 166460 4576 166580 4604
rect 166460 4536 166488 4576
rect 167178 4564 167184 4616
rect 167236 4564 167242 4616
rect 167454 4564 167460 4616
rect 167512 4564 167518 4616
rect 168929 4607 168987 4613
rect 168929 4573 168941 4607
rect 168975 4604 168987 4607
rect 169386 4604 169392 4616
rect 168975 4576 169392 4604
rect 168975 4573 168987 4576
rect 168929 4567 168987 4573
rect 169386 4564 169392 4576
rect 169444 4564 169450 4616
rect 176626 4604 176654 4644
rect 195946 4644 205864 4672
rect 195946 4604 195974 4644
rect 205836 4616 205864 4644
rect 176626 4576 195974 4604
rect 205634 4564 205640 4616
rect 205692 4564 205698 4616
rect 205729 4607 205787 4613
rect 205729 4573 205741 4607
rect 205775 4573 205787 4607
rect 205729 4567 205787 4573
rect 160296 4508 166488 4536
rect 155184 4440 157334 4468
rect 155184 4428 155190 4440
rect 160370 4428 160376 4480
rect 160428 4428 160434 4480
rect 165982 4428 165988 4480
rect 166040 4428 166046 4480
rect 166460 4468 166488 4508
rect 169846 4496 169852 4548
rect 169904 4536 169910 4548
rect 205744 4536 205772 4567
rect 205818 4564 205824 4616
rect 205876 4564 205882 4616
rect 205928 4536 205956 4712
rect 206646 4700 206652 4712
rect 206704 4740 206710 4752
rect 210142 4740 210148 4752
rect 206704 4712 210148 4740
rect 206704 4700 206710 4712
rect 210142 4700 210148 4712
rect 210200 4700 210206 4752
rect 212166 4700 212172 4752
rect 212224 4700 212230 4752
rect 212537 4743 212595 4749
rect 212537 4709 212549 4743
rect 212583 4740 212595 4743
rect 212583 4712 213592 4740
rect 212583 4709 212595 4712
rect 212537 4703 212595 4709
rect 206462 4632 206468 4684
rect 206520 4632 206526 4684
rect 211430 4672 211436 4684
rect 208320 4644 211436 4672
rect 207934 4564 207940 4616
rect 207992 4604 207998 4616
rect 208320 4604 208348 4644
rect 211430 4632 211436 4644
rect 211488 4632 211494 4684
rect 212626 4632 212632 4684
rect 212684 4672 212690 4684
rect 212813 4675 212871 4681
rect 212813 4672 212825 4675
rect 212684 4644 212825 4672
rect 212684 4632 212690 4644
rect 212813 4641 212825 4644
rect 212859 4641 212871 4675
rect 212813 4635 212871 4641
rect 213454 4632 213460 4684
rect 213512 4632 213518 4684
rect 213564 4672 213592 4712
rect 214558 4700 214564 4752
rect 214616 4740 214622 4752
rect 219986 4740 219992 4752
rect 214616 4712 219992 4740
rect 214616 4700 214622 4712
rect 219986 4700 219992 4712
rect 220044 4700 220050 4752
rect 220814 4700 220820 4752
rect 220872 4740 220878 4752
rect 220872 4712 221872 4740
rect 220872 4700 220878 4712
rect 213850 4675 213908 4681
rect 213850 4672 213862 4675
rect 213564 4644 213862 4672
rect 213850 4641 213862 4644
rect 213896 4672 213908 4675
rect 213896 4644 214604 4672
rect 213896 4641 213908 4644
rect 213850 4635 213908 4641
rect 207992 4576 208348 4604
rect 207992 4564 207998 4576
rect 208670 4564 208676 4616
rect 208728 4604 208734 4616
rect 208857 4607 208915 4613
rect 208857 4604 208869 4607
rect 208728 4576 208869 4604
rect 208728 4564 208734 4576
rect 208857 4573 208869 4576
rect 208903 4573 208915 4607
rect 208857 4567 208915 4573
rect 208949 4607 209007 4613
rect 208949 4573 208961 4607
rect 208995 4573 209007 4607
rect 208949 4567 209007 4573
rect 169904 4508 205956 4536
rect 206005 4539 206063 4545
rect 169904 4496 169910 4508
rect 206005 4505 206017 4539
rect 206051 4536 206063 4539
rect 206649 4539 206707 4545
rect 206649 4536 206661 4539
rect 206051 4508 206661 4536
rect 206051 4505 206063 4508
rect 206005 4499 206063 4505
rect 206649 4505 206661 4508
rect 206695 4505 206707 4539
rect 206649 4499 206707 4505
rect 207566 4496 207572 4548
rect 207624 4536 207630 4548
rect 208305 4539 208363 4545
rect 208305 4536 208317 4539
rect 207624 4508 208317 4536
rect 207624 4496 207630 4508
rect 208305 4505 208317 4508
rect 208351 4536 208363 4539
rect 208578 4536 208584 4548
rect 208351 4508 208584 4536
rect 208351 4505 208363 4508
rect 208305 4499 208363 4505
rect 208578 4496 208584 4508
rect 208636 4496 208642 4548
rect 208964 4536 208992 4567
rect 209038 4564 209044 4616
rect 209096 4604 209102 4616
rect 209958 4604 209964 4616
rect 209096 4576 209964 4604
rect 209096 4564 209102 4576
rect 209958 4564 209964 4576
rect 210016 4604 210022 4616
rect 210510 4604 210516 4616
rect 210016 4576 210516 4604
rect 210016 4564 210022 4576
rect 210510 4564 210516 4576
rect 210568 4564 210574 4616
rect 211338 4564 211344 4616
rect 211396 4604 211402 4616
rect 211525 4607 211583 4613
rect 211525 4604 211537 4607
rect 211396 4576 211537 4604
rect 211396 4564 211402 4576
rect 211525 4573 211537 4576
rect 211571 4573 211583 4607
rect 211525 4567 211583 4573
rect 211614 4564 211620 4616
rect 211672 4564 211678 4616
rect 211706 4564 211712 4616
rect 211764 4604 211770 4616
rect 211801 4607 211859 4613
rect 211801 4604 211813 4607
rect 211764 4576 211813 4604
rect 211764 4564 211770 4576
rect 211801 4573 211813 4576
rect 211847 4573 211859 4607
rect 211801 4567 211859 4573
rect 212994 4564 213000 4616
rect 213052 4564 213058 4616
rect 213730 4564 213736 4616
rect 213788 4564 213794 4616
rect 214006 4564 214012 4616
rect 214064 4564 214070 4616
rect 208872 4508 210096 4536
rect 208872 4480 208900 4508
rect 167178 4468 167184 4480
rect 166460 4440 167184 4468
rect 167178 4428 167184 4440
rect 167236 4428 167242 4480
rect 167270 4428 167276 4480
rect 167328 4468 167334 4480
rect 187602 4468 187608 4480
rect 167328 4440 187608 4468
rect 167328 4428 167334 4440
rect 187602 4428 187608 4440
rect 187660 4428 187666 4480
rect 208854 4428 208860 4480
rect 208912 4428 208918 4480
rect 209225 4471 209283 4477
rect 209225 4437 209237 4471
rect 209271 4468 209283 4471
rect 209958 4468 209964 4480
rect 209271 4440 209964 4468
rect 209271 4437 209283 4440
rect 209225 4431 209283 4437
rect 209958 4428 209964 4440
rect 210016 4428 210022 4480
rect 210068 4468 210096 4508
rect 210142 4496 210148 4548
rect 210200 4496 210206 4548
rect 214576 4536 214604 4644
rect 214742 4632 214748 4684
rect 214800 4672 214806 4684
rect 215389 4675 215447 4681
rect 215389 4672 215401 4675
rect 214800 4644 215401 4672
rect 214800 4632 214806 4644
rect 215389 4641 215401 4644
rect 215435 4641 215447 4675
rect 215389 4635 215447 4641
rect 217962 4632 217968 4684
rect 218020 4632 218026 4684
rect 218146 4632 218152 4684
rect 218204 4632 218210 4684
rect 218422 4632 218428 4684
rect 218480 4672 218486 4684
rect 219066 4672 219072 4684
rect 218480 4644 219072 4672
rect 218480 4632 218486 4644
rect 219066 4632 219072 4644
rect 219124 4632 219130 4684
rect 219434 4632 219440 4684
rect 219492 4632 219498 4684
rect 220354 4632 220360 4684
rect 220412 4672 220418 4684
rect 221093 4675 221151 4681
rect 221093 4672 221105 4675
rect 220412 4644 221105 4672
rect 220412 4632 220418 4644
rect 221093 4641 221105 4644
rect 221139 4641 221151 4675
rect 221734 4672 221740 4684
rect 221093 4635 221151 4641
rect 221200 4644 221740 4672
rect 214653 4607 214711 4613
rect 214653 4573 214665 4607
rect 214699 4604 214711 4607
rect 215205 4607 215263 4613
rect 215205 4604 215217 4607
rect 214699 4576 215217 4604
rect 214699 4573 214711 4576
rect 214653 4567 214711 4573
rect 215205 4573 215217 4576
rect 215251 4573 215263 4607
rect 220541 4607 220599 4613
rect 220541 4604 220553 4607
rect 215205 4567 215263 4573
rect 219360 4576 220553 4604
rect 216398 4536 216404 4548
rect 214576 4508 216404 4536
rect 216398 4496 216404 4508
rect 216456 4496 216462 4548
rect 217042 4496 217048 4548
rect 217100 4496 217106 4548
rect 217962 4496 217968 4548
rect 218020 4536 218026 4548
rect 218330 4536 218336 4548
rect 218020 4508 218336 4536
rect 218020 4496 218026 4508
rect 218330 4496 218336 4508
rect 218388 4496 218394 4548
rect 218422 4496 218428 4548
rect 218480 4536 218486 4548
rect 218698 4536 218704 4548
rect 218480 4508 218704 4536
rect 218480 4496 218486 4508
rect 218698 4496 218704 4508
rect 218756 4496 218762 4548
rect 218882 4496 218888 4548
rect 218940 4536 218946 4548
rect 219360 4536 219388 4576
rect 220541 4573 220553 4576
rect 220587 4573 220599 4607
rect 220541 4567 220599 4573
rect 220722 4564 220728 4616
rect 220780 4604 220786 4616
rect 221200 4604 221228 4644
rect 221734 4632 221740 4644
rect 221792 4632 221798 4684
rect 221844 4672 221872 4712
rect 223758 4700 223764 4752
rect 223816 4740 223822 4752
rect 224126 4740 224132 4752
rect 223816 4712 224132 4740
rect 223816 4700 223822 4712
rect 224126 4700 224132 4712
rect 224184 4700 224190 4752
rect 224328 4740 224356 4768
rect 224678 4740 224684 4752
rect 224328 4712 224684 4740
rect 224678 4700 224684 4712
rect 224736 4700 224742 4752
rect 224880 4740 224908 4780
rect 224954 4768 224960 4820
rect 225012 4808 225018 4820
rect 228082 4808 228088 4820
rect 225012 4780 228088 4808
rect 225012 4768 225018 4780
rect 228082 4768 228088 4780
rect 228140 4768 228146 4820
rect 228266 4768 228272 4820
rect 228324 4808 228330 4820
rect 245562 4808 245568 4820
rect 228324 4780 245568 4808
rect 228324 4768 228330 4780
rect 245562 4768 245568 4780
rect 245620 4768 245626 4820
rect 246482 4768 246488 4820
rect 246540 4808 246546 4820
rect 246942 4808 246948 4820
rect 246540 4780 246948 4808
rect 246540 4768 246546 4780
rect 246942 4768 246948 4780
rect 247000 4808 247006 4820
rect 248046 4808 248052 4820
rect 247000 4780 248052 4808
rect 247000 4768 247006 4780
rect 248046 4768 248052 4780
rect 248104 4808 248110 4820
rect 251174 4808 251180 4820
rect 248104 4780 251180 4808
rect 248104 4768 248110 4780
rect 251174 4768 251180 4780
rect 251232 4808 251238 4820
rect 251545 4811 251603 4817
rect 251545 4808 251557 4811
rect 251232 4780 251557 4808
rect 251232 4768 251238 4780
rect 251545 4777 251557 4780
rect 251591 4808 251603 4811
rect 252462 4808 252468 4820
rect 251591 4780 252468 4808
rect 251591 4777 251603 4780
rect 251545 4771 251603 4777
rect 252462 4768 252468 4780
rect 252520 4768 252526 4820
rect 252557 4811 252615 4817
rect 252557 4777 252569 4811
rect 252603 4808 252615 4811
rect 253014 4808 253020 4820
rect 252603 4780 253020 4808
rect 252603 4777 252615 4780
rect 252557 4771 252615 4777
rect 253014 4768 253020 4780
rect 253072 4768 253078 4820
rect 253198 4768 253204 4820
rect 253256 4808 253262 4820
rect 253256 4780 257844 4808
rect 253256 4768 253262 4780
rect 225414 4740 225420 4752
rect 224880 4712 225420 4740
rect 225414 4700 225420 4712
rect 225472 4700 225478 4752
rect 227806 4700 227812 4752
rect 227864 4740 227870 4752
rect 244737 4743 244795 4749
rect 227864 4712 244688 4740
rect 227864 4700 227870 4712
rect 244660 4672 244688 4712
rect 244737 4709 244749 4743
rect 244783 4740 244795 4743
rect 247494 4740 247500 4752
rect 244783 4712 247500 4740
rect 244783 4709 244795 4712
rect 244737 4703 244795 4709
rect 247494 4700 247500 4712
rect 247552 4700 247558 4752
rect 248230 4700 248236 4752
rect 248288 4740 248294 4752
rect 253106 4740 253112 4752
rect 248288 4712 250300 4740
rect 248288 4700 248294 4712
rect 247589 4675 247647 4681
rect 221844 4644 234614 4672
rect 244660 4644 245700 4672
rect 220780 4576 221228 4604
rect 221277 4607 221335 4613
rect 220780 4564 220786 4576
rect 221277 4573 221289 4607
rect 221323 4573 221335 4607
rect 221277 4567 221335 4573
rect 218940 4508 219388 4536
rect 218940 4496 218946 4508
rect 219526 4496 219532 4548
rect 219584 4536 219590 4548
rect 220630 4536 220636 4548
rect 219584 4508 220636 4536
rect 219584 4496 219590 4508
rect 220630 4496 220636 4508
rect 220688 4496 220694 4548
rect 210234 4468 210240 4480
rect 210068 4440 210240 4468
rect 210234 4428 210240 4440
rect 210292 4428 210298 4480
rect 210326 4428 210332 4480
rect 210384 4468 210390 4480
rect 215110 4468 215116 4480
rect 210384 4440 215116 4468
rect 210384 4428 210390 4440
rect 215110 4428 215116 4440
rect 215168 4428 215174 4480
rect 216214 4428 216220 4480
rect 216272 4468 216278 4480
rect 220170 4468 220176 4480
rect 216272 4440 220176 4468
rect 216272 4428 216278 4440
rect 220170 4428 220176 4440
rect 220228 4428 220234 4480
rect 220262 4428 220268 4480
rect 220320 4468 220326 4480
rect 220357 4471 220415 4477
rect 220357 4468 220369 4471
rect 220320 4440 220369 4468
rect 220320 4428 220326 4440
rect 220357 4437 220369 4440
rect 220403 4437 220415 4471
rect 221292 4468 221320 4567
rect 222010 4564 222016 4616
rect 222068 4564 222074 4616
rect 222102 4564 222108 4616
rect 222160 4613 222166 4616
rect 222160 4607 222188 4613
rect 222176 4573 222188 4607
rect 222160 4567 222188 4573
rect 222160 4564 222166 4567
rect 222286 4564 222292 4616
rect 222344 4564 222350 4616
rect 223206 4564 223212 4616
rect 223264 4604 223270 4616
rect 223669 4607 223727 4613
rect 223669 4604 223681 4607
rect 223264 4576 223681 4604
rect 223264 4564 223270 4576
rect 223669 4573 223681 4576
rect 223715 4573 223727 4607
rect 223669 4567 223727 4573
rect 223758 4564 223764 4616
rect 223816 4604 223822 4616
rect 223853 4607 223911 4613
rect 223853 4604 223865 4607
rect 223816 4576 223865 4604
rect 223816 4564 223822 4576
rect 223853 4573 223865 4576
rect 223899 4573 223911 4607
rect 224681 4607 224739 4613
rect 224681 4604 224693 4607
rect 223853 4567 223911 4573
rect 223960 4576 224693 4604
rect 222838 4496 222844 4548
rect 222896 4536 222902 4548
rect 223393 4539 223451 4545
rect 223393 4536 223405 4539
rect 222896 4508 223405 4536
rect 222896 4496 222902 4508
rect 223393 4505 223405 4508
rect 223439 4505 223451 4539
rect 223393 4499 223451 4505
rect 223482 4496 223488 4548
rect 223540 4536 223546 4548
rect 223960 4536 223988 4576
rect 224681 4573 224693 4576
rect 224727 4573 224739 4607
rect 224681 4567 224739 4573
rect 224770 4564 224776 4616
rect 224828 4604 224834 4616
rect 225509 4607 225567 4613
rect 225509 4604 225521 4607
rect 224828 4576 225521 4604
rect 224828 4564 224834 4576
rect 225509 4573 225521 4576
rect 225555 4573 225567 4607
rect 225509 4567 225567 4573
rect 227346 4564 227352 4616
rect 227404 4604 227410 4616
rect 227806 4604 227812 4616
rect 227404 4576 227812 4604
rect 227404 4564 227410 4576
rect 227806 4564 227812 4576
rect 227864 4564 227870 4616
rect 223540 4508 223988 4536
rect 223540 4496 223546 4508
rect 224126 4496 224132 4548
rect 224184 4536 224190 4548
rect 225693 4539 225751 4545
rect 225693 4536 225705 4539
rect 224184 4508 225705 4536
rect 224184 4496 224190 4508
rect 225693 4505 225705 4508
rect 225739 4505 225751 4539
rect 234586 4536 234614 4644
rect 244918 4564 244924 4616
rect 244976 4564 244982 4616
rect 245562 4564 245568 4616
rect 245620 4564 245626 4616
rect 245672 4604 245700 4644
rect 247589 4641 247601 4675
rect 247635 4672 247647 4675
rect 247678 4672 247684 4684
rect 247635 4644 247684 4672
rect 247635 4641 247647 4644
rect 247589 4635 247647 4641
rect 247678 4632 247684 4644
rect 247736 4632 247742 4684
rect 249058 4632 249064 4684
rect 249116 4632 249122 4684
rect 245672 4576 246804 4604
rect 246298 4536 246304 4548
rect 234586 4508 246304 4536
rect 225693 4499 225751 4505
rect 246298 4496 246304 4508
rect 246356 4496 246362 4548
rect 246574 4496 246580 4548
rect 246632 4536 246638 4548
rect 246669 4539 246727 4545
rect 246669 4536 246681 4539
rect 246632 4508 246681 4536
rect 246632 4496 246638 4508
rect 246669 4505 246681 4508
rect 246715 4505 246727 4539
rect 246776 4536 246804 4576
rect 246850 4564 246856 4616
rect 246908 4564 246914 4616
rect 246942 4564 246948 4616
rect 247000 4604 247006 4616
rect 247126 4604 247132 4616
rect 247000 4576 247132 4604
rect 247000 4564 247006 4576
rect 247126 4564 247132 4576
rect 247184 4604 247190 4616
rect 247184 4576 247448 4604
rect 247184 4564 247190 4576
rect 247310 4536 247316 4548
rect 246776 4508 247316 4536
rect 246669 4499 246727 4505
rect 247310 4496 247316 4508
rect 247368 4496 247374 4548
rect 247420 4536 247448 4576
rect 247770 4564 247776 4616
rect 247828 4604 247834 4616
rect 247865 4607 247923 4613
rect 247865 4604 247877 4607
rect 247828 4576 247877 4604
rect 247828 4564 247834 4576
rect 247865 4573 247877 4576
rect 247911 4604 247923 4607
rect 247911 4576 248368 4604
rect 247911 4573 247923 4576
rect 247865 4567 247923 4573
rect 248230 4536 248236 4548
rect 247420 4508 248236 4536
rect 248230 4496 248236 4508
rect 248288 4496 248294 4548
rect 248340 4536 248368 4576
rect 248874 4564 248880 4616
rect 248932 4564 248938 4616
rect 250272 4604 250300 4712
rect 250732 4712 253112 4740
rect 250732 4681 250760 4712
rect 253106 4700 253112 4712
rect 253164 4700 253170 4752
rect 254486 4740 254492 4752
rect 253308 4712 254492 4740
rect 250717 4675 250775 4681
rect 250717 4641 250729 4675
rect 250763 4641 250775 4675
rect 250717 4635 250775 4641
rect 251453 4675 251511 4681
rect 251453 4641 251465 4675
rect 251499 4672 251511 4675
rect 251634 4672 251640 4684
rect 251499 4644 251640 4672
rect 251499 4641 251511 4644
rect 251453 4635 251511 4641
rect 251634 4632 251640 4644
rect 251692 4632 251698 4684
rect 252741 4675 252799 4681
rect 252741 4641 252753 4675
rect 252787 4672 252799 4675
rect 253014 4672 253020 4684
rect 252787 4644 253020 4672
rect 252787 4641 252799 4644
rect 252741 4635 252799 4641
rect 253014 4632 253020 4644
rect 253072 4632 253078 4684
rect 251545 4607 251603 4613
rect 251545 4604 251557 4607
rect 250272 4576 251557 4604
rect 251545 4573 251557 4576
rect 251591 4573 251603 4607
rect 251545 4567 251603 4573
rect 251652 4576 252692 4604
rect 251266 4536 251272 4548
rect 248340 4508 251272 4536
rect 251266 4496 251272 4508
rect 251324 4496 251330 4548
rect 251358 4496 251364 4548
rect 251416 4536 251422 4548
rect 251560 4536 251588 4567
rect 251416 4508 251588 4536
rect 251416 4496 251422 4508
rect 222102 4468 222108 4480
rect 221292 4440 222108 4468
rect 220357 4431 220415 4437
rect 222102 4428 222108 4440
rect 222160 4428 222166 4480
rect 222286 4428 222292 4480
rect 222344 4468 222350 4480
rect 223114 4468 223120 4480
rect 222344 4440 223120 4468
rect 222344 4428 222350 4440
rect 223114 4428 223120 4440
rect 223172 4428 223178 4480
rect 224034 4428 224040 4480
rect 224092 4428 224098 4480
rect 224586 4428 224592 4480
rect 224644 4468 224650 4480
rect 227530 4468 227536 4480
rect 224644 4440 227536 4468
rect 224644 4428 224650 4440
rect 227530 4428 227536 4440
rect 227588 4428 227594 4480
rect 245378 4428 245384 4480
rect 245436 4428 245442 4480
rect 247126 4428 247132 4480
rect 247184 4428 247190 4480
rect 249702 4428 249708 4480
rect 249760 4468 249766 4480
rect 251652 4468 251680 4576
rect 252554 4496 252560 4548
rect 252612 4496 252618 4548
rect 252664 4536 252692 4576
rect 252830 4564 252836 4616
rect 252888 4604 252894 4616
rect 253308 4604 253336 4712
rect 254486 4700 254492 4712
rect 254544 4700 254550 4752
rect 257816 4740 257844 4780
rect 258626 4768 258632 4820
rect 258684 4808 258690 4820
rect 258721 4811 258779 4817
rect 258721 4808 258733 4811
rect 258684 4780 258733 4808
rect 258684 4768 258690 4780
rect 258721 4777 258733 4780
rect 258767 4777 258779 4811
rect 258721 4771 258779 4777
rect 259178 4768 259184 4820
rect 259236 4768 259242 4820
rect 260282 4768 260288 4820
rect 260340 4808 260346 4820
rect 264701 4811 264759 4817
rect 260340 4780 263594 4808
rect 260340 4768 260346 4780
rect 263566 4740 263594 4780
rect 264701 4777 264713 4811
rect 264747 4808 264759 4811
rect 265158 4808 265164 4820
rect 264747 4780 265164 4808
rect 264747 4777 264759 4780
rect 264701 4771 264759 4777
rect 265158 4768 265164 4780
rect 265216 4768 265222 4820
rect 265342 4768 265348 4820
rect 265400 4768 265406 4820
rect 265710 4768 265716 4820
rect 265768 4808 265774 4820
rect 265989 4811 266047 4817
rect 265989 4808 266001 4811
rect 265768 4780 266001 4808
rect 265768 4768 265774 4780
rect 265989 4777 266001 4780
rect 266035 4777 266047 4811
rect 265989 4771 266047 4777
rect 266906 4768 266912 4820
rect 266964 4808 266970 4820
rect 269022 4808 269028 4820
rect 266964 4780 269028 4808
rect 266964 4768 266970 4780
rect 269022 4768 269028 4780
rect 269080 4768 269086 4820
rect 270310 4768 270316 4820
rect 270368 4808 270374 4820
rect 270681 4811 270739 4817
rect 270681 4808 270693 4811
rect 270368 4780 270693 4808
rect 270368 4768 270374 4780
rect 270681 4777 270693 4780
rect 270727 4777 270739 4811
rect 270681 4771 270739 4777
rect 272150 4740 272156 4752
rect 257816 4712 261800 4740
rect 263566 4712 272156 4740
rect 256602 4632 256608 4684
rect 256660 4632 256666 4684
rect 257338 4632 257344 4684
rect 257396 4672 257402 4684
rect 257396 4644 257844 4672
rect 257396 4632 257402 4644
rect 252888 4576 253336 4604
rect 253385 4607 253443 4613
rect 252888 4564 252894 4576
rect 253385 4573 253397 4607
rect 253431 4573 253443 4607
rect 253385 4567 253443 4573
rect 252664 4508 252876 4536
rect 249760 4440 251680 4468
rect 251729 4471 251787 4477
rect 249760 4428 249766 4440
rect 251729 4437 251741 4471
rect 251775 4468 251787 4471
rect 252738 4468 252744 4480
rect 251775 4440 252744 4468
rect 251775 4437 251787 4440
rect 251729 4431 251787 4437
rect 252738 4428 252744 4440
rect 252796 4428 252802 4480
rect 252848 4468 252876 4508
rect 252922 4496 252928 4548
rect 252980 4496 252986 4548
rect 253400 4468 253428 4567
rect 255866 4564 255872 4616
rect 255924 4564 255930 4616
rect 256418 4564 256424 4616
rect 256476 4564 256482 4616
rect 257816 4604 257844 4644
rect 258718 4632 258724 4684
rect 258776 4672 258782 4684
rect 258813 4675 258871 4681
rect 258813 4672 258825 4675
rect 258776 4644 258825 4672
rect 258776 4632 258782 4644
rect 258813 4641 258825 4644
rect 258859 4641 258871 4675
rect 258813 4635 258871 4641
rect 258997 4607 259055 4613
rect 257816 4576 258764 4604
rect 253569 4539 253627 4545
rect 253569 4505 253581 4539
rect 253615 4536 253627 4539
rect 255225 4539 255283 4545
rect 253615 4508 253934 4536
rect 253615 4505 253627 4508
rect 253569 4499 253627 4505
rect 252848 4440 253428 4468
rect 253906 4468 253934 4508
rect 255225 4505 255237 4539
rect 255271 4536 255283 4539
rect 255271 4508 258212 4536
rect 255271 4505 255283 4508
rect 255225 4499 255283 4505
rect 255685 4471 255743 4477
rect 255685 4468 255697 4471
rect 253906 4440 255697 4468
rect 255685 4437 255697 4440
rect 255731 4437 255743 4471
rect 258184 4468 258212 4508
rect 258258 4496 258264 4548
rect 258316 4496 258322 4548
rect 258736 4545 258764 4576
rect 258997 4573 259009 4607
rect 259043 4604 259055 4607
rect 259362 4604 259368 4616
rect 259043 4576 259368 4604
rect 259043 4573 259055 4576
rect 258997 4567 259055 4573
rect 259362 4564 259368 4576
rect 259420 4564 259426 4616
rect 259822 4564 259828 4616
rect 259880 4564 259886 4616
rect 261772 4613 261800 4712
rect 272150 4700 272156 4712
rect 272208 4700 272214 4752
rect 268470 4672 268476 4684
rect 265544 4644 268476 4672
rect 261757 4607 261815 4613
rect 261757 4573 261769 4607
rect 261803 4573 261815 4607
rect 261757 4567 261815 4573
rect 264241 4607 264299 4613
rect 264241 4573 264253 4607
rect 264287 4604 264299 4607
rect 264330 4604 264336 4616
rect 264287 4576 264336 4604
rect 264287 4573 264299 4576
rect 264241 4567 264299 4573
rect 264330 4564 264336 4576
rect 264388 4564 264394 4616
rect 264885 4607 264943 4613
rect 264885 4573 264897 4607
rect 264931 4604 264943 4607
rect 265066 4604 265072 4616
rect 264931 4576 265072 4604
rect 264931 4573 264943 4576
rect 264885 4567 264943 4573
rect 265066 4564 265072 4576
rect 265124 4564 265130 4616
rect 265544 4613 265572 4644
rect 268470 4632 268476 4644
rect 268528 4632 268534 4684
rect 270037 4675 270095 4681
rect 270037 4672 270049 4675
rect 268580 4644 270049 4672
rect 265529 4607 265587 4613
rect 265529 4573 265541 4607
rect 265575 4573 265587 4607
rect 265529 4567 265587 4573
rect 266170 4564 266176 4616
rect 266228 4564 266234 4616
rect 266909 4607 266967 4613
rect 266909 4573 266921 4607
rect 266955 4604 266967 4607
rect 267642 4604 267648 4616
rect 266955 4576 267648 4604
rect 266955 4573 266967 4576
rect 266909 4567 266967 4573
rect 267642 4564 267648 4576
rect 267700 4564 267706 4616
rect 268580 4613 268608 4644
rect 270037 4641 270049 4644
rect 270083 4641 270095 4675
rect 270037 4635 270095 4641
rect 268565 4607 268623 4613
rect 268565 4573 268577 4607
rect 268611 4573 268623 4607
rect 268565 4567 268623 4573
rect 269206 4564 269212 4616
rect 269264 4604 269270 4616
rect 269669 4607 269727 4613
rect 269669 4604 269681 4607
rect 269264 4576 269681 4604
rect 269264 4564 269270 4576
rect 269669 4573 269681 4576
rect 269715 4573 269727 4607
rect 269669 4567 269727 4573
rect 269850 4564 269856 4616
rect 269908 4564 269914 4616
rect 270497 4607 270555 4613
rect 270497 4573 270509 4607
rect 270543 4604 270555 4607
rect 271046 4604 271052 4616
rect 270543 4576 271052 4604
rect 270543 4573 270555 4576
rect 270497 4567 270555 4573
rect 271046 4564 271052 4576
rect 271104 4564 271110 4616
rect 271138 4564 271144 4616
rect 271196 4604 271202 4616
rect 271966 4604 271972 4616
rect 271196 4576 271972 4604
rect 271196 4564 271202 4576
rect 271966 4564 271972 4576
rect 272024 4564 272030 4616
rect 258721 4539 258779 4545
rect 258721 4505 258733 4539
rect 258767 4536 258779 4539
rect 259178 4536 259184 4548
rect 258767 4508 259184 4536
rect 258767 4505 258779 4508
rect 258721 4499 258779 4505
rect 259178 4496 259184 4508
rect 259236 4496 259242 4548
rect 260834 4536 260840 4548
rect 259564 4508 260840 4536
rect 259564 4468 259592 4508
rect 260834 4496 260840 4508
rect 260892 4496 260898 4548
rect 263594 4496 263600 4548
rect 263652 4536 263658 4548
rect 267182 4536 267188 4548
rect 263652 4508 267188 4536
rect 263652 4496 263658 4508
rect 267182 4496 267188 4508
rect 267240 4496 267246 4548
rect 267274 4496 267280 4548
rect 267332 4496 267338 4548
rect 267550 4496 267556 4548
rect 267608 4536 267614 4548
rect 268933 4539 268991 4545
rect 268933 4536 268945 4539
rect 267608 4508 268945 4536
rect 267608 4496 267614 4508
rect 268933 4505 268945 4508
rect 268979 4505 268991 4539
rect 268933 4499 268991 4505
rect 269022 4496 269028 4548
rect 269080 4536 269086 4548
rect 271690 4536 271696 4548
rect 269080 4508 271696 4536
rect 269080 4496 269086 4508
rect 271690 4496 271696 4508
rect 271748 4496 271754 4548
rect 258184 4440 259592 4468
rect 259641 4471 259699 4477
rect 255685 4431 255743 4437
rect 259641 4437 259653 4471
rect 259687 4468 259699 4471
rect 259822 4468 259828 4480
rect 259687 4440 259828 4468
rect 259687 4437 259699 4440
rect 259641 4431 259699 4437
rect 259822 4428 259828 4440
rect 259880 4428 259886 4480
rect 261570 4428 261576 4480
rect 261628 4428 261634 4480
rect 264057 4471 264115 4477
rect 264057 4437 264069 4471
rect 264103 4468 264115 4471
rect 269758 4468 269764 4480
rect 264103 4440 269764 4468
rect 264103 4437 264115 4440
rect 264057 4431 264115 4437
rect 269758 4428 269764 4440
rect 269816 4428 269822 4480
rect 270402 4428 270408 4480
rect 270460 4468 270466 4480
rect 271046 4468 271052 4480
rect 270460 4440 271052 4468
rect 270460 4428 270466 4440
rect 271046 4428 271052 4440
rect 271104 4428 271110 4480
rect 1104 4378 271651 4400
rect 1104 4326 68546 4378
rect 68598 4326 68610 4378
rect 68662 4326 68674 4378
rect 68726 4326 68738 4378
rect 68790 4326 68802 4378
rect 68854 4326 136143 4378
rect 136195 4326 136207 4378
rect 136259 4326 136271 4378
rect 136323 4326 136335 4378
rect 136387 4326 136399 4378
rect 136451 4326 203740 4378
rect 203792 4326 203804 4378
rect 203856 4326 203868 4378
rect 203920 4326 203932 4378
rect 203984 4326 203996 4378
rect 204048 4326 271337 4378
rect 271389 4326 271401 4378
rect 271453 4326 271465 4378
rect 271517 4326 271529 4378
rect 271581 4326 271593 4378
rect 271645 4326 271651 4378
rect 1104 4304 271651 4326
rect 38378 4264 38384 4276
rect 36832 4236 38384 4264
rect 4430 4156 4436 4208
rect 4488 4196 4494 4208
rect 36832 4196 36860 4236
rect 38378 4224 38384 4236
rect 38436 4224 38442 4276
rect 41785 4267 41843 4273
rect 41785 4233 41797 4267
rect 41831 4264 41843 4267
rect 41874 4264 41880 4276
rect 41831 4236 41880 4264
rect 41831 4233 41843 4236
rect 41785 4227 41843 4233
rect 41874 4224 41880 4236
rect 41932 4224 41938 4276
rect 45738 4264 45744 4276
rect 44836 4236 45744 4264
rect 4488 4168 36860 4196
rect 4488 4156 4494 4168
rect 18046 4088 18052 4140
rect 18104 4128 18110 4140
rect 36722 4128 36728 4140
rect 18104 4100 36728 4128
rect 18104 4088 18110 4100
rect 36722 4088 36728 4100
rect 36780 4088 36786 4140
rect 36832 4137 36860 4168
rect 37645 4199 37703 4205
rect 37645 4165 37657 4199
rect 37691 4196 37703 4199
rect 37826 4196 37832 4208
rect 37691 4168 37832 4196
rect 37691 4165 37703 4168
rect 37645 4159 37703 4165
rect 37826 4156 37832 4168
rect 37884 4156 37890 4208
rect 38654 4196 38660 4208
rect 37936 4168 38660 4196
rect 37936 4137 37964 4168
rect 38654 4156 38660 4168
rect 38712 4156 38718 4208
rect 38746 4156 38752 4208
rect 38804 4196 38810 4208
rect 39301 4199 39359 4205
rect 39301 4196 39313 4199
rect 38804 4168 39313 4196
rect 38804 4156 38810 4168
rect 39301 4165 39313 4168
rect 39347 4165 39359 4199
rect 39301 4159 39359 4165
rect 41693 4199 41751 4205
rect 41693 4165 41705 4199
rect 41739 4196 41751 4199
rect 44358 4196 44364 4208
rect 41739 4168 44364 4196
rect 41739 4165 41751 4168
rect 41693 4159 41751 4165
rect 44358 4156 44364 4168
rect 44416 4156 44422 4208
rect 44450 4156 44456 4208
rect 44508 4156 44514 4208
rect 44836 4205 44864 4236
rect 45738 4224 45744 4236
rect 45796 4224 45802 4276
rect 48406 4224 48412 4276
rect 48464 4264 48470 4276
rect 49605 4267 49663 4273
rect 49605 4264 49617 4267
rect 48464 4236 49617 4264
rect 48464 4224 48470 4236
rect 49605 4233 49617 4236
rect 49651 4233 49663 4267
rect 49605 4227 49663 4233
rect 49786 4224 49792 4276
rect 49844 4224 49850 4276
rect 50525 4267 50583 4273
rect 50525 4233 50537 4267
rect 50571 4264 50583 4267
rect 51074 4264 51080 4276
rect 50571 4236 51080 4264
rect 50571 4233 50583 4236
rect 50525 4227 50583 4233
rect 51074 4224 51080 4236
rect 51132 4224 51138 4276
rect 55858 4224 55864 4276
rect 55916 4264 55922 4276
rect 100662 4264 100668 4276
rect 55916 4236 100668 4264
rect 55916 4224 55922 4236
rect 100662 4224 100668 4236
rect 100720 4224 100726 4276
rect 105814 4224 105820 4276
rect 105872 4264 105878 4276
rect 110785 4267 110843 4273
rect 105872 4236 110736 4264
rect 105872 4224 105878 4236
rect 44821 4199 44879 4205
rect 44821 4196 44833 4199
rect 44652 4168 44833 4196
rect 36817 4131 36875 4137
rect 36817 4097 36829 4131
rect 36863 4097 36875 4131
rect 36817 4091 36875 4097
rect 37921 4131 37979 4137
rect 37921 4097 37933 4131
rect 37967 4097 37979 4131
rect 37921 4091 37979 4097
rect 38010 4088 38016 4140
rect 38068 4088 38074 4140
rect 38378 4088 38384 4140
rect 38436 4128 38442 4140
rect 39669 4131 39727 4137
rect 39669 4128 39681 4131
rect 38436 4100 39681 4128
rect 38436 4088 38442 4100
rect 39669 4097 39681 4100
rect 39715 4097 39727 4131
rect 39669 4091 39727 4097
rect 42610 4088 42616 4140
rect 42668 4088 42674 4140
rect 43346 4088 43352 4140
rect 43404 4128 43410 4140
rect 44652 4128 44680 4168
rect 44821 4165 44833 4168
rect 44867 4165 44879 4199
rect 44821 4159 44879 4165
rect 45554 4156 45560 4208
rect 45612 4156 45618 4208
rect 48501 4199 48559 4205
rect 48501 4165 48513 4199
rect 48547 4196 48559 4199
rect 49142 4196 49148 4208
rect 48547 4168 49148 4196
rect 48547 4165 48559 4168
rect 48501 4159 48559 4165
rect 49142 4156 49148 4168
rect 49200 4156 49206 4208
rect 49237 4199 49295 4205
rect 49237 4165 49249 4199
rect 49283 4196 49295 4199
rect 49510 4196 49516 4208
rect 49283 4168 49516 4196
rect 49283 4165 49295 4168
rect 49237 4159 49295 4165
rect 49510 4156 49516 4168
rect 49568 4156 49574 4208
rect 50801 4199 50859 4205
rect 50264 4168 50752 4196
rect 43404 4100 44680 4128
rect 43404 4088 43410 4100
rect 44726 4088 44732 4140
rect 44784 4088 44790 4140
rect 45094 4088 45100 4140
rect 45152 4128 45158 4140
rect 45189 4131 45247 4137
rect 45189 4128 45201 4131
rect 45152 4100 45201 4128
rect 45152 4088 45158 4100
rect 45189 4097 45201 4100
rect 45235 4097 45247 4131
rect 45189 4091 45247 4097
rect 48590 4088 48596 4140
rect 48648 4128 48654 4140
rect 48777 4131 48835 4137
rect 48777 4128 48789 4131
rect 48648 4100 48789 4128
rect 48648 4088 48654 4100
rect 48777 4097 48789 4100
rect 48823 4097 48835 4131
rect 48777 4091 48835 4097
rect 48869 4131 48927 4137
rect 48869 4097 48881 4131
rect 48915 4128 48927 4131
rect 49050 4128 49056 4140
rect 48915 4100 49056 4128
rect 48915 4097 48927 4100
rect 48869 4091 48927 4097
rect 49050 4088 49056 4100
rect 49108 4128 49114 4140
rect 50264 4128 50292 4168
rect 49108 4100 50292 4128
rect 50724 4128 50752 4168
rect 50801 4165 50813 4199
rect 50847 4196 50859 4199
rect 50847 4168 51028 4196
rect 50847 4165 50859 4168
rect 50801 4159 50859 4165
rect 50890 4128 50896 4140
rect 50724 4100 50896 4128
rect 49108 4088 49114 4100
rect 50890 4088 50896 4100
rect 50948 4088 50954 4140
rect 51000 4128 51028 4168
rect 51166 4156 51172 4208
rect 51224 4196 51230 4208
rect 51261 4199 51319 4205
rect 51261 4196 51273 4199
rect 51224 4168 51273 4196
rect 51224 4156 51230 4168
rect 51261 4165 51273 4168
rect 51307 4165 51319 4199
rect 51261 4159 51319 4165
rect 51629 4199 51687 4205
rect 51629 4165 51641 4199
rect 51675 4196 51687 4199
rect 51718 4196 51724 4208
rect 51675 4168 51724 4196
rect 51675 4165 51687 4168
rect 51629 4159 51687 4165
rect 51718 4156 51724 4168
rect 51776 4156 51782 4208
rect 94498 4156 94504 4208
rect 94556 4196 94562 4208
rect 94556 4168 98592 4196
rect 94556 4156 94562 4168
rect 51810 4128 51816 4140
rect 51000 4100 51816 4128
rect 51810 4088 51816 4100
rect 51868 4088 51874 4140
rect 66901 4131 66959 4137
rect 66901 4097 66913 4131
rect 66947 4097 66959 4131
rect 92566 4128 92572 4140
rect 66901 4091 66959 4097
rect 80026 4100 92572 4128
rect 45468 4072 45520 4078
rect 12802 4020 12808 4072
rect 12860 4060 12866 4072
rect 36906 4060 36912 4072
rect 12860 4032 36912 4060
rect 12860 4020 12866 4032
rect 36906 4020 36912 4032
rect 36964 4020 36970 4072
rect 38470 4020 38476 4072
rect 38528 4020 38534 4072
rect 42518 4020 42524 4072
rect 42576 4060 42582 4072
rect 42797 4063 42855 4069
rect 42797 4060 42809 4063
rect 42576 4032 42809 4060
rect 42576 4020 42582 4032
rect 42797 4029 42809 4032
rect 42843 4029 42855 4063
rect 42797 4023 42855 4029
rect 47118 4020 47124 4072
rect 47176 4060 47182 4072
rect 47946 4060 47952 4072
rect 47176 4032 47952 4060
rect 47176 4020 47182 4032
rect 47946 4020 47952 4032
rect 48004 4060 48010 4072
rect 51626 4060 51632 4072
rect 48004 4032 48346 4060
rect 51566 4032 51632 4060
rect 48004 4020 48010 4032
rect 51626 4020 51632 4032
rect 51684 4060 51690 4072
rect 52086 4060 52092 4072
rect 51684 4032 52092 4060
rect 51684 4020 51690 4032
rect 52086 4020 52092 4032
rect 52144 4020 52150 4072
rect 66441 4063 66499 4069
rect 66441 4029 66453 4063
rect 66487 4060 66499 4063
rect 66916 4060 66944 4091
rect 80026 4060 80054 4100
rect 92566 4088 92572 4100
rect 92624 4088 92630 4140
rect 92934 4088 92940 4140
rect 92992 4088 92998 4140
rect 93578 4088 93584 4140
rect 93636 4088 93642 4140
rect 94590 4088 94596 4140
rect 94648 4088 94654 4140
rect 96338 4128 96344 4140
rect 95988 4100 96344 4128
rect 94406 4060 94412 4072
rect 66487 4032 80054 4060
rect 84488 4032 94412 4060
rect 66487 4029 66499 4032
rect 66441 4023 66499 4029
rect 45468 4014 45520 4020
rect 8018 3952 8024 4004
rect 8076 3992 8082 4004
rect 36538 3992 36544 4004
rect 8076 3964 36544 3992
rect 8076 3952 8082 3964
rect 36538 3952 36544 3964
rect 36596 3952 36602 4004
rect 36814 3952 36820 4004
rect 36872 3992 36878 4004
rect 37366 3992 37372 4004
rect 36872 3964 37372 3992
rect 36872 3952 36878 3964
rect 37366 3952 37372 3964
rect 37424 3952 37430 4004
rect 38930 3952 38936 4004
rect 38988 3952 38994 4004
rect 39022 3952 39028 4004
rect 39080 3992 39086 4004
rect 44082 3992 44088 4004
rect 39080 3964 44088 3992
rect 39080 3952 39086 3964
rect 44082 3952 44088 3964
rect 44140 3952 44146 4004
rect 51813 3995 51871 4001
rect 51813 3961 51825 3995
rect 51859 3992 51871 3995
rect 84488 3992 84516 4032
rect 94406 4020 94412 4032
rect 94464 4020 94470 4072
rect 94774 4020 94780 4072
rect 94832 4020 94838 4072
rect 95142 4020 95148 4072
rect 95200 4060 95206 4072
rect 95988 4060 96016 4100
rect 96338 4088 96344 4100
rect 96396 4088 96402 4140
rect 98564 4128 98592 4168
rect 98638 4156 98644 4208
rect 98696 4196 98702 4208
rect 98733 4199 98791 4205
rect 98733 4196 98745 4199
rect 98696 4168 98745 4196
rect 98696 4156 98702 4168
rect 98733 4165 98745 4168
rect 98779 4196 98791 4199
rect 99190 4196 99196 4208
rect 98779 4168 99196 4196
rect 98779 4165 98791 4168
rect 98733 4159 98791 4165
rect 99190 4156 99196 4168
rect 99248 4156 99254 4208
rect 101490 4196 101496 4208
rect 99300 4168 101496 4196
rect 99300 4128 99328 4168
rect 101490 4156 101496 4168
rect 101548 4156 101554 4208
rect 105538 4196 105544 4208
rect 104728 4168 105544 4196
rect 98564 4100 99328 4128
rect 102042 4088 102048 4140
rect 102100 4088 102106 4140
rect 104728 4137 104756 4168
rect 105538 4156 105544 4168
rect 105596 4156 105602 4208
rect 105998 4196 106004 4208
rect 105740 4168 106004 4196
rect 104713 4131 104771 4137
rect 104713 4097 104725 4131
rect 104759 4097 104771 4131
rect 105740 4128 105768 4168
rect 105998 4156 106004 4168
rect 106056 4156 106062 4208
rect 106274 4156 106280 4208
rect 106332 4196 106338 4208
rect 106918 4196 106924 4208
rect 106332 4168 106924 4196
rect 106332 4156 106338 4168
rect 106918 4156 106924 4168
rect 106976 4156 106982 4208
rect 108114 4156 108120 4208
rect 108172 4196 108178 4208
rect 110708 4196 110736 4236
rect 110785 4233 110797 4267
rect 110831 4264 110843 4267
rect 111610 4264 111616 4276
rect 110831 4236 111616 4264
rect 110831 4233 110843 4236
rect 110785 4227 110843 4233
rect 111610 4224 111616 4236
rect 111668 4224 111674 4276
rect 118234 4264 118240 4276
rect 111720 4236 118240 4264
rect 111720 4196 111748 4236
rect 118234 4224 118240 4236
rect 118292 4224 118298 4276
rect 137986 4236 147674 4264
rect 108172 4168 110276 4196
rect 110708 4168 111748 4196
rect 108172 4156 108178 4168
rect 108500 4137 108528 4168
rect 110248 4140 110276 4168
rect 116670 4156 116676 4208
rect 116728 4196 116734 4208
rect 116728 4168 117268 4196
rect 116728 4156 116734 4168
rect 104713 4091 104771 4097
rect 104912 4100 105768 4128
rect 108485 4131 108543 4137
rect 95200 4032 96016 4060
rect 95200 4020 95206 4032
rect 96154 4020 96160 4072
rect 96212 4020 96218 4072
rect 96890 4020 96896 4072
rect 96948 4020 96954 4072
rect 97077 4063 97135 4069
rect 97077 4029 97089 4063
rect 97123 4029 97135 4063
rect 97077 4023 97135 4029
rect 51859 3964 84516 3992
rect 51859 3961 51871 3964
rect 51813 3955 51871 3961
rect 89714 3952 89720 4004
rect 89772 3992 89778 4004
rect 93210 3992 93216 4004
rect 89772 3964 93216 3992
rect 89772 3952 89778 3964
rect 93210 3952 93216 3964
rect 93268 3952 93274 4004
rect 93397 3995 93455 4001
rect 93397 3961 93409 3995
rect 93443 3992 93455 3995
rect 96706 3992 96712 4004
rect 93443 3964 96712 3992
rect 93443 3961 93455 3964
rect 93397 3955 93455 3961
rect 96706 3952 96712 3964
rect 96764 3952 96770 4004
rect 97092 3992 97120 4023
rect 98270 4020 98276 4072
rect 98328 4060 98334 4072
rect 99285 4063 99343 4069
rect 99285 4060 99297 4063
rect 98328 4032 99297 4060
rect 98328 4020 98334 4032
rect 99285 4029 99297 4032
rect 99331 4029 99343 4063
rect 99285 4023 99343 4029
rect 99469 4063 99527 4069
rect 99469 4029 99481 4063
rect 99515 4029 99527 4063
rect 99469 4023 99527 4029
rect 101125 4063 101183 4069
rect 101125 4029 101137 4063
rect 101171 4060 101183 4063
rect 101214 4060 101220 4072
rect 101171 4032 101220 4060
rect 101171 4029 101183 4032
rect 101125 4023 101183 4029
rect 97810 3992 97816 4004
rect 97092 3964 97816 3992
rect 97810 3952 97816 3964
rect 97868 3952 97874 4004
rect 99484 3992 99512 4023
rect 101214 4020 101220 4032
rect 101272 4020 101278 4072
rect 102229 4063 102287 4069
rect 102229 4029 102241 4063
rect 102275 4060 102287 4063
rect 102962 4060 102968 4072
rect 102275 4032 102968 4060
rect 102275 4029 102287 4032
rect 102229 4023 102287 4029
rect 102962 4020 102968 4032
rect 103020 4020 103026 4072
rect 103885 4063 103943 4069
rect 103885 4029 103897 4063
rect 103931 4060 103943 4063
rect 104912 4060 104940 4100
rect 108485 4097 108497 4131
rect 108531 4097 108543 4131
rect 108485 4091 108543 4097
rect 108758 4088 108764 4140
rect 108816 4128 108822 4140
rect 109773 4131 109831 4137
rect 108816 4100 109540 4128
rect 108816 4088 108822 4100
rect 103931 4032 104940 4060
rect 104989 4063 105047 4069
rect 103931 4029 103943 4032
rect 103885 4023 103943 4029
rect 104989 4029 105001 4063
rect 105035 4060 105047 4063
rect 105170 4060 105176 4072
rect 105035 4032 105176 4060
rect 105035 4029 105047 4032
rect 104989 4023 105047 4029
rect 105170 4020 105176 4032
rect 105228 4020 105234 4072
rect 105354 4020 105360 4072
rect 105412 4060 105418 4072
rect 105725 4063 105783 4069
rect 105725 4060 105737 4063
rect 105412 4032 105737 4060
rect 105412 4020 105418 4032
rect 105725 4029 105737 4032
rect 105771 4029 105783 4063
rect 105725 4023 105783 4029
rect 105906 4020 105912 4072
rect 105964 4020 105970 4072
rect 105998 4020 106004 4072
rect 106056 4060 106062 4072
rect 107565 4063 107623 4069
rect 107565 4060 107577 4063
rect 106056 4032 107577 4060
rect 106056 4020 106062 4032
rect 107565 4029 107577 4032
rect 107611 4060 107623 4063
rect 108114 4060 108120 4072
rect 107611 4032 108120 4060
rect 107611 4029 107623 4032
rect 107565 4023 107623 4029
rect 108114 4020 108120 4032
rect 108172 4020 108178 4072
rect 108850 4020 108856 4072
rect 108908 4060 108914 4072
rect 109512 4060 109540 4100
rect 109773 4097 109785 4131
rect 109819 4128 109831 4131
rect 109954 4128 109960 4140
rect 109819 4100 109960 4128
rect 109819 4097 109831 4100
rect 109773 4091 109831 4097
rect 109954 4088 109960 4100
rect 110012 4088 110018 4140
rect 110230 4088 110236 4140
rect 110288 4088 110294 4140
rect 114186 4088 114192 4140
rect 114244 4088 114250 4140
rect 117038 4088 117044 4140
rect 117096 4088 117102 4140
rect 117240 4128 117268 4168
rect 120074 4156 120080 4208
rect 120132 4196 120138 4208
rect 122098 4196 122104 4208
rect 120132 4168 122104 4196
rect 120132 4156 120138 4168
rect 122098 4156 122104 4168
rect 122156 4156 122162 4208
rect 137986 4196 138014 4236
rect 137296 4168 138014 4196
rect 117240 4100 117360 4128
rect 110506 4060 110512 4072
rect 108908 4032 109448 4060
rect 109512 4032 110512 4060
rect 108908 4020 108914 4032
rect 97920 3964 99512 3992
rect 28994 3884 29000 3936
rect 29052 3924 29058 3936
rect 36722 3924 36728 3936
rect 29052 3896 36728 3924
rect 29052 3884 29058 3896
rect 36722 3884 36728 3896
rect 36780 3884 36786 3936
rect 41138 3884 41144 3936
rect 41196 3924 41202 3936
rect 41874 3924 41880 3936
rect 41196 3896 41880 3924
rect 41196 3884 41202 3896
rect 41874 3884 41880 3896
rect 41932 3884 41938 3936
rect 42426 3884 42432 3936
rect 42484 3924 42490 3936
rect 44450 3924 44456 3936
rect 42484 3896 44456 3924
rect 42484 3884 42490 3896
rect 44450 3884 44456 3896
rect 44508 3884 44514 3936
rect 45738 3884 45744 3936
rect 45796 3884 45802 3936
rect 47670 3884 47676 3936
rect 47728 3924 47734 3936
rect 47949 3927 48007 3933
rect 47949 3924 47961 3927
rect 47728 3896 47961 3924
rect 47728 3884 47734 3896
rect 47949 3893 47961 3896
rect 47995 3924 48007 3927
rect 48406 3924 48412 3936
rect 47995 3896 48412 3924
rect 47995 3893 48007 3896
rect 47949 3887 48007 3893
rect 48406 3884 48412 3896
rect 48464 3884 48470 3936
rect 66714 3884 66720 3936
rect 66772 3884 66778 3936
rect 92753 3927 92811 3933
rect 92753 3893 92765 3927
rect 92799 3924 92811 3927
rect 93302 3924 93308 3936
rect 92799 3896 93308 3924
rect 92799 3893 92811 3896
rect 92753 3887 92811 3893
rect 93302 3884 93308 3896
rect 93360 3884 93366 3936
rect 95234 3884 95240 3936
rect 95292 3924 95298 3936
rect 97920 3924 97948 3964
rect 102870 3952 102876 4004
rect 102928 3992 102934 4004
rect 102928 3964 104940 3992
rect 102928 3952 102934 3964
rect 95292 3896 97948 3924
rect 95292 3884 95298 3896
rect 100202 3884 100208 3936
rect 100260 3924 100266 3936
rect 104158 3924 104164 3936
rect 100260 3896 104164 3924
rect 100260 3884 100266 3896
rect 104158 3884 104164 3896
rect 104216 3884 104222 3936
rect 104342 3884 104348 3936
rect 104400 3924 104406 3936
rect 104805 3927 104863 3933
rect 104805 3924 104817 3927
rect 104400 3896 104817 3924
rect 104400 3884 104406 3896
rect 104805 3893 104817 3896
rect 104851 3893 104863 3927
rect 104912 3924 104940 3964
rect 105262 3952 105268 4004
rect 105320 3952 105326 4004
rect 108758 3992 108764 4004
rect 105372 3964 108764 3992
rect 105372 3924 105400 3964
rect 108758 3952 108764 3964
rect 108816 3952 108822 4004
rect 104912 3896 105400 3924
rect 104805 3887 104863 3893
rect 105446 3884 105452 3936
rect 105504 3924 105510 3936
rect 107838 3924 107844 3936
rect 105504 3896 107844 3924
rect 105504 3884 105510 3896
rect 107838 3884 107844 3896
rect 107896 3884 107902 3936
rect 108850 3884 108856 3936
rect 108908 3884 108914 3936
rect 109037 3927 109095 3933
rect 109037 3893 109049 3927
rect 109083 3924 109095 3927
rect 109310 3924 109316 3936
rect 109083 3896 109316 3924
rect 109083 3893 109095 3896
rect 109037 3887 109095 3893
rect 109310 3884 109316 3896
rect 109368 3884 109374 3936
rect 109420 3924 109448 4032
rect 110506 4020 110512 4032
rect 110564 4020 110570 4072
rect 110782 4020 110788 4072
rect 110840 4060 110846 4072
rect 111150 4060 111156 4072
rect 110840 4032 111156 4060
rect 110840 4020 110846 4032
rect 111150 4020 111156 4032
rect 111208 4020 111214 4072
rect 111610 4020 111616 4072
rect 111668 4020 111674 4072
rect 111794 4020 111800 4072
rect 111852 4020 111858 4072
rect 111978 4020 111984 4072
rect 112036 4060 112042 4072
rect 112073 4063 112131 4069
rect 112073 4060 112085 4063
rect 112036 4032 112085 4060
rect 112036 4020 112042 4032
rect 112073 4029 112085 4032
rect 112119 4060 112131 4063
rect 114554 4060 114560 4072
rect 112119 4032 114560 4060
rect 112119 4029 112131 4032
rect 112073 4023 112131 4029
rect 114554 4020 114560 4032
rect 114612 4020 114618 4072
rect 114738 4020 114744 4072
rect 114796 4020 114802 4072
rect 114925 4063 114983 4069
rect 114925 4029 114937 4063
rect 114971 4029 114983 4063
rect 114925 4023 114983 4029
rect 116581 4063 116639 4069
rect 116581 4029 116593 4063
rect 116627 4029 116639 4063
rect 116581 4023 116639 4029
rect 109589 3995 109647 4001
rect 109589 3961 109601 3995
rect 109635 3992 109647 3995
rect 112162 3992 112168 4004
rect 109635 3964 112168 3992
rect 109635 3961 109647 3964
rect 109589 3955 109647 3961
rect 112162 3952 112168 3964
rect 112220 3952 112226 4004
rect 114005 3995 114063 4001
rect 114005 3961 114017 3995
rect 114051 3992 114063 3995
rect 114940 3992 114968 4023
rect 114051 3964 114968 3992
rect 114051 3961 114063 3964
rect 114005 3955 114063 3961
rect 109770 3924 109776 3936
rect 109420 3896 109776 3924
rect 109770 3884 109776 3896
rect 109828 3924 109834 3936
rect 110322 3924 110328 3936
rect 109828 3896 110328 3924
rect 109828 3884 109834 3896
rect 110322 3884 110328 3896
rect 110380 3924 110386 3936
rect 110601 3927 110659 3933
rect 110601 3924 110613 3927
rect 110380 3896 110613 3924
rect 110380 3884 110386 3896
rect 110601 3893 110613 3896
rect 110647 3924 110659 3927
rect 111702 3924 111708 3936
rect 110647 3896 111708 3924
rect 110647 3893 110659 3896
rect 110601 3887 110659 3893
rect 111702 3884 111708 3896
rect 111760 3884 111766 3936
rect 116596 3924 116624 4023
rect 117222 4020 117228 4072
rect 117280 4020 117286 4072
rect 117332 4060 117360 4100
rect 118234 4088 118240 4140
rect 118292 4088 118298 4140
rect 120442 4088 120448 4140
rect 120500 4088 120506 4140
rect 120813 4131 120871 4137
rect 120813 4097 120825 4131
rect 120859 4128 120871 4131
rect 120994 4128 121000 4140
rect 120859 4100 121000 4128
rect 120859 4097 120871 4100
rect 120813 4091 120871 4097
rect 120994 4088 121000 4100
rect 121052 4088 121058 4140
rect 117685 4063 117743 4069
rect 117685 4060 117697 4063
rect 117332 4032 117697 4060
rect 117685 4029 117697 4032
rect 117731 4029 117743 4063
rect 117685 4023 117743 4029
rect 117958 4020 117964 4072
rect 118016 4020 118022 4072
rect 118050 4020 118056 4072
rect 118108 4069 118114 4072
rect 118108 4063 118136 4069
rect 118124 4029 118136 4063
rect 118108 4023 118136 4029
rect 118108 4020 118114 4023
rect 121454 4020 121460 4072
rect 121512 4020 121518 4072
rect 121641 4063 121699 4069
rect 121641 4029 121653 4063
rect 121687 4060 121699 4063
rect 122466 4060 122472 4072
rect 121687 4032 122472 4060
rect 121687 4029 121699 4032
rect 121641 4023 121699 4029
rect 122466 4020 122472 4032
rect 122524 4020 122530 4072
rect 123297 4063 123355 4069
rect 123297 4029 123309 4063
rect 123343 4060 123355 4063
rect 123343 4032 128354 4060
rect 123343 4029 123355 4032
rect 123297 4023 123355 4029
rect 120258 3992 120264 4004
rect 118666 3964 120264 3992
rect 118666 3924 118694 3964
rect 120258 3952 120264 3964
rect 120316 3952 120322 4004
rect 120997 3995 121055 4001
rect 120997 3961 121009 3995
rect 121043 3992 121055 3995
rect 121914 3992 121920 4004
rect 121043 3964 121920 3992
rect 121043 3961 121055 3964
rect 120997 3955 121055 3961
rect 121914 3952 121920 3964
rect 121972 3952 121978 4004
rect 122006 3952 122012 4004
rect 122064 3992 122070 4004
rect 123312 3992 123340 4023
rect 122064 3964 123340 3992
rect 128326 3992 128354 4032
rect 137296 3992 137324 4168
rect 138842 4156 138848 4208
rect 138900 4196 138906 4208
rect 141142 4196 141148 4208
rect 138900 4168 141148 4196
rect 138900 4156 138906 4168
rect 141142 4156 141148 4168
rect 141200 4156 141206 4208
rect 142706 4156 142712 4208
rect 142764 4196 142770 4208
rect 142764 4168 145052 4196
rect 142764 4156 142770 4168
rect 138385 4131 138443 4137
rect 138385 4097 138397 4131
rect 138431 4128 138443 4131
rect 139394 4128 139400 4140
rect 138431 4100 139400 4128
rect 138431 4097 138443 4100
rect 138385 4091 138443 4097
rect 139394 4088 139400 4100
rect 139452 4088 139458 4140
rect 141878 4088 141884 4140
rect 141936 4128 141942 4140
rect 142801 4131 142859 4137
rect 142801 4128 142813 4131
rect 141936 4100 142813 4128
rect 141936 4088 141942 4100
rect 142801 4097 142813 4100
rect 142847 4128 142859 4131
rect 142982 4128 142988 4140
rect 142847 4100 142988 4128
rect 142847 4097 142859 4100
rect 142801 4091 142859 4097
rect 142982 4088 142988 4100
rect 143040 4128 143046 4140
rect 145024 4137 145052 4168
rect 145098 4156 145104 4208
rect 145156 4196 145162 4208
rect 147646 4196 147674 4236
rect 148410 4224 148416 4276
rect 148468 4264 148474 4276
rect 148505 4267 148563 4273
rect 148505 4264 148517 4267
rect 148468 4236 148517 4264
rect 148468 4224 148474 4236
rect 148505 4233 148517 4236
rect 148551 4233 148563 4267
rect 148505 4227 148563 4233
rect 150986 4224 150992 4276
rect 151044 4264 151050 4276
rect 153838 4264 153844 4276
rect 151044 4236 153844 4264
rect 151044 4224 151050 4236
rect 153838 4224 153844 4236
rect 153896 4224 153902 4276
rect 155037 4267 155095 4273
rect 155037 4233 155049 4267
rect 155083 4264 155095 4267
rect 155678 4264 155684 4276
rect 155083 4236 155684 4264
rect 155083 4233 155095 4236
rect 155037 4227 155095 4233
rect 155678 4224 155684 4236
rect 155736 4224 155742 4276
rect 165982 4224 165988 4276
rect 166040 4264 166046 4276
rect 167270 4264 167276 4276
rect 166040 4236 167276 4264
rect 166040 4224 166046 4236
rect 167270 4224 167276 4236
rect 167328 4224 167334 4276
rect 167362 4224 167368 4276
rect 167420 4264 167426 4276
rect 170858 4264 170864 4276
rect 167420 4236 170864 4264
rect 167420 4224 167426 4236
rect 170858 4224 170864 4236
rect 170916 4224 170922 4276
rect 176654 4224 176660 4276
rect 176712 4264 176718 4276
rect 209314 4264 209320 4276
rect 176712 4236 209320 4264
rect 176712 4224 176718 4236
rect 209314 4224 209320 4236
rect 209372 4224 209378 4276
rect 210142 4224 210148 4276
rect 210200 4264 210206 4276
rect 215938 4264 215944 4276
rect 210200 4236 215944 4264
rect 210200 4224 210206 4236
rect 150342 4196 150348 4208
rect 145156 4168 145880 4196
rect 147646 4168 150348 4196
rect 145156 4156 145162 4168
rect 143813 4131 143871 4137
rect 143813 4128 143825 4131
rect 143040 4100 143825 4128
rect 143040 4088 143046 4100
rect 143813 4097 143825 4100
rect 143859 4097 143871 4131
rect 143813 4091 143871 4097
rect 145009 4131 145067 4137
rect 145009 4097 145021 4131
rect 145055 4097 145067 4131
rect 145852 4128 145880 4168
rect 150342 4156 150348 4168
rect 150400 4156 150406 4208
rect 152826 4196 152832 4208
rect 150728 4168 152832 4196
rect 145852 4100 146064 4128
rect 145009 4091 145067 4097
rect 138661 4063 138719 4069
rect 138661 4029 138673 4063
rect 138707 4060 138719 4063
rect 139026 4060 139032 4072
rect 138707 4032 139032 4060
rect 138707 4029 138719 4032
rect 138661 4023 138719 4029
rect 139026 4020 139032 4032
rect 139084 4060 139090 4072
rect 139673 4063 139731 4069
rect 139673 4060 139685 4063
rect 139084 4032 139685 4060
rect 139084 4020 139090 4032
rect 139673 4029 139685 4032
rect 139719 4060 139731 4063
rect 139762 4060 139768 4072
rect 139719 4032 139768 4060
rect 139719 4029 139731 4032
rect 139673 4023 139731 4029
rect 139762 4020 139768 4032
rect 139820 4020 139826 4072
rect 140501 4063 140559 4069
rect 140501 4029 140513 4063
rect 140547 4029 140559 4063
rect 140501 4023 140559 4029
rect 139486 3992 139492 4004
rect 128326 3964 137324 3992
rect 138768 3964 139492 3992
rect 122064 3952 122070 3964
rect 116596 3896 118694 3924
rect 118881 3927 118939 3933
rect 118881 3893 118893 3927
rect 118927 3924 118939 3927
rect 120074 3924 120080 3936
rect 118927 3896 120080 3924
rect 118927 3893 118939 3896
rect 118881 3887 118939 3893
rect 120074 3884 120080 3896
rect 120132 3884 120138 3936
rect 120813 3927 120871 3933
rect 120813 3893 120825 3927
rect 120859 3924 120871 3927
rect 120902 3924 120908 3936
rect 120859 3896 120908 3924
rect 120859 3893 120871 3896
rect 120813 3887 120871 3893
rect 120902 3884 120908 3896
rect 120960 3884 120966 3936
rect 138768 3933 138796 3964
rect 139486 3952 139492 3964
rect 139544 3992 139550 4004
rect 140516 3992 140544 4023
rect 140682 4020 140688 4072
rect 140740 4020 140746 4072
rect 140958 4020 140964 4072
rect 141016 4020 141022 4072
rect 142522 4020 142528 4072
rect 142580 4060 142586 4072
rect 143077 4063 143135 4069
rect 143077 4060 143089 4063
rect 142580 4032 143089 4060
rect 142580 4020 142586 4032
rect 143077 4029 143089 4032
rect 143123 4060 143135 4063
rect 144089 4063 144147 4069
rect 144089 4060 144101 4063
rect 143123 4032 144101 4060
rect 143123 4029 143135 4032
rect 143077 4023 143135 4029
rect 144089 4029 144101 4032
rect 144135 4029 144147 4063
rect 144089 4023 144147 4029
rect 144730 4020 144736 4072
rect 144788 4060 144794 4072
rect 145653 4063 145711 4069
rect 145653 4060 145665 4063
rect 144788 4032 145665 4060
rect 144788 4020 144794 4032
rect 145653 4029 145665 4032
rect 145699 4029 145711 4063
rect 145653 4023 145711 4029
rect 145834 4020 145840 4072
rect 145892 4020 145898 4072
rect 146036 4060 146064 4100
rect 146846 4088 146852 4140
rect 146904 4088 146910 4140
rect 147490 4088 147496 4140
rect 147548 4088 147554 4140
rect 147950 4088 147956 4140
rect 148008 4128 148014 4140
rect 148965 4131 149023 4137
rect 148965 4128 148977 4131
rect 148008 4100 148977 4128
rect 148008 4088 148014 4100
rect 148965 4097 148977 4100
rect 149011 4128 149023 4131
rect 149146 4128 149152 4140
rect 149011 4100 149152 4128
rect 149011 4097 149023 4100
rect 148965 4091 149023 4097
rect 149146 4088 149152 4100
rect 149204 4088 149210 4140
rect 150253 4131 150311 4137
rect 150253 4097 150265 4131
rect 150299 4128 150311 4131
rect 150728 4128 150756 4168
rect 152826 4156 152832 4168
rect 152884 4156 152890 4208
rect 154942 4156 154948 4208
rect 155000 4156 155006 4208
rect 156230 4156 156236 4208
rect 156288 4196 156294 4208
rect 160278 4196 160284 4208
rect 156288 4168 160284 4196
rect 156288 4156 156294 4168
rect 160278 4156 160284 4168
rect 160336 4156 160342 4208
rect 161290 4156 161296 4208
rect 161348 4196 161354 4208
rect 163590 4196 163596 4208
rect 161348 4168 163596 4196
rect 161348 4156 161354 4168
rect 163590 4156 163596 4168
rect 163648 4156 163654 4208
rect 167178 4156 167184 4208
rect 167236 4196 167242 4208
rect 168006 4196 168012 4208
rect 167236 4168 168012 4196
rect 167236 4156 167242 4168
rect 168006 4156 168012 4168
rect 168064 4156 168070 4208
rect 205634 4156 205640 4208
rect 205692 4196 205698 4208
rect 205821 4199 205879 4205
rect 205821 4196 205833 4199
rect 205692 4168 205833 4196
rect 205692 4156 205698 4168
rect 205821 4165 205833 4168
rect 205867 4196 205879 4199
rect 215570 4196 215576 4208
rect 205867 4168 215576 4196
rect 205867 4165 205879 4168
rect 205821 4159 205879 4165
rect 215570 4156 215576 4168
rect 215628 4156 215634 4208
rect 215772 4205 215800 4236
rect 215938 4224 215944 4236
rect 215996 4224 216002 4276
rect 216766 4224 216772 4276
rect 216824 4264 216830 4276
rect 220906 4264 220912 4276
rect 216824 4236 220912 4264
rect 216824 4224 216830 4236
rect 220906 4224 220912 4236
rect 220964 4224 220970 4276
rect 220998 4224 221004 4276
rect 221056 4264 221062 4276
rect 221056 4236 222332 4264
rect 221056 4224 221062 4236
rect 215757 4199 215815 4205
rect 215757 4165 215769 4199
rect 215803 4165 215815 4199
rect 215757 4159 215815 4165
rect 216306 4156 216312 4208
rect 216364 4196 216370 4208
rect 216677 4199 216735 4205
rect 216677 4196 216689 4199
rect 216364 4168 216689 4196
rect 216364 4156 216370 4168
rect 216677 4165 216689 4168
rect 216723 4165 216735 4199
rect 217045 4199 217103 4205
rect 217045 4196 217057 4199
rect 216677 4159 216735 4165
rect 216784 4168 217057 4196
rect 150299 4100 150756 4128
rect 150299 4097 150311 4100
rect 150253 4091 150311 4097
rect 150802 4088 150808 4140
rect 150860 4088 150866 4140
rect 153194 4088 153200 4140
rect 153252 4088 153258 4140
rect 146202 4060 146208 4072
rect 146036 4032 146208 4060
rect 146202 4020 146208 4032
rect 146260 4060 146266 4072
rect 146297 4063 146355 4069
rect 146297 4060 146309 4063
rect 146260 4032 146309 4060
rect 146260 4020 146266 4032
rect 146297 4029 146309 4032
rect 146343 4029 146355 4063
rect 146573 4063 146631 4069
rect 146573 4060 146585 4063
rect 146297 4023 146355 4029
rect 146404 4032 146585 4060
rect 142154 3992 142160 4004
rect 139544 3964 139624 3992
rect 140516 3964 142160 3992
rect 139544 3952 139550 3964
rect 138753 3927 138811 3933
rect 138753 3893 138765 3927
rect 138799 3893 138811 3927
rect 138753 3887 138811 3893
rect 138934 3884 138940 3936
rect 138992 3884 138998 3936
rect 139596 3933 139624 3964
rect 142154 3952 142160 3964
rect 142212 3952 142218 4004
rect 142264 3964 143028 3992
rect 139581 3927 139639 3933
rect 139581 3893 139593 3927
rect 139627 3893 139639 3927
rect 139581 3887 139639 3893
rect 139670 3884 139676 3936
rect 139728 3924 139734 3936
rect 139949 3927 140007 3933
rect 139949 3924 139961 3927
rect 139728 3896 139961 3924
rect 139728 3884 139734 3896
rect 139949 3893 139961 3896
rect 139995 3893 140007 3927
rect 139949 3887 140007 3893
rect 140774 3884 140780 3936
rect 140832 3924 140838 3936
rect 142264 3924 142292 3964
rect 140832 3896 142292 3924
rect 140832 3884 140838 3896
rect 142338 3884 142344 3936
rect 142396 3924 142402 3936
rect 142893 3927 142951 3933
rect 142893 3924 142905 3927
rect 142396 3896 142905 3924
rect 142396 3884 142402 3896
rect 142893 3893 142905 3896
rect 142939 3893 142951 3927
rect 143000 3924 143028 3964
rect 143258 3952 143264 4004
rect 143316 3992 143322 4004
rect 144365 3995 144423 4001
rect 144365 3992 144377 3995
rect 143316 3964 144377 3992
rect 143316 3952 143322 3964
rect 144365 3961 144377 3964
rect 144411 3961 144423 3995
rect 144365 3955 144423 3961
rect 143353 3927 143411 3933
rect 143353 3924 143365 3927
rect 143000 3896 143365 3924
rect 142893 3887 142951 3893
rect 143353 3893 143365 3896
rect 143399 3893 143411 3927
rect 143353 3887 143411 3893
rect 143442 3884 143448 3936
rect 143500 3924 143506 3936
rect 143905 3927 143963 3933
rect 143905 3924 143917 3927
rect 143500 3896 143917 3924
rect 143500 3884 143506 3896
rect 143905 3893 143917 3896
rect 143951 3893 143963 3927
rect 143905 3887 143963 3893
rect 144825 3927 144883 3933
rect 144825 3893 144837 3927
rect 144871 3924 144883 3927
rect 145558 3924 145564 3936
rect 144871 3896 145564 3924
rect 144871 3893 144883 3896
rect 144825 3887 144883 3893
rect 145558 3884 145564 3896
rect 145616 3884 145622 3936
rect 146404 3924 146432 4032
rect 146573 4029 146585 4032
rect 146619 4029 146631 4063
rect 146573 4023 146631 4029
rect 146711 4063 146769 4069
rect 146711 4029 146723 4063
rect 146757 4060 146769 4063
rect 148229 4063 148287 4069
rect 146757 4032 148180 4060
rect 146757 4029 146769 4032
rect 146711 4023 146769 4029
rect 147858 3992 147864 4004
rect 147232 3964 147864 3992
rect 147232 3924 147260 3964
rect 147858 3952 147864 3964
rect 147916 3952 147922 4004
rect 148152 3992 148180 4032
rect 148229 4029 148241 4063
rect 148275 4060 148287 4063
rect 149054 4060 149060 4072
rect 148275 4032 149060 4060
rect 148275 4029 148287 4032
rect 148229 4023 148287 4029
rect 149054 4020 149060 4032
rect 149112 4060 149118 4072
rect 149241 4063 149299 4069
rect 149241 4060 149253 4063
rect 149112 4032 149253 4060
rect 149112 4020 149118 4032
rect 149241 4029 149253 4032
rect 149287 4060 149299 4063
rect 149422 4060 149428 4072
rect 149287 4032 149428 4060
rect 149287 4029 149299 4032
rect 149241 4023 149299 4029
rect 149422 4020 149428 4032
rect 149480 4020 149486 4072
rect 150989 4063 151047 4069
rect 150989 4060 151001 4063
rect 150084 4032 151001 4060
rect 149974 3992 149980 4004
rect 148152 3964 149980 3992
rect 149974 3952 149980 3964
rect 150032 3952 150038 4004
rect 150084 4001 150112 4032
rect 150989 4029 151001 4032
rect 151035 4029 151047 4063
rect 150989 4023 151047 4029
rect 151998 4020 152004 4072
rect 152056 4020 152062 4072
rect 153381 4063 153439 4069
rect 153381 4029 153393 4063
rect 153427 4060 153439 4063
rect 153470 4060 153476 4072
rect 153427 4032 153476 4060
rect 153427 4029 153439 4032
rect 153381 4023 153439 4029
rect 153470 4020 153476 4032
rect 153528 4020 153534 4072
rect 153841 4063 153899 4069
rect 153841 4029 153853 4063
rect 153887 4060 153899 4063
rect 153930 4060 153936 4072
rect 153887 4032 153936 4060
rect 153887 4029 153899 4032
rect 153841 4023 153899 4029
rect 153930 4020 153936 4032
rect 153988 4020 153994 4072
rect 154114 4020 154120 4072
rect 154172 4020 154178 4072
rect 154206 4020 154212 4072
rect 154264 4069 154270 4072
rect 154264 4063 154292 4069
rect 154280 4029 154292 4063
rect 154264 4023 154292 4029
rect 154393 4063 154451 4069
rect 154393 4029 154405 4063
rect 154439 4060 154451 4063
rect 154960 4060 154988 4156
rect 164326 4128 164332 4140
rect 159652 4100 164332 4128
rect 154439 4032 154988 4060
rect 154439 4029 154451 4032
rect 154393 4023 154451 4029
rect 154264 4020 154270 4023
rect 155218 4020 155224 4072
rect 155276 4060 155282 4072
rect 155957 4063 156015 4069
rect 155957 4060 155969 4063
rect 155276 4032 155969 4060
rect 155276 4020 155282 4032
rect 155957 4029 155969 4032
rect 156003 4029 156015 4063
rect 155957 4023 156015 4029
rect 156141 4063 156199 4069
rect 156141 4029 156153 4063
rect 156187 4060 156199 4063
rect 156230 4060 156236 4072
rect 156187 4032 156236 4060
rect 156187 4029 156199 4032
rect 156141 4023 156199 4029
rect 156230 4020 156236 4032
rect 156288 4020 156294 4072
rect 157058 4020 157064 4072
rect 157116 4020 157122 4072
rect 158257 4063 158315 4069
rect 158257 4029 158269 4063
rect 158303 4029 158315 4063
rect 158257 4023 158315 4029
rect 150069 3995 150127 4001
rect 150069 3961 150081 3995
rect 150115 3961 150127 3995
rect 150069 3955 150127 3961
rect 152182 3952 152188 4004
rect 152240 3992 152246 4004
rect 152240 3964 152872 3992
rect 152240 3952 152246 3964
rect 146404 3896 147260 3924
rect 147306 3884 147312 3936
rect 147364 3924 147370 3936
rect 148045 3927 148103 3933
rect 148045 3924 148057 3927
rect 147364 3896 148057 3924
rect 147364 3884 147370 3896
rect 148045 3893 148057 3896
rect 148091 3924 148103 3927
rect 149057 3927 149115 3933
rect 149057 3924 149069 3927
rect 148091 3896 149069 3924
rect 148091 3893 148103 3896
rect 148045 3887 148103 3893
rect 149057 3893 149069 3896
rect 149103 3924 149115 3927
rect 149238 3924 149244 3936
rect 149103 3896 149244 3924
rect 149103 3893 149115 3896
rect 149057 3887 149115 3893
rect 149238 3884 149244 3896
rect 149296 3884 149302 3936
rect 149517 3927 149575 3933
rect 149517 3893 149529 3927
rect 149563 3924 149575 3927
rect 152734 3924 152740 3936
rect 149563 3896 152740 3924
rect 149563 3893 149575 3896
rect 149517 3887 149575 3893
rect 152734 3884 152740 3896
rect 152792 3884 152798 3936
rect 152844 3924 152872 3964
rect 154942 3952 154948 4004
rect 155000 3992 155006 4004
rect 158162 3992 158168 4004
rect 155000 3964 158168 3992
rect 155000 3952 155006 3964
rect 158162 3952 158168 3964
rect 158220 3952 158226 4004
rect 158272 3992 158300 4023
rect 158438 4020 158444 4072
rect 158496 4020 158502 4072
rect 158530 4020 158536 4072
rect 158588 4060 158594 4072
rect 159652 4060 159680 4100
rect 164326 4088 164332 4100
rect 164384 4088 164390 4140
rect 167641 4131 167699 4137
rect 167641 4097 167653 4131
rect 167687 4128 167699 4131
rect 167730 4128 167736 4140
rect 167687 4100 167736 4128
rect 167687 4097 167699 4100
rect 167641 4091 167699 4097
rect 167730 4088 167736 4100
rect 167788 4088 167794 4140
rect 168024 4128 168052 4156
rect 168101 4131 168159 4137
rect 168101 4128 168113 4131
rect 168024 4100 168113 4128
rect 168101 4097 168113 4100
rect 168147 4097 168159 4131
rect 168101 4091 168159 4097
rect 190454 4088 190460 4140
rect 190512 4088 190518 4140
rect 206005 4131 206063 4137
rect 206005 4097 206017 4131
rect 206051 4128 206063 4131
rect 206554 4128 206560 4140
rect 206051 4100 206560 4128
rect 206051 4097 206063 4100
rect 206005 4091 206063 4097
rect 206554 4088 206560 4100
rect 206612 4088 206618 4140
rect 206646 4088 206652 4140
rect 206704 4088 206710 4140
rect 206738 4088 206744 4140
rect 206796 4088 206802 4140
rect 213178 4088 213184 4140
rect 213236 4088 213242 4140
rect 158588 4032 159680 4060
rect 158588 4020 158594 4032
rect 160002 4020 160008 4072
rect 160060 4020 160066 4072
rect 168009 4063 168067 4069
rect 168009 4029 168021 4063
rect 168055 4060 168067 4063
rect 168190 4060 168196 4072
rect 168055 4032 168196 4060
rect 168055 4029 168067 4032
rect 168009 4023 168067 4029
rect 168190 4020 168196 4032
rect 168248 4020 168254 4072
rect 176626 4032 206876 4060
rect 160370 3992 160376 4004
rect 158272 3964 160376 3992
rect 160370 3952 160376 3964
rect 160428 3952 160434 4004
rect 161382 3952 161388 4004
rect 161440 3992 161446 4004
rect 176626 3992 176654 4032
rect 161440 3964 176654 3992
rect 161440 3952 161446 3964
rect 154574 3924 154580 3936
rect 152844 3896 154580 3924
rect 154574 3884 154580 3896
rect 154632 3884 154638 3936
rect 158530 3884 158536 3936
rect 158588 3924 158594 3936
rect 164234 3924 164240 3936
rect 158588 3896 164240 3924
rect 158588 3884 158594 3896
rect 164234 3884 164240 3896
rect 164292 3884 164298 3936
rect 164326 3884 164332 3936
rect 164384 3924 164390 3936
rect 167362 3924 167368 3936
rect 164384 3896 167368 3924
rect 164384 3884 164390 3896
rect 167362 3884 167368 3896
rect 167420 3884 167426 3936
rect 167454 3884 167460 3936
rect 167512 3924 167518 3936
rect 167733 3927 167791 3933
rect 167733 3924 167745 3927
rect 167512 3896 167745 3924
rect 167512 3884 167518 3896
rect 167733 3893 167745 3896
rect 167779 3893 167791 3927
rect 167733 3887 167791 3893
rect 168282 3884 168288 3936
rect 168340 3884 168346 3936
rect 190273 3927 190331 3933
rect 190273 3893 190285 3927
rect 190319 3924 190331 3927
rect 191190 3924 191196 3936
rect 190319 3896 191196 3924
rect 190319 3893 190331 3896
rect 190273 3887 190331 3893
rect 191190 3884 191196 3896
rect 191248 3884 191254 3936
rect 206848 3924 206876 4032
rect 207474 4020 207480 4072
rect 207532 4020 207538 4072
rect 207661 4063 207719 4069
rect 207661 4029 207673 4063
rect 207707 4029 207719 4063
rect 207661 4023 207719 4029
rect 206925 3995 206983 4001
rect 206925 3961 206937 3995
rect 206971 3992 206983 3995
rect 207676 3992 207704 4023
rect 209314 4020 209320 4072
rect 209372 4020 209378 4072
rect 209774 4020 209780 4072
rect 209832 4020 209838 4072
rect 209958 4020 209964 4072
rect 210016 4020 210022 4072
rect 210237 4063 210295 4069
rect 210237 4029 210249 4063
rect 210283 4029 210295 4063
rect 210237 4023 210295 4029
rect 206971 3964 207704 3992
rect 206971 3961 206983 3964
rect 206925 3955 206983 3961
rect 208302 3952 208308 4004
rect 208360 3992 208366 4004
rect 209222 3992 209228 4004
rect 208360 3964 209228 3992
rect 208360 3952 208366 3964
rect 209222 3952 209228 3964
rect 209280 3952 209286 4004
rect 210252 3992 210280 4023
rect 212074 4020 212080 4072
rect 212132 4060 212138 4072
rect 213365 4063 213423 4069
rect 213365 4060 213377 4063
rect 212132 4032 213377 4060
rect 212132 4020 212138 4032
rect 213365 4029 213377 4032
rect 213411 4029 213423 4063
rect 213365 4023 213423 4029
rect 213914 4020 213920 4072
rect 213972 4060 213978 4072
rect 216582 4060 216588 4072
rect 213972 4032 216588 4060
rect 213972 4020 213978 4032
rect 216582 4020 216588 4032
rect 216640 4020 216646 4072
rect 216674 4020 216680 4072
rect 216732 4060 216738 4072
rect 216784 4060 216812 4168
rect 217045 4165 217057 4168
rect 217091 4196 217103 4199
rect 217870 4196 217876 4208
rect 217091 4168 217876 4196
rect 217091 4165 217103 4168
rect 217045 4159 217103 4165
rect 217870 4156 217876 4168
rect 217928 4156 217934 4208
rect 216950 4088 216956 4140
rect 217008 4128 217014 4140
rect 217965 4131 218023 4137
rect 217965 4128 217977 4131
rect 217008 4100 217977 4128
rect 217008 4088 217014 4100
rect 217965 4097 217977 4100
rect 218011 4097 218023 4131
rect 217965 4091 218023 4097
rect 220262 4088 220268 4140
rect 220320 4088 220326 4140
rect 222304 4128 222332 4236
rect 223298 4224 223304 4276
rect 223356 4264 223362 4276
rect 223356 4236 224954 4264
rect 223356 4224 223362 4236
rect 224926 4196 224954 4236
rect 225138 4224 225144 4276
rect 225196 4264 225202 4276
rect 242986 4264 242992 4276
rect 225196 4236 242992 4264
rect 225196 4224 225202 4236
rect 242986 4224 242992 4236
rect 243044 4224 243050 4276
rect 244369 4267 244427 4273
rect 244369 4233 244381 4267
rect 244415 4233 244427 4267
rect 244369 4227 244427 4233
rect 226978 4196 226984 4208
rect 224926 4168 226984 4196
rect 226978 4156 226984 4168
rect 227036 4156 227042 4208
rect 222933 4131 222991 4137
rect 222933 4128 222945 4131
rect 222304 4100 222945 4128
rect 222933 4097 222945 4100
rect 222979 4097 222991 4131
rect 223853 4131 223911 4137
rect 223853 4106 223865 4131
rect 223899 4106 223911 4131
rect 223991 4131 224049 4137
rect 222933 4091 222991 4097
rect 216732 4032 216812 4060
rect 216732 4020 216738 4032
rect 217686 4020 217692 4072
rect 217744 4060 217750 4072
rect 217781 4063 217839 4069
rect 217781 4060 217793 4063
rect 217744 4032 217793 4060
rect 217744 4020 217750 4032
rect 217781 4029 217793 4032
rect 217827 4029 217839 4063
rect 217781 4023 217839 4029
rect 218146 4020 218152 4072
rect 218204 4060 218210 4072
rect 218422 4060 218428 4072
rect 218204 4032 218428 4060
rect 218204 4020 218210 4032
rect 218422 4020 218428 4032
rect 218480 4020 218486 4072
rect 218698 4020 218704 4072
rect 218756 4020 218762 4072
rect 218790 4020 218796 4072
rect 218848 4069 218854 4072
rect 218848 4063 218876 4069
rect 218864 4029 218876 4063
rect 218848 4023 218876 4029
rect 218848 4020 218854 4023
rect 218974 4020 218980 4072
rect 219032 4060 219038 4072
rect 219158 4060 219164 4072
rect 219032 4032 219164 4060
rect 219032 4020 219038 4032
rect 219158 4020 219164 4032
rect 219216 4020 219222 4072
rect 219342 4020 219348 4072
rect 219400 4060 219406 4072
rect 220081 4063 220139 4069
rect 220081 4060 220093 4063
rect 219400 4032 220093 4060
rect 219400 4020 219406 4032
rect 220081 4029 220093 4032
rect 220127 4029 220139 4063
rect 220081 4023 220139 4029
rect 220998 4020 221004 4072
rect 221056 4020 221062 4072
rect 221182 4069 221188 4072
rect 221139 4063 221188 4069
rect 221139 4029 221151 4063
rect 221185 4029 221188 4063
rect 221139 4023 221188 4029
rect 221182 4020 221188 4023
rect 221240 4020 221246 4072
rect 221277 4063 221335 4069
rect 221277 4029 221289 4063
rect 221323 4060 221335 4063
rect 221918 4060 221924 4072
rect 221323 4032 221924 4060
rect 221323 4029 221335 4032
rect 221277 4023 221335 4029
rect 221918 4020 221924 4032
rect 221976 4060 221982 4072
rect 222286 4060 222292 4072
rect 221976 4032 222292 4060
rect 221976 4020 221982 4032
rect 222286 4020 222292 4032
rect 222344 4020 222350 4072
rect 223117 4063 223175 4069
rect 223117 4029 223129 4063
rect 223163 4060 223175 4063
rect 223298 4060 223304 4072
rect 223163 4032 223304 4060
rect 223163 4029 223175 4032
rect 223117 4023 223175 4029
rect 223298 4020 223304 4032
rect 223356 4020 223362 4072
rect 223574 4020 223580 4072
rect 223632 4020 223638 4072
rect 223850 4054 223856 4106
rect 223908 4054 223914 4106
rect 223991 4097 224003 4131
rect 224037 4097 224049 4131
rect 223991 4091 224049 4097
rect 224006 4060 224034 4091
rect 224126 4088 224132 4140
rect 224184 4088 224190 4140
rect 224770 4088 224776 4140
rect 224828 4088 224834 4140
rect 227254 4088 227260 4140
rect 227312 4128 227318 4140
rect 236549 4131 236607 4137
rect 236549 4128 236561 4131
rect 227312 4100 236561 4128
rect 227312 4088 227318 4100
rect 236549 4097 236561 4100
rect 236595 4097 236607 4131
rect 236549 4091 236607 4097
rect 225233 4063 225291 4069
rect 224006 4032 225184 4060
rect 211798 3992 211804 4004
rect 209608 3964 211804 3992
rect 209608 3924 209636 3964
rect 211798 3952 211804 3964
rect 211856 3952 211862 4004
rect 213178 3952 213184 4004
rect 213236 3992 213242 4004
rect 215294 3992 215300 4004
rect 213236 3964 215300 3992
rect 213236 3952 213242 3964
rect 215294 3952 215300 3964
rect 215352 3952 215358 4004
rect 217962 3992 217968 4004
rect 215956 3964 217968 3992
rect 206848 3896 209636 3924
rect 209682 3884 209688 3936
rect 209740 3924 209746 3936
rect 215956 3924 215984 3964
rect 217962 3952 217968 3964
rect 218020 3952 218026 4004
rect 219802 3952 219808 4004
rect 219860 3992 219866 4004
rect 220354 3992 220360 4004
rect 219860 3964 220360 3992
rect 219860 3952 219866 3964
rect 220354 3952 220360 3964
rect 220412 3992 220418 4004
rect 220722 3992 220728 4004
rect 220412 3964 220728 3992
rect 220412 3952 220418 3964
rect 220722 3952 220728 3964
rect 220780 3952 220786 4004
rect 209740 3896 215984 3924
rect 209740 3884 209746 3896
rect 216030 3884 216036 3936
rect 216088 3884 216094 3936
rect 217410 3884 217416 3936
rect 217468 3924 217474 3936
rect 219621 3927 219679 3933
rect 219621 3924 219633 3927
rect 217468 3896 219633 3924
rect 217468 3884 217474 3896
rect 219621 3893 219633 3896
rect 219667 3893 219679 3927
rect 219621 3887 219679 3893
rect 221090 3884 221096 3936
rect 221148 3924 221154 3936
rect 221921 3927 221979 3933
rect 221921 3924 221933 3927
rect 221148 3896 221933 3924
rect 221148 3884 221154 3896
rect 221921 3893 221933 3896
rect 221967 3893 221979 3927
rect 221921 3887 221979 3893
rect 222102 3884 222108 3936
rect 222160 3924 222166 3936
rect 224770 3924 224776 3936
rect 222160 3896 224776 3924
rect 222160 3884 222166 3896
rect 224770 3884 224776 3896
rect 224828 3884 224834 3936
rect 225156 3933 225184 4032
rect 225233 4029 225245 4063
rect 225279 4029 225291 4063
rect 225233 4023 225291 4029
rect 225248 3992 225276 4023
rect 225414 4020 225420 4072
rect 225472 4020 225478 4072
rect 226702 4020 226708 4072
rect 226760 4020 226766 4072
rect 227622 4020 227628 4072
rect 227680 4060 227686 4072
rect 229830 4060 229836 4072
rect 227680 4032 229836 4060
rect 227680 4020 227686 4032
rect 229830 4020 229836 4032
rect 229888 4020 229894 4072
rect 236825 4063 236883 4069
rect 236825 4029 236837 4063
rect 236871 4060 236883 4063
rect 242894 4060 242900 4072
rect 236871 4032 242900 4060
rect 236871 4029 236883 4032
rect 236825 4023 236883 4029
rect 242894 4020 242900 4032
rect 242952 4020 242958 4072
rect 244384 4060 244412 4227
rect 247034 4224 247040 4276
rect 247092 4264 247098 4276
rect 247092 4236 258028 4264
rect 247092 4224 247098 4236
rect 244936 4168 246436 4196
rect 244553 4131 244611 4137
rect 244553 4097 244565 4131
rect 244599 4128 244611 4131
rect 244936 4128 244964 4168
rect 244599 4100 244964 4128
rect 244599 4097 244611 4100
rect 244553 4091 244611 4097
rect 245010 4088 245016 4140
rect 245068 4137 245074 4140
rect 245068 4091 245076 4137
rect 246408 4128 246436 4168
rect 246850 4156 246856 4208
rect 246908 4196 246914 4208
rect 246908 4168 247632 4196
rect 246908 4156 246914 4168
rect 247604 4140 247632 4168
rect 251266 4156 251272 4208
rect 251324 4196 251330 4208
rect 251324 4168 252508 4196
rect 251324 4156 251330 4168
rect 247126 4128 247132 4140
rect 246408 4100 247132 4128
rect 245068 4088 245074 4091
rect 247126 4088 247132 4100
rect 247184 4088 247190 4140
rect 247218 4088 247224 4140
rect 247276 4128 247282 4140
rect 247313 4131 247371 4137
rect 247313 4128 247325 4131
rect 247276 4100 247325 4128
rect 247276 4088 247282 4100
rect 247313 4097 247325 4100
rect 247359 4097 247371 4131
rect 247313 4091 247371 4097
rect 247586 4088 247592 4140
rect 247644 4088 247650 4140
rect 250990 4088 250996 4140
rect 251048 4088 251054 4140
rect 252480 4128 252508 4168
rect 252554 4156 252560 4208
rect 252612 4196 252618 4208
rect 252833 4199 252891 4205
rect 252833 4196 252845 4199
rect 252612 4168 252845 4196
rect 252612 4156 252618 4168
rect 252833 4165 252845 4168
rect 252879 4196 252891 4199
rect 252879 4168 253796 4196
rect 252879 4165 252891 4168
rect 252833 4159 252891 4165
rect 252646 4128 252652 4140
rect 252480 4100 252652 4128
rect 252646 4088 252652 4100
rect 252704 4088 252710 4140
rect 252922 4088 252928 4140
rect 252980 4128 252986 4140
rect 253109 4131 253167 4137
rect 253109 4128 253121 4131
rect 252980 4100 253121 4128
rect 252980 4088 252986 4100
rect 253109 4097 253121 4100
rect 253155 4128 253167 4131
rect 253658 4128 253664 4140
rect 253155 4100 253664 4128
rect 253155 4097 253167 4100
rect 253109 4091 253167 4097
rect 253658 4088 253664 4100
rect 253716 4088 253722 4140
rect 253768 4128 253796 4168
rect 253842 4156 253848 4208
rect 253900 4196 253906 4208
rect 257890 4196 257896 4208
rect 253900 4168 254440 4196
rect 253900 4156 253906 4168
rect 254118 4128 254124 4140
rect 253768 4100 254124 4128
rect 254118 4088 254124 4100
rect 254176 4088 254182 4140
rect 254412 4137 254440 4168
rect 257264 4168 257896 4196
rect 254397 4131 254455 4137
rect 254397 4097 254409 4131
rect 254443 4097 254455 4131
rect 254397 4091 254455 4097
rect 256881 4131 256939 4137
rect 256881 4097 256893 4131
rect 256927 4128 256939 4131
rect 257264 4128 257292 4168
rect 257890 4156 257896 4168
rect 257948 4156 257954 4208
rect 258000 4196 258028 4236
rect 258258 4224 258264 4276
rect 258316 4264 258322 4276
rect 266262 4264 266268 4276
rect 258316 4236 266268 4264
rect 258316 4224 258322 4236
rect 266262 4224 266268 4236
rect 266320 4224 266326 4276
rect 266446 4224 266452 4276
rect 266504 4264 266510 4276
rect 267277 4267 267335 4273
rect 267277 4264 267289 4267
rect 266504 4236 267289 4264
rect 266504 4224 266510 4236
rect 267277 4233 267289 4236
rect 267323 4233 267335 4267
rect 267277 4227 267335 4233
rect 268562 4224 268568 4276
rect 268620 4224 268626 4276
rect 270770 4224 270776 4276
rect 270828 4224 270834 4276
rect 258534 4196 258540 4208
rect 258000 4168 258540 4196
rect 258534 4156 258540 4168
rect 258592 4156 258598 4208
rect 259822 4156 259828 4208
rect 259880 4156 259886 4208
rect 267734 4196 267740 4208
rect 265820 4168 267740 4196
rect 256927 4100 257292 4128
rect 256927 4097 256939 4100
rect 256881 4091 256939 4097
rect 257338 4088 257344 4140
rect 257396 4088 257402 4140
rect 257430 4088 257436 4140
rect 257488 4128 257494 4140
rect 257525 4131 257583 4137
rect 257525 4128 257537 4131
rect 257488 4100 257537 4128
rect 257488 4088 257494 4100
rect 257525 4097 257537 4100
rect 257571 4097 257583 4131
rect 257525 4091 257583 4097
rect 257614 4088 257620 4140
rect 257672 4088 257678 4140
rect 258445 4131 258503 4137
rect 258445 4128 258457 4131
rect 257724 4100 258457 4128
rect 245197 4063 245255 4069
rect 245197 4060 245209 4063
rect 244384 4032 245209 4060
rect 245197 4029 245209 4032
rect 245243 4029 245255 4063
rect 245197 4023 245255 4029
rect 246853 4063 246911 4069
rect 246853 4029 246865 4063
rect 246899 4060 246911 4063
rect 248414 4060 248420 4072
rect 246899 4032 248420 4060
rect 246899 4029 246911 4032
rect 246853 4023 246911 4029
rect 248414 4020 248420 4032
rect 248472 4020 248478 4072
rect 248690 4020 248696 4072
rect 248748 4020 248754 4072
rect 248877 4063 248935 4069
rect 248877 4029 248889 4063
rect 248923 4060 248935 4063
rect 249426 4060 249432 4072
rect 248923 4032 249432 4060
rect 248923 4029 248935 4032
rect 248877 4023 248935 4029
rect 249426 4020 249432 4032
rect 249484 4020 249490 4072
rect 250533 4063 250591 4069
rect 250533 4029 250545 4063
rect 250579 4060 250591 4063
rect 250806 4060 250812 4072
rect 250579 4032 250812 4060
rect 250579 4029 250591 4032
rect 250533 4023 250591 4029
rect 250806 4020 250812 4032
rect 250864 4020 250870 4072
rect 251269 4063 251327 4069
rect 251269 4029 251281 4063
rect 251315 4060 251327 4063
rect 251358 4060 251364 4072
rect 251315 4032 251364 4060
rect 251315 4029 251327 4032
rect 251269 4023 251327 4029
rect 251358 4020 251364 4032
rect 251416 4020 251422 4072
rect 253014 4020 253020 4072
rect 253072 4060 253078 4072
rect 254305 4063 254363 4069
rect 254305 4060 254317 4063
rect 253072 4032 254317 4060
rect 253072 4020 253078 4032
rect 254305 4029 254317 4032
rect 254351 4060 254363 4063
rect 254578 4060 254584 4072
rect 254351 4032 254584 4060
rect 254351 4029 254363 4032
rect 254305 4023 254363 4029
rect 254578 4020 254584 4032
rect 254636 4020 254642 4072
rect 255041 4063 255099 4069
rect 255041 4029 255053 4063
rect 255087 4029 255099 4063
rect 255041 4023 255099 4029
rect 255225 4063 255283 4069
rect 255225 4029 255237 4063
rect 255271 4060 255283 4063
rect 257062 4060 257068 4072
rect 255271 4032 257068 4060
rect 255271 4029 255283 4032
rect 255225 4023 255283 4029
rect 227346 3992 227352 4004
rect 225248 3964 227352 3992
rect 227346 3952 227352 3964
rect 227404 3952 227410 4004
rect 227438 3952 227444 4004
rect 227496 3992 227502 4004
rect 244182 3992 244188 4004
rect 227496 3964 244188 3992
rect 227496 3952 227502 3964
rect 244182 3952 244188 3964
rect 244240 3952 244246 4004
rect 244458 3952 244464 4004
rect 244516 3992 244522 4004
rect 255056 3992 255084 4023
rect 257062 4020 257068 4032
rect 257120 4020 257126 4072
rect 257724 4060 257752 4100
rect 258445 4097 258457 4100
rect 258491 4097 258503 4131
rect 258445 4091 258503 4097
rect 258997 4131 259055 4137
rect 258997 4097 259009 4131
rect 259043 4097 259055 4131
rect 258997 4091 259055 4097
rect 259012 4060 259040 4091
rect 261754 4088 261760 4140
rect 261812 4128 261818 4140
rect 265161 4131 265219 4137
rect 261812 4100 265020 4128
rect 261812 4088 261818 4100
rect 257172 4032 257752 4060
rect 257816 4032 259040 4060
rect 244516 3964 255084 3992
rect 244516 3952 244522 3964
rect 225141 3927 225199 3933
rect 225141 3893 225153 3927
rect 225187 3924 225199 3927
rect 228174 3924 228180 3936
rect 225187 3896 228180 3924
rect 225187 3893 225199 3896
rect 225141 3887 225199 3893
rect 228174 3884 228180 3896
rect 228232 3884 228238 3936
rect 229738 3884 229744 3936
rect 229796 3924 229802 3936
rect 244274 3924 244280 3936
rect 229796 3896 244280 3924
rect 229796 3884 229802 3896
rect 244274 3884 244280 3896
rect 244332 3884 244338 3936
rect 252830 3884 252836 3936
rect 252888 3884 252894 3936
rect 253293 3927 253351 3933
rect 253293 3893 253305 3927
rect 253339 3924 253351 3927
rect 254026 3924 254032 3936
rect 253339 3896 254032 3924
rect 253339 3893 253351 3896
rect 253293 3887 253351 3893
rect 254026 3884 254032 3896
rect 254084 3884 254090 3936
rect 254118 3884 254124 3936
rect 254176 3884 254182 3936
rect 254581 3927 254639 3933
rect 254581 3893 254593 3927
rect 254627 3924 254639 3927
rect 257172 3924 257200 4032
rect 257816 4001 257844 4032
rect 259270 4020 259276 4072
rect 259328 4060 259334 4072
rect 259641 4063 259699 4069
rect 259641 4060 259653 4063
rect 259328 4032 259653 4060
rect 259328 4020 259334 4032
rect 259641 4029 259653 4032
rect 259687 4029 259699 4063
rect 259641 4023 259699 4029
rect 260742 4020 260748 4072
rect 260800 4020 260806 4072
rect 257801 3995 257859 4001
rect 257801 3961 257813 3995
rect 257847 3961 257859 3995
rect 257801 3955 257859 3961
rect 257890 3952 257896 4004
rect 257948 3992 257954 4004
rect 264992 3992 265020 4100
rect 265161 4097 265173 4131
rect 265207 4128 265219 4131
rect 265526 4128 265532 4140
rect 265207 4100 265532 4128
rect 265207 4097 265219 4100
rect 265161 4091 265219 4097
rect 265526 4088 265532 4100
rect 265584 4088 265590 4140
rect 265820 4137 265848 4168
rect 267734 4156 267740 4168
rect 267792 4156 267798 4208
rect 265805 4131 265863 4137
rect 265805 4097 265817 4131
rect 265851 4097 265863 4131
rect 265805 4091 265863 4097
rect 266449 4131 266507 4137
rect 266449 4097 266461 4131
rect 266495 4128 266507 4131
rect 266906 4128 266912 4140
rect 266495 4100 266912 4128
rect 266495 4097 266507 4100
rect 266449 4091 266507 4097
rect 266906 4088 266912 4100
rect 266964 4088 266970 4140
rect 266998 4088 267004 4140
rect 267056 4088 267062 4140
rect 267090 4088 267096 4140
rect 267148 4128 267154 4140
rect 267921 4131 267979 4137
rect 267921 4128 267933 4131
rect 267148 4100 267933 4128
rect 267148 4088 267154 4100
rect 267921 4097 267933 4100
rect 267967 4097 267979 4131
rect 267921 4091 267979 4097
rect 269298 4088 269304 4140
rect 269356 4088 269362 4140
rect 270037 4131 270095 4137
rect 270037 4097 270049 4131
rect 270083 4128 270095 4131
rect 270862 4128 270868 4140
rect 270083 4100 270868 4128
rect 270083 4097 270095 4100
rect 270037 4091 270095 4097
rect 270862 4088 270868 4100
rect 270920 4088 270926 4140
rect 270957 4131 271015 4137
rect 270957 4097 270969 4131
rect 271003 4128 271015 4131
rect 272058 4128 272064 4140
rect 271003 4100 272064 4128
rect 271003 4097 271015 4100
rect 270957 4091 271015 4097
rect 272058 4088 272064 4100
rect 272116 4088 272122 4140
rect 267274 4020 267280 4072
rect 267332 4060 267338 4072
rect 267737 4063 267795 4069
rect 267737 4060 267749 4063
rect 267332 4032 267749 4060
rect 267332 4020 267338 4032
rect 267737 4029 267749 4032
rect 267783 4029 267795 4063
rect 267737 4023 267795 4029
rect 266265 3995 266323 4001
rect 266265 3992 266277 3995
rect 257948 3964 263594 3992
rect 264992 3964 266277 3992
rect 257948 3952 257954 3964
rect 254627 3896 257200 3924
rect 254627 3893 254639 3896
rect 254581 3887 254639 3893
rect 257338 3884 257344 3936
rect 257396 3884 257402 3936
rect 257430 3884 257436 3936
rect 257488 3924 257494 3936
rect 258261 3927 258319 3933
rect 258261 3924 258273 3927
rect 257488 3896 258273 3924
rect 257488 3884 257494 3896
rect 258261 3893 258273 3896
rect 258307 3893 258319 3927
rect 258261 3887 258319 3893
rect 258810 3884 258816 3936
rect 258868 3884 258874 3936
rect 259270 3884 259276 3936
rect 259328 3884 259334 3936
rect 261754 3884 261760 3936
rect 261812 3924 261818 3936
rect 262030 3924 262036 3936
rect 261812 3896 262036 3924
rect 261812 3884 261818 3896
rect 262030 3884 262036 3896
rect 262088 3884 262094 3936
rect 263566 3924 263594 3964
rect 266265 3961 266277 3964
rect 266311 3961 266323 3995
rect 266265 3955 266323 3961
rect 269482 3952 269488 4004
rect 269540 3952 269546 4004
rect 270221 3995 270279 4001
rect 270221 3961 270233 3995
rect 270267 3992 270279 3995
rect 270494 3992 270500 4004
rect 270267 3964 270500 3992
rect 270267 3961 270279 3964
rect 270221 3955 270279 3961
rect 270494 3952 270500 3964
rect 270552 3952 270558 4004
rect 264790 3924 264796 3936
rect 263566 3896 264796 3924
rect 264790 3884 264796 3896
rect 264848 3884 264854 3936
rect 264977 3927 265035 3933
rect 264977 3893 264989 3927
rect 265023 3924 265035 3927
rect 265802 3924 265808 3936
rect 265023 3896 265808 3924
rect 265023 3893 265035 3896
rect 264977 3887 265035 3893
rect 265802 3884 265808 3896
rect 265860 3884 265866 3936
rect 267734 3884 267740 3936
rect 267792 3924 267798 3936
rect 268105 3927 268163 3933
rect 268105 3924 268117 3927
rect 267792 3896 268117 3924
rect 267792 3884 267798 3896
rect 268105 3893 268117 3896
rect 268151 3893 268163 3927
rect 268105 3887 268163 3893
rect 1104 3834 271492 3856
rect 1104 3782 34748 3834
rect 34800 3782 34812 3834
rect 34864 3782 34876 3834
rect 34928 3782 34940 3834
rect 34992 3782 35004 3834
rect 35056 3782 102345 3834
rect 102397 3782 102409 3834
rect 102461 3782 102473 3834
rect 102525 3782 102537 3834
rect 102589 3782 102601 3834
rect 102653 3782 169942 3834
rect 169994 3782 170006 3834
rect 170058 3782 170070 3834
rect 170122 3782 170134 3834
rect 170186 3782 170198 3834
rect 170250 3782 237539 3834
rect 237591 3782 237603 3834
rect 237655 3782 237667 3834
rect 237719 3782 237731 3834
rect 237783 3782 237795 3834
rect 237847 3782 271492 3834
rect 1104 3760 271492 3782
rect 44450 3680 44456 3732
rect 44508 3720 44514 3732
rect 48130 3720 48136 3732
rect 44508 3692 48136 3720
rect 44508 3680 44514 3692
rect 48130 3680 48136 3692
rect 48188 3680 48194 3732
rect 92474 3720 92480 3732
rect 80026 3692 92480 3720
rect 67634 3612 67640 3664
rect 67692 3652 67698 3664
rect 68833 3655 68891 3661
rect 68833 3652 68845 3655
rect 67692 3624 68845 3652
rect 67692 3612 67698 3624
rect 68833 3621 68845 3624
rect 68879 3621 68891 3655
rect 68833 3615 68891 3621
rect 37372 3596 37424 3602
rect 38470 3584 38476 3596
rect 37424 3556 38476 3584
rect 38470 3544 38476 3556
rect 38528 3544 38534 3596
rect 42518 3584 42524 3596
rect 41814 3556 42524 3584
rect 37372 3538 37424 3544
rect 23198 3476 23204 3528
rect 23256 3516 23262 3528
rect 23385 3519 23443 3525
rect 23385 3516 23397 3519
rect 23256 3488 23397 3516
rect 23256 3476 23262 3488
rect 23385 3485 23397 3488
rect 23431 3485 23443 3519
rect 23385 3479 23443 3485
rect 36630 3476 36636 3528
rect 36688 3476 36694 3528
rect 36814 3476 36820 3528
rect 36872 3516 36878 3528
rect 37093 3519 37151 3525
rect 37093 3516 37105 3519
rect 36872 3488 37105 3516
rect 36872 3476 36878 3488
rect 37093 3485 37105 3488
rect 37139 3485 37151 3519
rect 37274 3516 37280 3528
rect 37093 3479 37151 3485
rect 37200 3488 37280 3516
rect 7374 3408 7380 3460
rect 7432 3448 7438 3460
rect 36725 3451 36783 3457
rect 7432 3420 36676 3448
rect 7432 3408 7438 3420
rect 23566 3340 23572 3392
rect 23624 3340 23630 3392
rect 36354 3340 36360 3392
rect 36412 3340 36418 3392
rect 36648 3380 36676 3420
rect 36725 3417 36737 3451
rect 36771 3448 36783 3451
rect 37200 3448 37228 3488
rect 37274 3476 37280 3488
rect 37332 3476 37338 3528
rect 41046 3476 41052 3528
rect 41104 3476 41110 3528
rect 41138 3476 41144 3528
rect 41196 3476 41202 3528
rect 41386 3488 41644 3516
rect 40221 3451 40279 3457
rect 40221 3448 40233 3451
rect 36771 3420 37228 3448
rect 37292 3420 40233 3448
rect 36771 3417 36783 3420
rect 36725 3411 36783 3417
rect 37292 3380 37320 3420
rect 40221 3417 40233 3420
rect 40267 3448 40279 3451
rect 41386 3448 41414 3488
rect 40267 3420 41414 3448
rect 40267 3417 40279 3420
rect 40221 3411 40279 3417
rect 41506 3408 41512 3460
rect 41564 3408 41570 3460
rect 41616 3448 41644 3488
rect 41877 3451 41935 3457
rect 41877 3448 41889 3451
rect 41616 3420 41889 3448
rect 41877 3417 41889 3420
rect 41923 3417 41935 3451
rect 41877 3411 41935 3417
rect 36648 3352 37320 3380
rect 37366 3340 37372 3392
rect 37424 3380 37430 3392
rect 37461 3383 37519 3389
rect 37461 3380 37473 3383
rect 37424 3352 37473 3380
rect 37424 3340 37430 3352
rect 37461 3349 37473 3352
rect 37507 3349 37519 3383
rect 37461 3343 37519 3349
rect 37645 3383 37703 3389
rect 37645 3349 37657 3383
rect 37691 3380 37703 3383
rect 39482 3380 39488 3392
rect 37691 3352 39488 3380
rect 37691 3349 37703 3352
rect 37645 3343 37703 3349
rect 39482 3340 39488 3352
rect 39540 3340 39546 3392
rect 40773 3383 40831 3389
rect 40773 3349 40785 3383
rect 40819 3380 40831 3383
rect 41230 3380 41236 3392
rect 40819 3352 41236 3380
rect 40819 3349 40831 3352
rect 40773 3343 40831 3349
rect 41230 3340 41236 3352
rect 41288 3340 41294 3392
rect 41322 3340 41328 3392
rect 41380 3380 41386 3392
rect 41984 3380 42012 3556
rect 42518 3544 42524 3556
rect 42576 3544 42582 3596
rect 45462 3584 45468 3596
rect 44298 3570 45468 3584
rect 44284 3556 45468 3570
rect 43533 3519 43591 3525
rect 43533 3485 43545 3519
rect 43579 3516 43591 3519
rect 43898 3516 43904 3528
rect 43579 3488 43904 3516
rect 43579 3485 43591 3488
rect 43533 3479 43591 3485
rect 43898 3476 43904 3488
rect 43956 3476 43962 3528
rect 43990 3476 43996 3528
rect 44048 3476 44054 3528
rect 43346 3408 43352 3460
rect 43404 3448 43410 3460
rect 43625 3451 43683 3457
rect 43625 3448 43637 3451
rect 43404 3420 43637 3448
rect 43404 3408 43410 3420
rect 43625 3417 43637 3420
rect 43671 3417 43683 3451
rect 43625 3411 43683 3417
rect 43806 3408 43812 3460
rect 43864 3448 43870 3460
rect 44284 3448 44312 3556
rect 45462 3544 45468 3556
rect 45520 3544 45526 3596
rect 47762 3544 47768 3596
rect 47820 3584 47826 3596
rect 47946 3584 47952 3596
rect 47820 3556 47952 3584
rect 47820 3544 47826 3556
rect 47946 3544 47952 3556
rect 48004 3584 48010 3596
rect 51626 3584 51632 3596
rect 48004 3570 48070 3584
rect 48004 3556 48084 3570
rect 51566 3556 51632 3584
rect 48004 3544 48010 3556
rect 48056 3516 48084 3556
rect 51626 3544 51632 3556
rect 51684 3544 51690 3596
rect 80026 3584 80054 3692
rect 92474 3680 92480 3692
rect 92532 3680 92538 3732
rect 92566 3680 92572 3732
rect 92624 3680 92630 3732
rect 95789 3723 95847 3729
rect 94056 3692 95740 3720
rect 92017 3655 92075 3661
rect 92017 3621 92029 3655
rect 92063 3652 92075 3655
rect 92198 3652 92204 3664
rect 92063 3624 92204 3652
rect 92063 3621 92075 3624
rect 92017 3615 92075 3621
rect 92198 3612 92204 3624
rect 92256 3652 92262 3664
rect 94056 3652 94084 3692
rect 92256 3624 94084 3652
rect 92256 3612 92262 3624
rect 94130 3612 94136 3664
rect 94188 3652 94194 3664
rect 94593 3655 94651 3661
rect 94593 3652 94605 3655
rect 94188 3624 94605 3652
rect 94188 3612 94194 3624
rect 94593 3621 94605 3624
rect 94639 3652 94651 3655
rect 94682 3652 94688 3664
rect 94639 3624 94688 3652
rect 94639 3621 94651 3624
rect 94593 3615 94651 3621
rect 94682 3612 94688 3624
rect 94740 3612 94746 3664
rect 94498 3584 94504 3596
rect 68756 3556 80054 3584
rect 89686 3556 94504 3584
rect 48774 3516 48780 3528
rect 48056 3488 48780 3516
rect 48774 3476 48780 3488
rect 48832 3476 48838 3528
rect 48958 3476 48964 3528
rect 49016 3476 49022 3528
rect 50430 3476 50436 3528
rect 50488 3516 50494 3528
rect 50801 3519 50859 3525
rect 50801 3516 50813 3519
rect 50488 3488 50813 3516
rect 50488 3476 50494 3488
rect 50801 3485 50813 3488
rect 50847 3485 50859 3519
rect 50801 3479 50859 3485
rect 50890 3476 50896 3528
rect 50948 3476 50954 3528
rect 68756 3525 68784 3556
rect 68741 3519 68799 3525
rect 51046 3488 64874 3516
rect 43864 3420 44312 3448
rect 43864 3408 43870 3420
rect 48222 3408 48228 3460
rect 48280 3408 48286 3460
rect 48406 3408 48412 3460
rect 48464 3448 48470 3460
rect 48501 3451 48559 3457
rect 48501 3448 48513 3451
rect 48464 3420 48513 3448
rect 48464 3408 48470 3420
rect 48501 3417 48513 3420
rect 48547 3417 48559 3451
rect 48501 3411 48559 3417
rect 48590 3408 48596 3460
rect 48648 3408 48654 3460
rect 51046 3448 51074 3488
rect 49252 3420 51074 3448
rect 51261 3451 51319 3457
rect 41380 3352 42012 3380
rect 41380 3340 41386 3352
rect 42058 3340 42064 3392
rect 42116 3340 42122 3392
rect 43257 3383 43315 3389
rect 43257 3349 43269 3383
rect 43303 3380 43315 3383
rect 43438 3380 43444 3392
rect 43303 3352 43444 3380
rect 43303 3349 43315 3352
rect 43257 3343 43315 3349
rect 43438 3340 43444 3352
rect 43496 3340 43502 3392
rect 44358 3340 44364 3392
rect 44416 3340 44422 3392
rect 44545 3383 44603 3389
rect 44545 3349 44557 3383
rect 44591 3380 44603 3383
rect 49252 3380 49280 3420
rect 51261 3417 51273 3451
rect 51307 3448 51319 3451
rect 51534 3448 51540 3460
rect 51307 3420 51540 3448
rect 51307 3417 51319 3420
rect 51261 3411 51319 3417
rect 51534 3408 51540 3420
rect 51592 3408 51598 3460
rect 64846 3448 64874 3488
rect 68741 3485 68753 3519
rect 68787 3485 68799 3519
rect 89686 3516 89714 3556
rect 94498 3544 94504 3556
rect 94556 3544 94562 3596
rect 94866 3544 94872 3596
rect 94924 3544 94930 3596
rect 95050 3593 95056 3596
rect 95007 3587 95056 3593
rect 95007 3553 95019 3587
rect 95053 3553 95056 3587
rect 95007 3547 95056 3553
rect 95050 3544 95056 3547
rect 95108 3544 95114 3596
rect 95145 3587 95203 3593
rect 95145 3553 95157 3587
rect 95191 3584 95203 3587
rect 95510 3584 95516 3596
rect 95191 3556 95516 3584
rect 95191 3553 95203 3556
rect 95145 3547 95203 3553
rect 95510 3544 95516 3556
rect 95568 3544 95574 3596
rect 68741 3479 68799 3485
rect 74506 3488 89714 3516
rect 74506 3448 74534 3488
rect 91922 3476 91928 3528
rect 91980 3476 91986 3528
rect 92753 3519 92811 3525
rect 92753 3485 92765 3519
rect 92799 3485 92811 3519
rect 92753 3479 92811 3485
rect 92658 3448 92664 3460
rect 64846 3420 74534 3448
rect 80026 3420 92664 3448
rect 44591 3352 49280 3380
rect 44591 3349 44603 3352
rect 44545 3343 44603 3349
rect 49326 3340 49332 3392
rect 49384 3340 49390 3392
rect 49510 3340 49516 3392
rect 49568 3340 49574 3392
rect 50430 3340 50436 3392
rect 50488 3380 50494 3392
rect 50525 3383 50583 3389
rect 50525 3380 50537 3383
rect 50488 3352 50537 3380
rect 50488 3340 50494 3352
rect 50525 3349 50537 3352
rect 50571 3349 50583 3383
rect 50525 3343 50583 3349
rect 51626 3340 51632 3392
rect 51684 3340 51690 3392
rect 51810 3340 51816 3392
rect 51868 3340 51874 3392
rect 52086 3340 52092 3392
rect 52144 3380 52150 3392
rect 80026 3380 80054 3420
rect 92658 3408 92664 3420
rect 92716 3408 92722 3460
rect 92768 3448 92796 3479
rect 93210 3476 93216 3528
rect 93268 3476 93274 3528
rect 93946 3476 93952 3528
rect 94004 3476 94010 3528
rect 94038 3476 94044 3528
rect 94096 3516 94102 3528
rect 94133 3519 94191 3525
rect 94133 3516 94145 3519
rect 94096 3488 94145 3516
rect 94096 3476 94102 3488
rect 94133 3485 94145 3488
rect 94179 3485 94191 3519
rect 94133 3479 94191 3485
rect 95712 3448 95740 3692
rect 95789 3689 95801 3723
rect 95835 3720 95847 3723
rect 96890 3720 96896 3732
rect 95835 3692 96896 3720
rect 95835 3689 95847 3692
rect 95789 3683 95847 3689
rect 96890 3680 96896 3692
rect 96948 3680 96954 3732
rect 96982 3680 96988 3732
rect 97040 3680 97046 3732
rect 101766 3680 101772 3732
rect 101824 3720 101830 3732
rect 101861 3723 101919 3729
rect 101861 3720 101873 3723
rect 101824 3692 101873 3720
rect 101824 3680 101830 3692
rect 101861 3689 101873 3692
rect 101907 3689 101919 3723
rect 101861 3683 101919 3689
rect 101950 3680 101956 3732
rect 102008 3720 102014 3732
rect 102229 3723 102287 3729
rect 102229 3720 102241 3723
rect 102008 3692 102241 3720
rect 102008 3680 102014 3692
rect 102229 3689 102241 3692
rect 102275 3689 102287 3723
rect 102229 3683 102287 3689
rect 105354 3680 105360 3732
rect 105412 3680 105418 3732
rect 106182 3680 106188 3732
rect 106240 3680 106246 3732
rect 106366 3680 106372 3732
rect 106424 3720 106430 3732
rect 106461 3723 106519 3729
rect 106461 3720 106473 3723
rect 106424 3692 106473 3720
rect 106424 3680 106430 3692
rect 106461 3689 106473 3692
rect 106507 3689 106519 3723
rect 106461 3683 106519 3689
rect 108758 3680 108764 3732
rect 108816 3720 108822 3732
rect 108816 3692 111380 3720
rect 108816 3680 108822 3692
rect 95970 3612 95976 3664
rect 96028 3652 96034 3664
rect 97718 3652 97724 3664
rect 96028 3624 97724 3652
rect 96028 3612 96034 3624
rect 97718 3612 97724 3624
rect 97776 3612 97782 3664
rect 100754 3612 100760 3664
rect 100812 3652 100818 3664
rect 102781 3655 102839 3661
rect 102781 3652 102793 3655
rect 100812 3624 102793 3652
rect 100812 3612 100818 3624
rect 102781 3621 102793 3624
rect 102827 3621 102839 3655
rect 102781 3615 102839 3621
rect 104158 3612 104164 3664
rect 104216 3612 104222 3664
rect 105170 3612 105176 3664
rect 105228 3652 105234 3664
rect 105228 3624 106044 3652
rect 105228 3612 105234 3624
rect 99101 3587 99159 3593
rect 99101 3584 99113 3587
rect 96816 3556 99113 3584
rect 96816 3528 96844 3556
rect 99101 3553 99113 3556
rect 99147 3553 99159 3587
rect 99101 3547 99159 3553
rect 99282 3544 99288 3596
rect 99340 3544 99346 3596
rect 101398 3544 101404 3596
rect 101456 3584 101462 3596
rect 101953 3587 102011 3593
rect 101953 3584 101965 3587
rect 101456 3556 101965 3584
rect 101456 3544 101462 3556
rect 101953 3553 101965 3556
rect 101999 3553 102011 3587
rect 101953 3547 102011 3553
rect 103698 3544 103704 3596
rect 103756 3544 103762 3596
rect 104434 3544 104440 3596
rect 104492 3544 104498 3596
rect 104551 3544 104557 3596
rect 104609 3544 104615 3596
rect 104713 3587 104771 3593
rect 104713 3553 104725 3587
rect 104759 3584 104771 3587
rect 105630 3584 105636 3596
rect 104759 3556 105636 3584
rect 104759 3553 104771 3556
rect 104713 3547 104771 3553
rect 105630 3544 105636 3556
rect 105688 3544 105694 3596
rect 96798 3476 96804 3528
rect 96856 3476 96862 3528
rect 96890 3476 96896 3528
rect 96948 3516 96954 3528
rect 96985 3519 97043 3525
rect 96985 3516 96997 3519
rect 96948 3488 96997 3516
rect 96948 3476 96954 3488
rect 96985 3485 96997 3488
rect 97031 3485 97043 3519
rect 96985 3479 97043 3485
rect 97169 3519 97227 3525
rect 97169 3485 97181 3519
rect 97215 3516 97227 3519
rect 97350 3516 97356 3528
rect 97215 3488 97356 3516
rect 97215 3485 97227 3488
rect 97169 3479 97227 3485
rect 97350 3476 97356 3488
rect 97408 3476 97414 3528
rect 97813 3519 97871 3525
rect 97813 3485 97825 3519
rect 97859 3485 97871 3519
rect 97813 3479 97871 3485
rect 98089 3519 98147 3525
rect 98089 3485 98101 3519
rect 98135 3485 98147 3519
rect 98089 3479 98147 3485
rect 97828 3448 97856 3479
rect 92768 3420 94084 3448
rect 95712 3420 97856 3448
rect 98104 3448 98132 3479
rect 101858 3476 101864 3528
rect 101916 3476 101922 3528
rect 102226 3476 102232 3528
rect 102284 3516 102290 3528
rect 102597 3519 102655 3525
rect 102597 3516 102609 3519
rect 102284 3488 102609 3516
rect 102284 3476 102290 3488
rect 102597 3485 102609 3488
rect 102643 3485 102655 3519
rect 102597 3479 102655 3485
rect 103517 3519 103575 3525
rect 103517 3485 103529 3519
rect 103563 3485 103575 3519
rect 103517 3479 103575 3485
rect 99374 3448 99380 3460
rect 98104 3420 99380 3448
rect 52144 3352 80054 3380
rect 93397 3383 93455 3389
rect 52144 3340 52150 3352
rect 93397 3349 93409 3383
rect 93443 3380 93455 3383
rect 93946 3380 93952 3392
rect 93443 3352 93952 3380
rect 93443 3349 93455 3352
rect 93397 3343 93455 3349
rect 93946 3340 93952 3352
rect 94004 3340 94010 3392
rect 94056 3380 94084 3420
rect 99374 3408 99380 3420
rect 99432 3408 99438 3460
rect 100938 3408 100944 3460
rect 100996 3408 101002 3460
rect 103146 3408 103152 3460
rect 103204 3448 103210 3460
rect 103532 3448 103560 3479
rect 105538 3476 105544 3528
rect 105596 3516 105602 3528
rect 105909 3519 105967 3525
rect 105909 3516 105921 3519
rect 105596 3488 105921 3516
rect 105596 3476 105602 3488
rect 105909 3485 105921 3488
rect 105955 3485 105967 3519
rect 106016 3516 106044 3624
rect 106550 3612 106556 3664
rect 106608 3652 106614 3664
rect 111352 3652 111380 3692
rect 111610 3680 111616 3732
rect 111668 3680 111674 3732
rect 111702 3680 111708 3732
rect 111760 3720 111766 3732
rect 119617 3723 119675 3729
rect 111760 3692 119568 3720
rect 111760 3680 111766 3692
rect 117406 3652 117412 3664
rect 106608 3624 108896 3652
rect 111352 3624 117412 3652
rect 106608 3612 106614 3624
rect 108868 3596 108896 3624
rect 117406 3612 117412 3624
rect 117464 3612 117470 3664
rect 118142 3612 118148 3664
rect 118200 3652 118206 3664
rect 118418 3652 118424 3664
rect 118200 3624 118424 3652
rect 118200 3612 118206 3624
rect 118418 3612 118424 3624
rect 118476 3612 118482 3664
rect 119540 3652 119568 3692
rect 119617 3689 119629 3723
rect 119663 3720 119675 3723
rect 121454 3720 121460 3732
rect 119663 3692 121460 3720
rect 119663 3689 119675 3692
rect 119617 3683 119675 3689
rect 121454 3680 121460 3692
rect 121512 3680 121518 3732
rect 122466 3680 122472 3732
rect 122524 3680 122530 3732
rect 138937 3723 138995 3729
rect 138937 3689 138949 3723
rect 138983 3720 138995 3723
rect 140682 3720 140688 3732
rect 138983 3692 140688 3720
rect 138983 3689 138995 3692
rect 138937 3683 138995 3689
rect 140682 3680 140688 3692
rect 140740 3680 140746 3732
rect 141973 3723 142031 3729
rect 141973 3689 141985 3723
rect 142019 3720 142031 3723
rect 142246 3720 142252 3732
rect 142019 3692 142252 3720
rect 142019 3689 142031 3692
rect 141973 3683 142031 3689
rect 120902 3652 120908 3664
rect 119540 3624 120908 3652
rect 120902 3612 120908 3624
rect 120960 3612 120966 3664
rect 128326 3624 138014 3652
rect 106090 3544 106096 3596
rect 106148 3584 106154 3596
rect 107197 3587 107255 3593
rect 107197 3584 107209 3587
rect 106148 3556 107209 3584
rect 106148 3544 106154 3556
rect 107197 3553 107209 3556
rect 107243 3553 107255 3587
rect 107197 3547 107255 3553
rect 108850 3544 108856 3596
rect 108908 3544 108914 3596
rect 109402 3544 109408 3596
rect 109460 3584 109466 3596
rect 109773 3587 109831 3593
rect 109773 3584 109785 3587
rect 109460 3556 109785 3584
rect 109460 3544 109466 3556
rect 109773 3553 109785 3556
rect 109819 3553 109831 3587
rect 109773 3547 109831 3553
rect 110414 3544 110420 3596
rect 110472 3544 110478 3596
rect 110690 3544 110696 3596
rect 110748 3544 110754 3596
rect 110969 3587 111027 3593
rect 110969 3553 110981 3587
rect 111015 3584 111027 3587
rect 111518 3584 111524 3596
rect 111015 3556 111524 3584
rect 111015 3553 111027 3556
rect 110969 3547 111027 3553
rect 111518 3544 111524 3556
rect 111576 3584 111582 3596
rect 111794 3584 111800 3596
rect 111576 3556 111800 3584
rect 111576 3544 111582 3556
rect 111794 3544 111800 3556
rect 111852 3544 111858 3596
rect 112165 3587 112223 3593
rect 112165 3553 112177 3587
rect 112211 3584 112223 3587
rect 112530 3584 112536 3596
rect 112211 3556 112536 3584
rect 112211 3553 112223 3556
rect 112165 3547 112223 3553
rect 112530 3544 112536 3556
rect 112588 3544 112594 3596
rect 113726 3544 113732 3596
rect 113784 3544 113790 3596
rect 114830 3544 114836 3596
rect 114888 3584 114894 3596
rect 115109 3587 115167 3593
rect 115109 3584 115121 3587
rect 114888 3556 115121 3584
rect 114888 3544 114894 3556
rect 115109 3553 115121 3556
rect 115155 3553 115167 3587
rect 115109 3547 115167 3553
rect 117682 3544 117688 3596
rect 117740 3584 117746 3596
rect 118510 3584 118516 3596
rect 117740 3556 118516 3584
rect 117740 3544 117746 3556
rect 118510 3544 118516 3556
rect 118568 3544 118574 3596
rect 118697 3587 118755 3593
rect 118697 3553 118709 3587
rect 118743 3584 118755 3587
rect 119154 3584 119160 3596
rect 118743 3556 119160 3584
rect 118743 3553 118755 3556
rect 118697 3547 118755 3553
rect 119154 3544 119160 3556
rect 119212 3544 119218 3596
rect 120074 3544 120080 3596
rect 120132 3544 120138 3596
rect 120261 3587 120319 3593
rect 120261 3553 120273 3587
rect 120307 3584 120319 3587
rect 122282 3584 122288 3596
rect 120307 3556 122288 3584
rect 120307 3553 120319 3556
rect 120261 3547 120319 3553
rect 122282 3544 122288 3556
rect 122340 3544 122346 3596
rect 106182 3516 106188 3528
rect 106016 3488 106188 3516
rect 105909 3479 105967 3485
rect 106182 3476 106188 3488
rect 106240 3476 106246 3528
rect 106274 3476 106280 3528
rect 106332 3516 106338 3528
rect 110874 3525 110880 3528
rect 107013 3519 107071 3525
rect 107013 3516 107025 3519
rect 106332 3488 107025 3516
rect 106332 3476 106338 3488
rect 107013 3485 107025 3488
rect 107059 3485 107071 3519
rect 107013 3479 107071 3485
rect 109957 3519 110015 3525
rect 109957 3485 109969 3519
rect 110003 3485 110015 3519
rect 109957 3479 110015 3485
rect 110831 3519 110880 3525
rect 110831 3485 110843 3519
rect 110877 3485 110880 3519
rect 110831 3479 110880 3485
rect 103204 3420 103560 3448
rect 103204 3408 103210 3420
rect 105722 3408 105728 3460
rect 105780 3448 105786 3460
rect 109972 3448 110000 3479
rect 110874 3476 110880 3479
rect 110932 3476 110938 3528
rect 114922 3476 114928 3528
rect 114980 3476 114986 3528
rect 117314 3476 117320 3528
rect 117372 3516 117378 3528
rect 117777 3519 117835 3525
rect 117777 3516 117789 3519
rect 117372 3488 117789 3516
rect 117372 3476 117378 3488
rect 117777 3485 117789 3488
rect 117823 3485 117835 3519
rect 117777 3479 117835 3485
rect 117866 3476 117872 3528
rect 117924 3516 117930 3528
rect 118878 3525 118884 3528
rect 117961 3519 118019 3525
rect 117961 3516 117973 3519
rect 117924 3488 117973 3516
rect 117924 3476 117930 3488
rect 117961 3485 117973 3488
rect 118007 3485 118019 3519
rect 117961 3479 118019 3485
rect 118835 3519 118884 3525
rect 118835 3485 118847 3519
rect 118881 3485 118884 3519
rect 118835 3479 118884 3485
rect 118878 3476 118884 3479
rect 118936 3476 118942 3528
rect 118970 3476 118976 3528
rect 119028 3476 119034 3528
rect 121917 3519 121975 3525
rect 121917 3485 121929 3519
rect 121963 3516 121975 3519
rect 122098 3516 122104 3528
rect 121963 3488 122104 3516
rect 121963 3485 121975 3488
rect 121917 3479 121975 3485
rect 122098 3476 122104 3488
rect 122156 3476 122162 3528
rect 122653 3519 122711 3525
rect 122653 3485 122665 3519
rect 122699 3516 122711 3519
rect 123018 3516 123024 3528
rect 122699 3488 123024 3516
rect 122699 3485 122711 3488
rect 122653 3479 122711 3485
rect 123018 3476 123024 3488
rect 123076 3476 123082 3528
rect 105780 3420 110000 3448
rect 105780 3408 105786 3420
rect 112162 3408 112168 3460
rect 112220 3448 112226 3460
rect 112349 3451 112407 3457
rect 112349 3448 112361 3451
rect 112220 3420 112361 3448
rect 112220 3408 112226 3420
rect 112349 3417 112361 3420
rect 112395 3417 112407 3451
rect 112349 3411 112407 3417
rect 116765 3451 116823 3457
rect 116765 3417 116777 3451
rect 116811 3417 116823 3451
rect 116765 3411 116823 3417
rect 97353 3383 97411 3389
rect 97353 3380 97365 3383
rect 94056 3352 97365 3380
rect 97353 3349 97365 3352
rect 97399 3349 97411 3383
rect 97353 3343 97411 3349
rect 98454 3340 98460 3392
rect 98512 3380 98518 3392
rect 103054 3380 103060 3392
rect 98512 3352 103060 3380
rect 98512 3340 98518 3352
rect 103054 3340 103060 3352
rect 103112 3340 103118 3392
rect 103698 3340 103704 3392
rect 103756 3380 103762 3392
rect 107654 3380 107660 3392
rect 103756 3352 107660 3380
rect 103756 3340 103762 3352
rect 107654 3340 107660 3352
rect 107712 3340 107718 3392
rect 110414 3340 110420 3392
rect 110472 3380 110478 3392
rect 111242 3380 111248 3392
rect 110472 3352 111248 3380
rect 110472 3340 110478 3352
rect 111242 3340 111248 3352
rect 111300 3340 111306 3392
rect 116780 3380 116808 3411
rect 119246 3380 119252 3392
rect 116780 3352 119252 3380
rect 119246 3340 119252 3352
rect 119304 3380 119310 3392
rect 128326 3380 128354 3624
rect 137986 3584 138014 3624
rect 139486 3612 139492 3664
rect 139544 3652 139550 3664
rect 141988 3652 142016 3683
rect 142246 3680 142252 3692
rect 142304 3680 142310 3732
rect 145834 3680 145840 3732
rect 145892 3720 145898 3732
rect 148229 3723 148287 3729
rect 148229 3720 148241 3723
rect 145892 3692 148241 3720
rect 145892 3680 145898 3692
rect 148229 3689 148241 3692
rect 148275 3689 148287 3723
rect 148229 3683 148287 3689
rect 149238 3680 149244 3732
rect 149296 3680 149302 3732
rect 151446 3720 151452 3732
rect 150728 3692 151452 3720
rect 139544 3624 142016 3652
rect 139544 3612 139550 3624
rect 144730 3612 144736 3664
rect 144788 3652 144794 3664
rect 145926 3652 145932 3664
rect 144788 3624 145932 3652
rect 144788 3612 144794 3624
rect 145926 3612 145932 3624
rect 145984 3612 145990 3664
rect 146680 3624 147628 3652
rect 146680 3584 146708 3624
rect 137986 3556 146708 3584
rect 147600 3600 147628 3624
rect 148502 3612 148508 3664
rect 148560 3652 148566 3664
rect 150728 3652 150756 3692
rect 151446 3680 151452 3692
rect 151504 3720 151510 3732
rect 151504 3692 154068 3720
rect 151504 3680 151510 3692
rect 148560 3624 150756 3652
rect 148560 3612 148566 3624
rect 150802 3612 150808 3664
rect 150860 3652 150866 3664
rect 152553 3655 152611 3661
rect 152553 3652 152565 3655
rect 150860 3624 152565 3652
rect 150860 3612 150866 3624
rect 152553 3621 152565 3624
rect 152599 3621 152611 3655
rect 152553 3615 152611 3621
rect 152826 3612 152832 3664
rect 152884 3652 152890 3664
rect 153654 3652 153660 3664
rect 152884 3624 153660 3652
rect 152884 3612 152890 3624
rect 153654 3612 153660 3624
rect 153712 3612 153718 3664
rect 154040 3661 154068 3692
rect 154298 3680 154304 3732
rect 154356 3720 154362 3732
rect 154356 3692 154988 3720
rect 154356 3680 154362 3692
rect 154025 3655 154083 3661
rect 154025 3621 154037 3655
rect 154071 3621 154083 3655
rect 154960 3652 154988 3692
rect 155218 3680 155224 3732
rect 155276 3680 155282 3732
rect 155328 3692 158760 3720
rect 155328 3652 155356 3692
rect 154960 3624 155356 3652
rect 154025 3615 154083 3621
rect 156322 3612 156328 3664
rect 156380 3612 156386 3664
rect 157260 3624 158668 3652
rect 147600 3584 147674 3600
rect 149514 3584 149520 3596
rect 147600 3572 149520 3584
rect 147646 3556 149520 3572
rect 149514 3544 149520 3556
rect 149572 3544 149578 3596
rect 150253 3587 150311 3593
rect 150253 3553 150265 3587
rect 150299 3584 150311 3587
rect 152642 3584 152648 3596
rect 150299 3556 152648 3584
rect 150299 3553 150311 3556
rect 150253 3547 150311 3553
rect 152642 3544 152648 3556
rect 152700 3544 152706 3596
rect 153378 3544 153384 3596
rect 153436 3544 153442 3596
rect 153565 3587 153623 3593
rect 153565 3553 153577 3587
rect 153611 3584 153623 3587
rect 153930 3584 153936 3596
rect 153611 3556 153936 3584
rect 153611 3553 153623 3556
rect 153565 3547 153623 3553
rect 153930 3544 153936 3556
rect 153988 3544 153994 3596
rect 154301 3587 154359 3593
rect 154301 3553 154313 3587
rect 154347 3584 154359 3587
rect 154942 3584 154948 3596
rect 154347 3556 154948 3584
rect 154347 3553 154359 3556
rect 154301 3547 154359 3553
rect 154942 3544 154948 3556
rect 155000 3544 155006 3596
rect 155218 3544 155224 3596
rect 155276 3584 155282 3596
rect 155865 3587 155923 3593
rect 155865 3584 155877 3587
rect 155276 3556 155877 3584
rect 155276 3544 155282 3556
rect 155865 3553 155877 3556
rect 155911 3553 155923 3587
rect 155865 3547 155923 3553
rect 156598 3544 156604 3596
rect 156656 3544 156662 3596
rect 156739 3587 156797 3593
rect 156739 3553 156751 3587
rect 156785 3584 156797 3587
rect 157260 3584 157288 3624
rect 156785 3556 157288 3584
rect 156785 3553 156797 3556
rect 156739 3547 156797 3553
rect 138477 3519 138535 3525
rect 138477 3485 138489 3519
rect 138523 3516 138535 3519
rect 138934 3516 138940 3528
rect 138523 3488 138940 3516
rect 138523 3485 138535 3488
rect 138477 3479 138535 3485
rect 138934 3476 138940 3488
rect 138992 3476 138998 3528
rect 139118 3476 139124 3528
rect 139176 3476 139182 3528
rect 139578 3476 139584 3528
rect 139636 3476 139642 3528
rect 141421 3519 141479 3525
rect 141421 3485 141433 3519
rect 141467 3516 141479 3519
rect 141510 3516 141516 3528
rect 141467 3488 141516 3516
rect 141467 3485 141479 3488
rect 141421 3479 141479 3485
rect 141510 3476 141516 3488
rect 141568 3476 141574 3528
rect 141602 3476 141608 3528
rect 141660 3516 141666 3528
rect 141878 3516 141884 3528
rect 141660 3488 141884 3516
rect 141660 3476 141666 3488
rect 141878 3476 141884 3488
rect 141936 3476 141942 3528
rect 142249 3519 142307 3525
rect 142249 3485 142261 3519
rect 142295 3485 142307 3519
rect 142249 3479 142307 3485
rect 139486 3408 139492 3460
rect 139544 3448 139550 3460
rect 139765 3451 139823 3457
rect 139765 3448 139777 3451
rect 139544 3420 139777 3448
rect 139544 3408 139550 3420
rect 139765 3417 139777 3420
rect 139811 3417 139823 3451
rect 139765 3411 139823 3417
rect 141970 3408 141976 3460
rect 142028 3448 142034 3460
rect 142264 3448 142292 3479
rect 142338 3476 142344 3528
rect 142396 3516 142402 3528
rect 143077 3519 143135 3525
rect 143077 3516 143089 3519
rect 142396 3488 143089 3516
rect 142396 3476 142402 3488
rect 143077 3485 143089 3488
rect 143123 3485 143135 3519
rect 143077 3479 143135 3485
rect 145377 3519 145435 3525
rect 145377 3485 145389 3519
rect 145423 3485 145435 3519
rect 148413 3519 148471 3525
rect 148413 3516 148425 3519
rect 145377 3479 145435 3485
rect 146772 3488 148425 3516
rect 142522 3448 142528 3460
rect 142028 3420 142528 3448
rect 142028 3408 142034 3420
rect 142522 3408 142528 3420
rect 142580 3408 142586 3460
rect 143258 3408 143264 3460
rect 143316 3408 143322 3460
rect 143626 3408 143632 3460
rect 143684 3448 143690 3460
rect 144822 3448 144828 3460
rect 143684 3420 144828 3448
rect 143684 3408 143690 3420
rect 144822 3408 144828 3420
rect 144880 3448 144886 3460
rect 144917 3451 144975 3457
rect 144917 3448 144929 3451
rect 144880 3420 144929 3448
rect 144880 3408 144886 3420
rect 144917 3417 144929 3420
rect 144963 3417 144975 3451
rect 144917 3411 144975 3417
rect 119304 3352 128354 3380
rect 119304 3340 119310 3352
rect 138290 3340 138296 3392
rect 138348 3340 138354 3392
rect 139026 3340 139032 3392
rect 139084 3380 139090 3392
rect 142433 3383 142491 3389
rect 142433 3380 142445 3383
rect 139084 3352 142445 3380
rect 139084 3340 139090 3352
rect 142433 3349 142445 3352
rect 142479 3349 142491 3383
rect 145392 3380 145420 3479
rect 145558 3408 145564 3460
rect 145616 3408 145622 3460
rect 145926 3408 145932 3460
rect 145984 3448 145990 3460
rect 146772 3448 146800 3488
rect 148413 3485 148425 3488
rect 148459 3485 148471 3519
rect 148413 3479 148471 3485
rect 149146 3476 149152 3528
rect 149204 3476 149210 3528
rect 149422 3476 149428 3528
rect 149480 3476 149486 3528
rect 152734 3476 152740 3528
rect 152792 3476 152798 3528
rect 153286 3476 153292 3528
rect 153344 3476 153350 3528
rect 154482 3525 154488 3528
rect 154439 3519 154488 3525
rect 154439 3485 154451 3519
rect 154485 3485 154488 3519
rect 154439 3479 154488 3485
rect 154482 3476 154488 3479
rect 154540 3476 154546 3528
rect 154574 3476 154580 3528
rect 154632 3476 154638 3528
rect 155586 3476 155592 3528
rect 155644 3516 155650 3528
rect 155681 3519 155739 3525
rect 155681 3516 155693 3519
rect 155644 3488 155693 3516
rect 155644 3476 155650 3488
rect 155681 3485 155693 3488
rect 155727 3485 155739 3519
rect 155681 3479 155739 3485
rect 156874 3476 156880 3528
rect 156932 3476 156938 3528
rect 145984 3420 146800 3448
rect 145984 3408 145990 3420
rect 147214 3408 147220 3460
rect 147272 3408 147278 3460
rect 149238 3408 149244 3460
rect 149296 3448 149302 3460
rect 149606 3448 149612 3460
rect 149296 3420 149612 3448
rect 149296 3408 149302 3420
rect 149606 3408 149612 3420
rect 149664 3408 149670 3460
rect 150434 3408 150440 3460
rect 150492 3408 150498 3460
rect 151722 3408 151728 3460
rect 151780 3448 151786 3460
rect 152093 3451 152151 3457
rect 152093 3448 152105 3451
rect 151780 3420 152105 3448
rect 151780 3408 151786 3420
rect 152093 3417 152105 3420
rect 152139 3448 152151 3451
rect 153304 3448 153332 3476
rect 152139 3420 153332 3448
rect 158640 3448 158668 3624
rect 158732 3525 158760 3692
rect 160094 3680 160100 3732
rect 160152 3720 160158 3732
rect 172698 3720 172704 3732
rect 160152 3692 172704 3720
rect 160152 3680 160158 3692
rect 172698 3680 172704 3692
rect 172756 3680 172762 3732
rect 207474 3680 207480 3732
rect 207532 3720 207538 3732
rect 208857 3723 208915 3729
rect 208857 3720 208869 3723
rect 207532 3692 208869 3720
rect 207532 3680 207538 3692
rect 208857 3689 208869 3692
rect 208903 3689 208915 3723
rect 208857 3683 208915 3689
rect 211338 3680 211344 3732
rect 211396 3720 211402 3732
rect 211396 3692 212655 3720
rect 211396 3680 211402 3692
rect 159634 3612 159640 3664
rect 159692 3652 159698 3664
rect 182082 3652 182088 3664
rect 159692 3624 182088 3652
rect 159692 3612 159698 3624
rect 182082 3612 182088 3624
rect 182140 3612 182146 3664
rect 208670 3612 208676 3664
rect 208728 3652 208734 3664
rect 208728 3624 210280 3652
rect 208728 3612 208734 3624
rect 168374 3584 168380 3596
rect 159468 3556 168380 3584
rect 158717 3519 158775 3525
rect 158717 3485 158729 3519
rect 158763 3485 158775 3519
rect 158717 3479 158775 3485
rect 159358 3476 159364 3528
rect 159416 3476 159422 3528
rect 159468 3448 159496 3556
rect 168374 3544 168380 3556
rect 168432 3544 168438 3596
rect 171778 3544 171784 3596
rect 171836 3584 171842 3596
rect 189718 3584 189724 3596
rect 171836 3556 189724 3584
rect 171836 3544 171842 3556
rect 189718 3544 189724 3556
rect 189776 3544 189782 3596
rect 207014 3544 207020 3596
rect 207072 3544 207078 3596
rect 207201 3587 207259 3593
rect 207201 3553 207213 3587
rect 207247 3584 207259 3587
rect 207566 3584 207572 3596
rect 207247 3556 207572 3584
rect 207247 3553 207259 3556
rect 207201 3547 207259 3553
rect 207566 3544 207572 3556
rect 207624 3544 207630 3596
rect 207658 3544 207664 3596
rect 207716 3544 207722 3596
rect 208075 3587 208133 3593
rect 208075 3553 208087 3587
rect 208121 3584 208133 3587
rect 209866 3584 209872 3596
rect 208121 3556 209872 3584
rect 208121 3553 208133 3556
rect 208075 3547 208133 3553
rect 209866 3544 209872 3556
rect 209924 3544 209930 3596
rect 210252 3584 210280 3624
rect 212074 3612 212080 3664
rect 212132 3612 212138 3664
rect 210252 3556 211384 3584
rect 167641 3519 167699 3525
rect 167641 3485 167653 3519
rect 167687 3516 167699 3519
rect 168282 3516 168288 3528
rect 167687 3488 168288 3516
rect 167687 3485 167699 3488
rect 167641 3479 167699 3485
rect 168282 3476 168288 3488
rect 168340 3476 168346 3528
rect 207934 3476 207940 3528
rect 207992 3476 207998 3528
rect 208210 3476 208216 3528
rect 208268 3476 208274 3528
rect 210252 3525 210280 3556
rect 211356 3528 211384 3556
rect 211540 3556 211844 3584
rect 211540 3528 211568 3556
rect 210237 3519 210295 3525
rect 210237 3485 210249 3519
rect 210283 3485 210295 3519
rect 210237 3479 210295 3485
rect 210326 3476 210332 3528
rect 210384 3476 210390 3528
rect 210510 3476 210516 3528
rect 210568 3516 210574 3528
rect 210970 3516 210976 3528
rect 210568 3488 210976 3516
rect 210568 3476 210574 3488
rect 210970 3476 210976 3488
rect 211028 3476 211034 3528
rect 211338 3476 211344 3528
rect 211396 3516 211402 3528
rect 211433 3519 211491 3525
rect 211433 3516 211445 3519
rect 211396 3488 211445 3516
rect 211396 3476 211402 3488
rect 211433 3485 211445 3488
rect 211479 3485 211491 3519
rect 211433 3479 211491 3485
rect 211522 3476 211528 3528
rect 211580 3476 211586 3528
rect 211706 3476 211712 3528
rect 211764 3476 211770 3528
rect 211816 3516 211844 3556
rect 212627 3526 212655 3692
rect 212994 3680 213000 3732
rect 213052 3720 213058 3732
rect 214377 3723 214435 3729
rect 214377 3720 214389 3723
rect 213052 3692 214389 3720
rect 213052 3680 213058 3692
rect 214377 3689 214389 3692
rect 214423 3689 214435 3723
rect 214377 3683 214435 3689
rect 218698 3680 218704 3732
rect 218756 3720 218762 3732
rect 224678 3720 224684 3732
rect 218756 3692 224684 3720
rect 218756 3680 218762 3692
rect 224678 3680 224684 3692
rect 224736 3680 224742 3732
rect 224788 3692 228128 3720
rect 214190 3612 214196 3664
rect 214248 3652 214254 3664
rect 215386 3652 215392 3664
rect 214248 3624 215392 3652
rect 214248 3612 214254 3624
rect 215386 3612 215392 3624
rect 215444 3612 215450 3664
rect 216030 3612 216036 3664
rect 216088 3652 216094 3664
rect 217962 3652 217968 3664
rect 216088 3624 217968 3652
rect 216088 3612 216094 3624
rect 216625 3584 216653 3624
rect 217962 3612 217968 3624
rect 218020 3612 218026 3664
rect 218514 3612 218520 3664
rect 218572 3652 218578 3664
rect 219526 3652 219532 3664
rect 218572 3624 219532 3652
rect 218572 3612 218578 3624
rect 219526 3612 219532 3624
rect 219584 3612 219590 3664
rect 219894 3612 219900 3664
rect 219952 3652 219958 3664
rect 220357 3655 220415 3661
rect 220357 3652 220369 3655
rect 219952 3624 220369 3652
rect 219952 3612 219958 3624
rect 220357 3621 220369 3624
rect 220403 3621 220415 3655
rect 220357 3615 220415 3621
rect 221182 3612 221188 3664
rect 221240 3652 221246 3664
rect 224788 3652 224816 3692
rect 221240 3624 224816 3652
rect 221240 3612 221246 3624
rect 227346 3612 227352 3664
rect 227404 3612 227410 3664
rect 227622 3612 227628 3664
rect 227680 3652 227686 3664
rect 228100 3652 228128 3692
rect 228174 3680 228180 3732
rect 228232 3720 228238 3732
rect 243630 3720 243636 3732
rect 228232 3692 243636 3720
rect 228232 3680 228238 3692
rect 243630 3680 243636 3692
rect 243688 3680 243694 3732
rect 244461 3723 244519 3729
rect 244461 3689 244473 3723
rect 244507 3720 244519 3723
rect 245381 3723 245439 3729
rect 245381 3720 245393 3723
rect 244507 3692 245393 3720
rect 244507 3689 244519 3692
rect 244461 3683 244519 3689
rect 245381 3689 245393 3692
rect 245427 3720 245439 3723
rect 245654 3720 245660 3732
rect 245427 3692 245660 3720
rect 245427 3689 245439 3692
rect 245381 3683 245439 3689
rect 245654 3680 245660 3692
rect 245712 3720 245718 3732
rect 246482 3720 246488 3732
rect 245712 3692 246488 3720
rect 245712 3680 245718 3692
rect 246482 3680 246488 3692
rect 246540 3680 246546 3732
rect 246666 3680 246672 3732
rect 246724 3680 246730 3732
rect 247586 3680 247592 3732
rect 247644 3720 247650 3732
rect 251634 3720 251640 3732
rect 247644 3692 251640 3720
rect 247644 3680 247650 3692
rect 251634 3680 251640 3692
rect 251692 3680 251698 3732
rect 252554 3680 252560 3732
rect 252612 3680 252618 3732
rect 252830 3680 252836 3732
rect 252888 3720 252894 3732
rect 254118 3720 254124 3732
rect 252888 3692 254124 3720
rect 252888 3680 252894 3692
rect 254118 3680 254124 3692
rect 254176 3680 254182 3732
rect 257338 3680 257344 3732
rect 257396 3720 257402 3732
rect 258626 3720 258632 3732
rect 257396 3692 258632 3720
rect 257396 3680 257402 3692
rect 258626 3680 258632 3692
rect 258684 3720 258690 3732
rect 258721 3723 258779 3729
rect 258721 3720 258733 3723
rect 258684 3692 258733 3720
rect 258684 3680 258690 3692
rect 258721 3689 258733 3692
rect 258767 3689 258779 3723
rect 258721 3683 258779 3689
rect 258994 3680 259000 3732
rect 259052 3720 259058 3732
rect 260561 3723 260619 3729
rect 260561 3720 260573 3723
rect 259052 3692 260573 3720
rect 259052 3680 259058 3692
rect 260561 3689 260573 3692
rect 260607 3689 260619 3723
rect 260561 3683 260619 3689
rect 264790 3680 264796 3732
rect 264848 3720 264854 3732
rect 267734 3720 267740 3732
rect 264848 3692 267740 3720
rect 264848 3680 264854 3692
rect 267734 3680 267740 3692
rect 267792 3680 267798 3732
rect 267921 3723 267979 3729
rect 267921 3689 267933 3723
rect 267967 3720 267979 3723
rect 268194 3720 268200 3732
rect 267967 3692 268200 3720
rect 267967 3689 267979 3692
rect 267921 3683 267979 3689
rect 268194 3680 268200 3692
rect 268252 3680 268258 3732
rect 268838 3680 268844 3732
rect 268896 3680 268902 3732
rect 269114 3680 269120 3732
rect 269172 3720 269178 3732
rect 269209 3723 269267 3729
rect 269209 3720 269221 3723
rect 269172 3692 269221 3720
rect 269172 3680 269178 3692
rect 269209 3689 269221 3692
rect 269255 3689 269267 3723
rect 269209 3683 269267 3689
rect 270037 3723 270095 3729
rect 270037 3689 270049 3723
rect 270083 3720 270095 3723
rect 270678 3720 270684 3732
rect 270083 3692 270684 3720
rect 270083 3689 270095 3692
rect 270037 3683 270095 3689
rect 270678 3680 270684 3692
rect 270736 3680 270742 3732
rect 229738 3652 229744 3664
rect 227680 3624 227760 3652
rect 228100 3624 229744 3652
rect 227680 3612 227686 3624
rect 216600 3556 216653 3584
rect 212627 3525 212672 3526
rect 212627 3519 212687 3525
rect 211816 3488 212580 3516
rect 212627 3498 212641 3519
rect 158640 3420 159496 3448
rect 152139 3417 152151 3420
rect 152093 3411 152151 3417
rect 161198 3408 161204 3460
rect 161256 3448 161262 3460
rect 187142 3448 187148 3460
rect 161256 3420 187148 3448
rect 161256 3408 161262 3420
rect 187142 3408 187148 3420
rect 187200 3408 187206 3460
rect 209222 3408 209228 3460
rect 209280 3448 209286 3460
rect 210142 3448 210148 3460
rect 209280 3420 210148 3448
rect 209280 3408 209286 3420
rect 210142 3408 210148 3420
rect 210200 3408 210206 3460
rect 146294 3380 146300 3392
rect 145392 3352 146300 3380
rect 142433 3343 142491 3349
rect 146294 3340 146300 3352
rect 146352 3340 146358 3392
rect 149701 3383 149759 3389
rect 149701 3349 149713 3383
rect 149747 3380 149759 3383
rect 152458 3380 152464 3392
rect 149747 3352 152464 3380
rect 149747 3349 149759 3352
rect 149701 3343 149759 3349
rect 152458 3340 152464 3352
rect 152516 3340 152522 3392
rect 153286 3340 153292 3392
rect 153344 3380 153350 3392
rect 155862 3380 155868 3392
rect 153344 3352 155868 3380
rect 153344 3340 153350 3352
rect 155862 3340 155868 3352
rect 155920 3340 155926 3392
rect 156138 3340 156144 3392
rect 156196 3380 156202 3392
rect 157521 3383 157579 3389
rect 157521 3380 157533 3383
rect 156196 3352 157533 3380
rect 156196 3340 156202 3352
rect 157521 3349 157533 3352
rect 157567 3349 157579 3383
rect 157521 3343 157579 3349
rect 158530 3340 158536 3392
rect 158588 3340 158594 3392
rect 158622 3340 158628 3392
rect 158680 3380 158686 3392
rect 159177 3383 159235 3389
rect 159177 3380 159189 3383
rect 158680 3352 159189 3380
rect 158680 3340 158686 3352
rect 159177 3349 159189 3352
rect 159223 3349 159235 3383
rect 159177 3343 159235 3349
rect 167730 3340 167736 3392
rect 167788 3340 167794 3392
rect 206738 3340 206744 3392
rect 206796 3380 206802 3392
rect 207934 3380 207940 3392
rect 206796 3352 207940 3380
rect 206796 3340 206802 3352
rect 207934 3340 207940 3352
rect 207992 3380 207998 3392
rect 209038 3380 209044 3392
rect 207992 3352 209044 3380
rect 207992 3340 207998 3352
rect 209038 3340 209044 3352
rect 209096 3340 209102 3392
rect 210344 3380 210372 3476
rect 210881 3451 210939 3457
rect 210881 3417 210893 3451
rect 210927 3448 210939 3451
rect 212350 3448 212356 3460
rect 210927 3420 212356 3448
rect 210927 3417 210939 3420
rect 210881 3411 210939 3417
rect 212350 3408 212356 3420
rect 212408 3408 212414 3460
rect 212552 3448 212580 3488
rect 212629 3485 212641 3498
rect 212675 3485 212687 3519
rect 212629 3479 212687 3485
rect 212721 3519 212779 3525
rect 212721 3485 212733 3519
rect 212767 3485 212779 3519
rect 212721 3479 212779 3485
rect 212736 3448 212764 3479
rect 212994 3476 213000 3528
rect 213052 3476 213058 3528
rect 213917 3519 213975 3525
rect 213917 3516 213929 3519
rect 213196 3488 213929 3516
rect 213196 3448 213224 3488
rect 213917 3485 213929 3488
rect 213963 3485 213975 3519
rect 213917 3479 213975 3485
rect 214006 3476 214012 3528
rect 214064 3516 214070 3528
rect 214561 3519 214619 3525
rect 214561 3516 214573 3519
rect 214064 3488 214573 3516
rect 214064 3476 214070 3488
rect 214561 3485 214573 3488
rect 214607 3485 214619 3519
rect 214561 3479 214619 3485
rect 215570 3476 215576 3528
rect 215628 3476 215634 3528
rect 215757 3519 215815 3525
rect 215757 3485 215769 3519
rect 215803 3516 215815 3519
rect 216490 3516 216496 3528
rect 215803 3488 216496 3516
rect 215803 3485 215815 3488
rect 215757 3479 215815 3485
rect 216490 3476 216496 3488
rect 216548 3476 216554 3528
rect 216600 3525 216628 3556
rect 217410 3544 217416 3596
rect 217468 3544 217474 3596
rect 221090 3544 221096 3596
rect 221148 3544 221154 3596
rect 221366 3544 221372 3596
rect 221424 3584 221430 3596
rect 221424 3556 222516 3584
rect 221424 3544 221430 3556
rect 216585 3519 216643 3525
rect 216585 3485 216597 3519
rect 216631 3485 216643 3519
rect 216585 3479 216643 3485
rect 216674 3476 216680 3528
rect 216732 3476 216738 3528
rect 220541 3519 220599 3525
rect 220541 3516 220553 3519
rect 218808 3488 220553 3516
rect 212552 3420 212764 3448
rect 213012 3420 213224 3448
rect 213273 3451 213331 3457
rect 211430 3380 211436 3392
rect 210344 3352 211436 3380
rect 211430 3340 211436 3352
rect 211488 3340 211494 3392
rect 211522 3340 211528 3392
rect 211580 3380 211586 3392
rect 213012 3380 213040 3420
rect 213273 3417 213285 3451
rect 213319 3448 213331 3451
rect 215110 3448 215116 3460
rect 213319 3420 215116 3448
rect 213319 3417 213331 3420
rect 213273 3411 213331 3417
rect 215110 3408 215116 3420
rect 215168 3408 215174 3460
rect 216861 3451 216919 3457
rect 216861 3417 216873 3451
rect 216907 3448 216919 3451
rect 217597 3451 217655 3457
rect 217597 3448 217609 3451
rect 216907 3420 217609 3448
rect 216907 3417 216919 3420
rect 216861 3411 216919 3417
rect 217597 3417 217609 3420
rect 217643 3417 217655 3451
rect 217597 3411 217655 3417
rect 217686 3408 217692 3460
rect 217744 3448 217750 3460
rect 218808 3448 218836 3488
rect 220541 3485 220553 3488
rect 220587 3485 220599 3519
rect 222488 3516 222516 3556
rect 222562 3544 222568 3596
rect 222620 3544 222626 3596
rect 222746 3544 222752 3596
rect 222804 3584 222810 3596
rect 222804 3556 223620 3584
rect 222804 3544 222810 3556
rect 223592 3525 223620 3556
rect 223942 3544 223948 3596
rect 224000 3584 224006 3596
rect 224129 3587 224187 3593
rect 224129 3584 224141 3587
rect 224000 3556 224141 3584
rect 224000 3544 224006 3556
rect 224129 3553 224141 3556
rect 224175 3553 224187 3587
rect 224129 3547 224187 3553
rect 224218 3544 224224 3596
rect 224276 3584 224282 3596
rect 225874 3584 225880 3596
rect 224276 3556 225880 3584
rect 224276 3544 224282 3556
rect 225874 3544 225880 3556
rect 225932 3584 225938 3596
rect 226153 3587 226211 3593
rect 226153 3584 226165 3587
rect 225932 3556 226165 3584
rect 225932 3544 225938 3556
rect 226153 3553 226165 3556
rect 226199 3553 226211 3587
rect 226153 3547 226211 3553
rect 226242 3544 226248 3596
rect 226300 3584 226306 3596
rect 226429 3587 226487 3593
rect 226429 3584 226441 3587
rect 226300 3556 226441 3584
rect 226300 3544 226306 3556
rect 226429 3553 226441 3556
rect 226475 3553 226487 3587
rect 226429 3547 226487 3553
rect 226567 3587 226625 3593
rect 226567 3553 226579 3587
rect 226613 3584 226625 3587
rect 227732 3584 227760 3624
rect 229738 3612 229744 3624
rect 229796 3612 229802 3664
rect 229830 3612 229836 3664
rect 229888 3652 229894 3664
rect 241790 3652 241796 3664
rect 229888 3624 241796 3652
rect 229888 3612 229894 3624
rect 241790 3612 241796 3624
rect 241848 3612 241854 3664
rect 244366 3612 244372 3664
rect 244424 3652 244430 3664
rect 253017 3655 253075 3661
rect 244424 3624 251588 3652
rect 244424 3612 244430 3624
rect 231854 3584 231860 3596
rect 226613 3556 227668 3584
rect 227732 3556 231860 3584
rect 226613 3553 226625 3556
rect 226567 3547 226625 3553
rect 223485 3519 223543 3525
rect 223485 3516 223497 3519
rect 222488 3488 223497 3516
rect 220541 3479 220599 3485
rect 223485 3485 223497 3488
rect 223531 3485 223543 3519
rect 223485 3479 223543 3485
rect 223577 3519 223635 3525
rect 223577 3485 223589 3519
rect 223623 3485 223635 3519
rect 223577 3479 223635 3485
rect 223758 3476 223764 3528
rect 223816 3476 223822 3528
rect 224034 3476 224040 3528
rect 224092 3516 224098 3528
rect 224589 3519 224647 3525
rect 224589 3516 224601 3519
rect 224092 3488 224601 3516
rect 224092 3476 224098 3488
rect 224589 3485 224601 3488
rect 224635 3485 224647 3519
rect 224589 3479 224647 3485
rect 225506 3476 225512 3528
rect 225564 3476 225570 3528
rect 225690 3476 225696 3528
rect 225748 3476 225754 3528
rect 226702 3476 226708 3528
rect 226760 3476 226766 3528
rect 217744 3420 218836 3448
rect 217744 3408 217750 3420
rect 219158 3408 219164 3460
rect 219216 3448 219222 3460
rect 219253 3451 219311 3457
rect 219253 3448 219265 3451
rect 219216 3420 219265 3448
rect 219216 3408 219222 3420
rect 219253 3417 219265 3420
rect 219299 3417 219311 3451
rect 219253 3411 219311 3417
rect 219618 3408 219624 3460
rect 219676 3448 219682 3460
rect 220814 3448 220820 3460
rect 219676 3420 220820 3448
rect 219676 3408 219682 3420
rect 220814 3408 220820 3420
rect 220872 3408 220878 3460
rect 220906 3408 220912 3460
rect 220964 3448 220970 3460
rect 221277 3451 221335 3457
rect 221277 3448 221289 3451
rect 220964 3420 221289 3448
rect 220964 3408 220970 3420
rect 221277 3417 221289 3420
rect 221323 3417 221335 3451
rect 221277 3411 221335 3417
rect 221458 3408 221464 3460
rect 221516 3448 221522 3460
rect 227640 3448 227668 3556
rect 231854 3544 231860 3556
rect 231912 3544 231918 3596
rect 238754 3584 238760 3596
rect 234586 3556 238760 3584
rect 227714 3476 227720 3528
rect 227772 3516 227778 3528
rect 234586 3516 234614 3556
rect 238754 3544 238760 3556
rect 238812 3544 238818 3596
rect 243998 3584 244004 3596
rect 241486 3556 244004 3584
rect 227772 3488 234614 3516
rect 227772 3476 227778 3488
rect 236270 3476 236276 3528
rect 236328 3516 236334 3528
rect 241486 3516 241514 3556
rect 243998 3544 244004 3556
rect 244056 3544 244062 3596
rect 244550 3584 244556 3596
rect 244384 3556 244556 3584
rect 244384 3525 244412 3556
rect 244550 3544 244556 3556
rect 244608 3584 244614 3596
rect 245289 3587 245347 3593
rect 245289 3584 245301 3587
rect 244608 3556 245301 3584
rect 244608 3544 244614 3556
rect 245289 3553 245301 3556
rect 245335 3584 245347 3587
rect 246393 3587 246451 3593
rect 246393 3584 246405 3587
rect 245335 3556 246405 3584
rect 245335 3553 245347 3556
rect 245289 3547 245347 3553
rect 246393 3553 246405 3556
rect 246439 3584 246451 3587
rect 246850 3584 246856 3596
rect 246439 3556 246856 3584
rect 246439 3553 246451 3556
rect 246393 3547 246451 3553
rect 246850 3544 246856 3556
rect 246908 3544 246914 3596
rect 247310 3544 247316 3596
rect 247368 3544 247374 3596
rect 248693 3587 248751 3593
rect 248693 3553 248705 3587
rect 248739 3584 248751 3587
rect 249242 3584 249248 3596
rect 248739 3556 249248 3584
rect 248739 3553 248751 3556
rect 248693 3547 248751 3553
rect 249242 3544 249248 3556
rect 249300 3544 249306 3596
rect 251560 3593 251588 3624
rect 253017 3621 253029 3655
rect 253063 3652 253075 3655
rect 253290 3652 253296 3664
rect 253063 3624 253296 3652
rect 253063 3621 253075 3624
rect 253017 3615 253075 3621
rect 253290 3612 253296 3624
rect 253348 3612 253354 3664
rect 268010 3652 268016 3664
rect 258276 3624 268016 3652
rect 251545 3587 251603 3593
rect 251545 3553 251557 3587
rect 251591 3553 251603 3587
rect 251545 3547 251603 3553
rect 251634 3544 251640 3596
rect 251692 3584 251698 3596
rect 252649 3587 252707 3593
rect 252649 3584 252661 3587
rect 251692 3556 252661 3584
rect 251692 3544 251698 3556
rect 252649 3553 252661 3556
rect 252695 3553 252707 3587
rect 252649 3547 252707 3553
rect 254026 3544 254032 3596
rect 254084 3544 254090 3596
rect 255130 3544 255136 3596
rect 255188 3584 255194 3596
rect 258276 3593 258304 3624
rect 268010 3612 268016 3624
rect 268068 3612 268074 3664
rect 268565 3655 268623 3661
rect 268565 3621 268577 3655
rect 268611 3621 268623 3655
rect 268565 3615 268623 3621
rect 255869 3587 255927 3593
rect 255188 3556 255452 3584
rect 255188 3544 255194 3556
rect 236328 3488 241514 3516
rect 244369 3519 244427 3525
rect 236328 3476 236334 3488
rect 244369 3485 244381 3519
rect 244415 3485 244427 3519
rect 244369 3479 244427 3485
rect 244461 3519 244519 3525
rect 244461 3485 244473 3519
rect 244507 3516 244519 3519
rect 245381 3519 245439 3525
rect 245381 3516 245393 3519
rect 244507 3488 245393 3516
rect 244507 3485 244519 3488
rect 244461 3479 244519 3485
rect 245381 3485 245393 3488
rect 245427 3516 245439 3519
rect 246485 3519 246543 3525
rect 246485 3516 246497 3519
rect 245427 3488 246497 3516
rect 245427 3485 245439 3488
rect 245381 3479 245439 3485
rect 246485 3485 246497 3488
rect 246531 3516 246543 3519
rect 246942 3516 246948 3528
rect 246531 3488 246948 3516
rect 246531 3485 246543 3488
rect 246485 3479 246543 3485
rect 221516 3420 224954 3448
rect 227640 3420 227760 3448
rect 221516 3408 221522 3420
rect 211580 3352 213040 3380
rect 211580 3340 211586 3352
rect 213730 3340 213736 3392
rect 213788 3340 213794 3392
rect 216582 3340 216588 3392
rect 216640 3380 216646 3392
rect 222102 3380 222108 3392
rect 216640 3352 222108 3380
rect 216640 3340 216646 3352
rect 222102 3340 222108 3352
rect 222160 3340 222166 3392
rect 223942 3340 223948 3392
rect 224000 3380 224006 3392
rect 224681 3383 224739 3389
rect 224681 3380 224693 3383
rect 224000 3352 224693 3380
rect 224000 3340 224006 3352
rect 224681 3349 224693 3352
rect 224727 3349 224739 3383
rect 224926 3380 224954 3420
rect 227732 3392 227760 3420
rect 243998 3408 244004 3460
rect 244056 3448 244062 3460
rect 244185 3451 244243 3457
rect 244185 3448 244197 3451
rect 244056 3420 244197 3448
rect 244056 3408 244062 3420
rect 244185 3417 244197 3420
rect 244231 3417 244243 3451
rect 244185 3411 244243 3417
rect 244274 3408 244280 3460
rect 244332 3448 244338 3460
rect 244476 3448 244504 3479
rect 246942 3476 246948 3488
rect 247000 3476 247006 3528
rect 247034 3476 247040 3528
rect 247092 3476 247098 3528
rect 248509 3519 248567 3525
rect 248509 3516 248521 3519
rect 248156 3488 248521 3516
rect 248156 3460 248184 3488
rect 248509 3485 248521 3488
rect 248555 3485 248567 3519
rect 248509 3479 248567 3485
rect 250990 3476 250996 3528
rect 251048 3516 251054 3528
rect 251269 3519 251327 3525
rect 251269 3516 251281 3519
rect 251048 3488 251281 3516
rect 251048 3476 251054 3488
rect 251269 3485 251281 3488
rect 251315 3485 251327 3519
rect 251269 3479 251327 3485
rect 251358 3476 251364 3528
rect 251416 3516 251422 3528
rect 252833 3519 252891 3525
rect 252833 3516 252845 3519
rect 251416 3488 252845 3516
rect 251416 3476 251422 3488
rect 252833 3485 252845 3488
rect 252879 3485 252891 3519
rect 255424 3516 255452 3556
rect 255869 3553 255881 3587
rect 255915 3584 255927 3587
rect 258261 3587 258319 3593
rect 255915 3556 258212 3584
rect 255915 3553 255927 3556
rect 255869 3547 255927 3553
rect 256421 3519 256479 3525
rect 256421 3516 256433 3519
rect 255424 3488 256433 3516
rect 252833 3479 252891 3485
rect 256421 3485 256433 3488
rect 256467 3485 256479 3519
rect 258184 3516 258212 3556
rect 258261 3553 258273 3587
rect 258307 3553 258319 3587
rect 258261 3547 258319 3553
rect 258718 3544 258724 3596
rect 258776 3584 258782 3596
rect 258813 3587 258871 3593
rect 258813 3584 258825 3587
rect 258776 3556 258825 3584
rect 258776 3544 258782 3556
rect 258813 3553 258825 3556
rect 258859 3553 258871 3587
rect 258813 3547 258871 3553
rect 258920 3556 263594 3584
rect 258920 3516 258948 3556
rect 258184 3488 258948 3516
rect 258997 3519 259055 3525
rect 256421 3479 256479 3485
rect 258997 3485 259009 3519
rect 259043 3516 259055 3519
rect 259362 3516 259368 3528
rect 259043 3488 259368 3516
rect 259043 3485 259055 3488
rect 258997 3479 259055 3485
rect 259362 3476 259368 3488
rect 259420 3476 259426 3528
rect 260377 3519 260435 3525
rect 260377 3485 260389 3519
rect 260423 3516 260435 3519
rect 260650 3516 260656 3528
rect 260423 3488 260656 3516
rect 260423 3485 260435 3488
rect 260377 3479 260435 3485
rect 260650 3476 260656 3488
rect 260708 3476 260714 3528
rect 263566 3516 263594 3556
rect 265894 3544 265900 3596
rect 265952 3584 265958 3596
rect 265989 3587 266047 3593
rect 265989 3584 266001 3587
rect 265952 3556 266001 3584
rect 265952 3544 265958 3556
rect 265989 3553 266001 3556
rect 266035 3553 266047 3587
rect 265989 3547 266047 3553
rect 266538 3544 266544 3596
rect 266596 3584 266602 3596
rect 268580 3584 268608 3615
rect 266596 3556 268608 3584
rect 266596 3544 266602 3556
rect 263566 3488 267412 3516
rect 245010 3448 245016 3460
rect 244332 3420 244504 3448
rect 244568 3420 245016 3448
rect 244332 3408 244338 3420
rect 225874 3380 225880 3392
rect 224926 3352 225880 3380
rect 224681 3343 224739 3349
rect 225874 3340 225880 3352
rect 225932 3340 225938 3392
rect 227714 3340 227720 3392
rect 227772 3340 227778 3392
rect 229738 3340 229744 3392
rect 229796 3380 229802 3392
rect 244568 3380 244596 3420
rect 245010 3408 245016 3420
rect 245068 3408 245074 3460
rect 245105 3451 245163 3457
rect 245105 3417 245117 3451
rect 245151 3448 245163 3451
rect 246209 3451 246267 3457
rect 246209 3448 246221 3451
rect 245151 3420 246221 3448
rect 245151 3417 245163 3420
rect 245105 3411 245163 3417
rect 246209 3417 246221 3420
rect 246255 3448 246267 3451
rect 246574 3448 246580 3460
rect 246255 3420 246580 3448
rect 246255 3417 246267 3420
rect 246209 3411 246267 3417
rect 229796 3352 244596 3380
rect 229796 3340 229802 3352
rect 244642 3340 244648 3392
rect 244700 3340 244706 3392
rect 244826 3340 244832 3392
rect 244884 3380 244890 3392
rect 245120 3380 245148 3411
rect 246574 3408 246580 3420
rect 246632 3448 246638 3460
rect 247218 3448 247224 3460
rect 246632 3420 247224 3448
rect 246632 3408 246638 3420
rect 247218 3408 247224 3420
rect 247276 3408 247282 3460
rect 248138 3408 248144 3460
rect 248196 3408 248202 3460
rect 250349 3451 250407 3457
rect 250349 3417 250361 3451
rect 250395 3417 250407 3451
rect 250349 3411 250407 3417
rect 252557 3451 252615 3457
rect 252557 3417 252569 3451
rect 252603 3448 252615 3451
rect 252646 3448 252652 3460
rect 252603 3420 252652 3448
rect 252603 3417 252615 3420
rect 252557 3411 252615 3417
rect 244884 3352 245148 3380
rect 244884 3340 244890 3352
rect 245562 3340 245568 3392
rect 245620 3340 245626 3392
rect 248414 3340 248420 3392
rect 248472 3380 248478 3392
rect 249610 3380 249616 3392
rect 248472 3352 249616 3380
rect 248472 3340 248478 3352
rect 249610 3340 249616 3352
rect 249668 3340 249674 3392
rect 250364 3380 250392 3411
rect 252646 3408 252652 3420
rect 252704 3408 252710 3460
rect 252940 3420 253152 3448
rect 252940 3380 252968 3420
rect 250364 3352 252968 3380
rect 253124 3380 253152 3420
rect 253934 3408 253940 3460
rect 253992 3448 253998 3460
rect 254213 3451 254271 3457
rect 254213 3448 254225 3451
rect 253992 3420 254225 3448
rect 253992 3408 253998 3420
rect 254213 3417 254225 3420
rect 254259 3417 254271 3451
rect 254213 3411 254271 3417
rect 254302 3408 254308 3460
rect 254360 3448 254366 3460
rect 256605 3451 256663 3457
rect 256605 3448 256617 3451
rect 254360 3420 256617 3448
rect 254360 3408 254366 3420
rect 256605 3417 256617 3420
rect 256651 3417 256663 3451
rect 256605 3411 256663 3417
rect 258721 3451 258779 3457
rect 258721 3417 258733 3451
rect 258767 3448 258779 3451
rect 259270 3448 259276 3460
rect 258767 3420 259276 3448
rect 258767 3417 258779 3420
rect 258721 3411 258779 3417
rect 259270 3408 259276 3420
rect 259328 3408 259334 3460
rect 259730 3408 259736 3460
rect 259788 3408 259794 3460
rect 267384 3448 267412 3488
rect 267458 3476 267464 3528
rect 267516 3476 267522 3528
rect 268102 3476 268108 3528
rect 268160 3476 268166 3528
rect 268746 3476 268752 3528
rect 268804 3476 268810 3528
rect 268856 3516 268884 3680
rect 270770 3612 270776 3664
rect 270828 3652 270834 3664
rect 271782 3652 271788 3664
rect 270828 3624 271788 3652
rect 270828 3612 270834 3624
rect 271782 3612 271788 3624
rect 271840 3612 271846 3664
rect 269393 3519 269451 3525
rect 269393 3516 269405 3519
rect 268856 3488 269405 3516
rect 269393 3485 269405 3488
rect 269439 3485 269451 3519
rect 269393 3479 269451 3485
rect 269853 3519 269911 3525
rect 269853 3485 269865 3519
rect 269899 3516 269911 3519
rect 270586 3516 270592 3528
rect 269899 3488 270592 3516
rect 269899 3485 269911 3488
rect 269853 3479 269911 3485
rect 270586 3476 270592 3488
rect 270644 3476 270650 3528
rect 270957 3519 271015 3525
rect 270957 3485 270969 3519
rect 271003 3516 271015 3519
rect 271874 3516 271880 3528
rect 271003 3488 271880 3516
rect 271003 3485 271015 3488
rect 270957 3479 271015 3485
rect 271874 3476 271880 3488
rect 271932 3476 271938 3528
rect 267918 3448 267924 3460
rect 265452 3420 267320 3448
rect 267384 3420 267924 3448
rect 254118 3380 254124 3392
rect 253124 3352 254124 3380
rect 254118 3340 254124 3352
rect 254176 3340 254182 3392
rect 258902 3340 258908 3392
rect 258960 3380 258966 3392
rect 259181 3383 259239 3389
rect 259181 3380 259193 3383
rect 258960 3352 259193 3380
rect 258960 3340 258966 3352
rect 259181 3349 259193 3352
rect 259227 3349 259239 3383
rect 259181 3343 259239 3349
rect 259825 3383 259883 3389
rect 259825 3349 259837 3383
rect 259871 3380 259883 3383
rect 260466 3380 260472 3392
rect 259871 3352 260472 3380
rect 259871 3349 259883 3352
rect 259825 3343 259883 3349
rect 260466 3340 260472 3352
rect 260524 3340 260530 3392
rect 262122 3340 262128 3392
rect 262180 3380 262186 3392
rect 265452 3380 265480 3420
rect 267292 3389 267320 3420
rect 267918 3408 267924 3420
rect 267976 3408 267982 3460
rect 271230 3448 271236 3460
rect 270788 3420 271236 3448
rect 262180 3352 265480 3380
rect 267277 3383 267335 3389
rect 262180 3340 262186 3352
rect 267277 3349 267289 3383
rect 267323 3349 267335 3383
rect 267277 3343 267335 3349
rect 267734 3340 267740 3392
rect 267792 3380 267798 3392
rect 268930 3380 268936 3392
rect 267792 3352 268936 3380
rect 267792 3340 267798 3352
rect 268930 3340 268936 3352
rect 268988 3340 268994 3392
rect 270788 3389 270816 3420
rect 271230 3408 271236 3420
rect 271288 3408 271294 3460
rect 270773 3383 270831 3389
rect 270773 3349 270785 3383
rect 270819 3349 270831 3383
rect 270773 3343 270831 3349
rect 271138 3340 271144 3392
rect 271196 3380 271202 3392
rect 272150 3380 272156 3392
rect 271196 3352 272156 3380
rect 271196 3340 271202 3352
rect 272150 3340 272156 3352
rect 272208 3340 272214 3392
rect 1104 3290 271651 3312
rect 1104 3238 68546 3290
rect 68598 3238 68610 3290
rect 68662 3238 68674 3290
rect 68726 3238 68738 3290
rect 68790 3238 68802 3290
rect 68854 3238 136143 3290
rect 136195 3238 136207 3290
rect 136259 3238 136271 3290
rect 136323 3238 136335 3290
rect 136387 3238 136399 3290
rect 136451 3238 203740 3290
rect 203792 3238 203804 3290
rect 203856 3238 203868 3290
rect 203920 3238 203932 3290
rect 203984 3238 203996 3290
rect 204048 3238 271337 3290
rect 271389 3238 271401 3290
rect 271453 3238 271465 3290
rect 271517 3238 271529 3290
rect 271581 3238 271593 3290
rect 271645 3238 271651 3290
rect 1104 3216 271651 3238
rect 23474 3136 23480 3188
rect 23532 3176 23538 3188
rect 38749 3179 38807 3185
rect 38749 3176 38761 3179
rect 23532 3148 38761 3176
rect 23532 3136 23538 3148
rect 38749 3145 38761 3148
rect 38795 3145 38807 3179
rect 38749 3139 38807 3145
rect 38933 3179 38991 3185
rect 38933 3145 38945 3179
rect 38979 3176 38991 3179
rect 39114 3176 39120 3188
rect 38979 3148 39120 3176
rect 38979 3145 38991 3148
rect 38933 3139 38991 3145
rect 39114 3136 39120 3148
rect 39172 3136 39178 3188
rect 39482 3136 39488 3188
rect 39540 3176 39546 3188
rect 42426 3176 42432 3188
rect 39540 3148 42432 3176
rect 39540 3136 39546 3148
rect 42426 3136 42432 3148
rect 42484 3136 42490 3188
rect 42536 3148 43760 3176
rect 24946 3068 24952 3120
rect 25004 3108 25010 3120
rect 25004 3080 37596 3108
rect 25004 3068 25010 3080
rect 22094 3000 22100 3052
rect 22152 3040 22158 3052
rect 22649 3043 22707 3049
rect 22649 3040 22661 3043
rect 22152 3012 22661 3040
rect 22152 3000 22158 3012
rect 22649 3009 22661 3012
rect 22695 3009 22707 3043
rect 22649 3003 22707 3009
rect 22833 3043 22891 3049
rect 22833 3009 22845 3043
rect 22879 3040 22891 3043
rect 23290 3040 23296 3052
rect 22879 3012 23296 3040
rect 22879 3009 22891 3012
rect 22833 3003 22891 3009
rect 23290 3000 23296 3012
rect 23348 3000 23354 3052
rect 23658 3000 23664 3052
rect 23716 3000 23722 3052
rect 24486 3000 24492 3052
rect 24544 3000 24550 3052
rect 24578 3000 24584 3052
rect 24636 3000 24642 3052
rect 25406 3000 25412 3052
rect 25464 3040 25470 3052
rect 25593 3043 25651 3049
rect 25593 3040 25605 3043
rect 25464 3012 25605 3040
rect 25464 3000 25470 3012
rect 25593 3009 25605 3012
rect 25639 3009 25651 3043
rect 25593 3003 25651 3009
rect 26234 3000 26240 3052
rect 26292 3040 26298 3052
rect 26329 3043 26387 3049
rect 26329 3040 26341 3043
rect 26292 3012 26341 3040
rect 26292 3000 26298 3012
rect 26329 3009 26341 3012
rect 26375 3009 26387 3043
rect 37568 3040 37596 3080
rect 37642 3068 37648 3120
rect 37700 3068 37706 3120
rect 37918 3068 37924 3120
rect 37976 3068 37982 3120
rect 38010 3068 38016 3120
rect 38068 3068 38074 3120
rect 39206 3068 39212 3120
rect 39264 3108 39270 3120
rect 42536 3108 42564 3148
rect 42981 3111 43039 3117
rect 39264 3080 42564 3108
rect 42720 3080 42932 3108
rect 39264 3068 39270 3080
rect 38381 3043 38439 3049
rect 38381 3040 38393 3043
rect 37568 3012 38393 3040
rect 26329 3003 26387 3009
rect 38381 3009 38393 3012
rect 38427 3009 38439 3043
rect 38381 3003 38439 3009
rect 38562 3000 38568 3052
rect 38620 3040 38626 3052
rect 42720 3040 42748 3080
rect 38620 3012 42748 3040
rect 42904 3040 42932 3080
rect 42981 3077 42993 3111
rect 43027 3108 43039 3111
rect 43162 3108 43168 3120
rect 43027 3080 43168 3108
rect 43027 3077 43039 3080
rect 42981 3071 43039 3077
rect 43162 3068 43168 3080
rect 43220 3068 43226 3120
rect 43254 3068 43260 3120
rect 43312 3068 43318 3120
rect 43346 3068 43352 3120
rect 43404 3068 43410 3120
rect 43732 3117 43760 3148
rect 44082 3136 44088 3188
rect 44140 3136 44146 3188
rect 44269 3179 44327 3185
rect 44269 3145 44281 3179
rect 44315 3176 44327 3179
rect 47486 3176 47492 3188
rect 44315 3148 47492 3176
rect 44315 3145 44327 3148
rect 44269 3139 44327 3145
rect 47486 3136 47492 3148
rect 47544 3136 47550 3188
rect 49510 3136 49516 3188
rect 49568 3176 49574 3188
rect 93026 3176 93032 3188
rect 49568 3148 93032 3176
rect 49568 3136 49574 3148
rect 93026 3136 93032 3148
rect 93084 3136 93090 3188
rect 93302 3136 93308 3188
rect 93360 3176 93366 3188
rect 93360 3148 95372 3176
rect 93360 3136 93366 3148
rect 43717 3111 43775 3117
rect 43717 3077 43729 3111
rect 43763 3077 43775 3111
rect 43717 3071 43775 3077
rect 47946 3068 47952 3120
rect 48004 3068 48010 3120
rect 49050 3068 49056 3120
rect 49108 3068 49114 3120
rect 51810 3068 51816 3120
rect 51868 3108 51874 3120
rect 91186 3108 91192 3120
rect 51868 3080 91192 3108
rect 51868 3068 51874 3080
rect 91186 3068 91192 3080
rect 91244 3068 91250 3120
rect 95237 3111 95295 3117
rect 95237 3108 95249 3111
rect 93320 3080 95249 3108
rect 42904 3012 44128 3040
rect 38620 3000 38626 3012
rect 31938 2932 31944 2984
rect 31996 2972 32002 2984
rect 32309 2975 32367 2981
rect 32309 2972 32321 2975
rect 31996 2944 32321 2972
rect 31996 2932 32002 2944
rect 32309 2941 32321 2944
rect 32355 2941 32367 2975
rect 32309 2935 32367 2941
rect 38470 2932 38476 2984
rect 38528 2932 38534 2984
rect 40586 2932 40592 2984
rect 40644 2972 40650 2984
rect 41138 2972 41144 2984
rect 40644 2944 41144 2972
rect 40644 2932 40650 2944
rect 41138 2932 41144 2944
rect 41196 2932 41202 2984
rect 43806 2932 43812 2984
rect 43864 2932 43870 2984
rect 44100 2972 44128 3012
rect 48038 3000 48044 3052
rect 48096 3040 48102 3052
rect 48218 3043 48276 3049
rect 48218 3040 48230 3043
rect 48096 3012 48230 3040
rect 48096 3000 48102 3012
rect 48218 3009 48230 3012
rect 48264 3009 48276 3043
rect 48218 3003 48276 3009
rect 48317 3043 48375 3049
rect 48317 3009 48329 3043
rect 48363 3040 48375 3043
rect 48498 3040 48504 3052
rect 48363 3012 48504 3040
rect 48363 3009 48375 3012
rect 48317 3003 48375 3009
rect 48498 3000 48504 3012
rect 48556 3000 48562 3052
rect 48682 3000 48688 3052
rect 48740 3000 48746 3052
rect 49142 3000 49148 3052
rect 49200 3040 49206 3052
rect 49605 3043 49663 3049
rect 49605 3040 49617 3043
rect 49200 3012 49617 3040
rect 49200 3000 49206 3012
rect 49605 3009 49617 3012
rect 49651 3009 49663 3043
rect 49605 3003 49663 3009
rect 54297 3043 54355 3049
rect 54297 3009 54309 3043
rect 54343 3040 54355 3043
rect 54662 3040 54668 3052
rect 54343 3012 54668 3040
rect 54343 3009 54355 3012
rect 54297 3003 54355 3009
rect 54662 3000 54668 3012
rect 54720 3000 54726 3052
rect 89346 3000 89352 3052
rect 89404 3000 89410 3052
rect 90637 3043 90695 3049
rect 90637 3009 90649 3043
rect 90683 3040 90695 3043
rect 90910 3040 90916 3052
rect 90683 3012 90916 3040
rect 90683 3009 90695 3012
rect 90637 3003 90695 3009
rect 90910 3000 90916 3012
rect 90968 3000 90974 3052
rect 91830 3000 91836 3052
rect 91888 3000 91894 3052
rect 93320 3049 93348 3080
rect 95237 3077 95249 3080
rect 95283 3077 95295 3111
rect 95344 3108 95372 3148
rect 96430 3136 96436 3188
rect 96488 3136 96494 3188
rect 96522 3136 96528 3188
rect 96580 3176 96586 3188
rect 96580 3148 97212 3176
rect 96580 3136 96586 3148
rect 97077 3111 97135 3117
rect 97077 3108 97089 3111
rect 95344 3080 97089 3108
rect 95237 3071 95295 3077
rect 97077 3077 97089 3080
rect 97123 3077 97135 3111
rect 97184 3108 97212 3148
rect 97258 3136 97264 3188
rect 97316 3176 97322 3188
rect 97626 3176 97632 3188
rect 97316 3148 97632 3176
rect 97316 3136 97322 3148
rect 97626 3136 97632 3148
rect 97684 3136 97690 3188
rect 97902 3136 97908 3188
rect 97960 3176 97966 3188
rect 97960 3148 104664 3176
rect 97960 3136 97966 3148
rect 97184 3080 99374 3108
rect 97077 3071 97135 3077
rect 92569 3043 92627 3049
rect 92569 3009 92581 3043
rect 92615 3009 92627 3043
rect 92569 3003 92627 3009
rect 93305 3043 93363 3049
rect 93305 3009 93317 3043
rect 93351 3009 93363 3043
rect 93305 3003 93363 3009
rect 47768 2984 47820 2990
rect 47670 2972 47676 2984
rect 44100 2944 47676 2972
rect 47670 2932 47676 2944
rect 47728 2932 47734 2984
rect 66346 2932 66352 2984
rect 66404 2932 66410 2984
rect 92584 2972 92612 3003
rect 94130 3000 94136 3052
rect 94188 3000 94194 3052
rect 94314 3000 94320 3052
rect 94372 3040 94378 3052
rect 94498 3040 94504 3052
rect 94372 3012 94504 3040
rect 94372 3000 94378 3012
rect 94498 3000 94504 3012
rect 94556 3000 94562 3052
rect 94958 3000 94964 3052
rect 95016 3000 95022 3052
rect 95053 3043 95111 3049
rect 95053 3009 95065 3043
rect 95099 3040 95111 3043
rect 96249 3043 96307 3049
rect 96249 3040 96261 3043
rect 95099 3012 96261 3040
rect 95099 3009 95111 3012
rect 95053 3003 95111 3009
rect 96249 3009 96261 3012
rect 96295 3040 96307 3043
rect 96338 3040 96344 3052
rect 96295 3012 96344 3040
rect 96295 3009 96307 3012
rect 96249 3003 96307 3009
rect 96338 3000 96344 3012
rect 96396 3040 96402 3052
rect 96396 3012 96568 3040
rect 96396 3000 96402 3012
rect 93394 2972 93400 2984
rect 92584 2944 93400 2972
rect 93394 2932 93400 2944
rect 93452 2932 93458 2984
rect 96065 2975 96123 2981
rect 96065 2941 96077 2975
rect 96111 2972 96123 2975
rect 96154 2972 96160 2984
rect 96111 2944 96160 2972
rect 96111 2941 96123 2944
rect 96065 2935 96123 2941
rect 96154 2932 96160 2944
rect 96212 2932 96218 2984
rect 47768 2926 47820 2932
rect 19242 2864 19248 2916
rect 19300 2904 19306 2916
rect 25958 2904 25964 2916
rect 19300 2876 25964 2904
rect 19300 2864 19306 2876
rect 25958 2864 25964 2876
rect 26016 2864 26022 2916
rect 44174 2864 44180 2916
rect 44232 2904 44238 2916
rect 44637 2907 44695 2913
rect 44637 2904 44649 2907
rect 44232 2876 44649 2904
rect 44232 2864 44238 2876
rect 44637 2873 44649 2876
rect 44683 2873 44695 2907
rect 44637 2867 44695 2873
rect 49234 2864 49240 2916
rect 49292 2864 49298 2916
rect 93489 2907 93547 2913
rect 93489 2873 93501 2907
rect 93535 2904 93547 2907
rect 95418 2904 95424 2916
rect 93535 2876 95424 2904
rect 93535 2873 93547 2876
rect 93489 2867 93547 2873
rect 95418 2864 95424 2876
rect 95476 2864 95482 2916
rect 95694 2864 95700 2916
rect 95752 2904 95758 2916
rect 96430 2904 96436 2916
rect 95752 2876 96436 2904
rect 95752 2864 95758 2876
rect 96430 2864 96436 2876
rect 96488 2864 96494 2916
rect 96540 2904 96568 3012
rect 96614 3000 96620 3052
rect 96672 3040 96678 3052
rect 96893 3043 96951 3049
rect 96893 3040 96905 3043
rect 96672 3012 96905 3040
rect 96672 3000 96678 3012
rect 96893 3009 96905 3012
rect 96939 3009 96951 3043
rect 99346 3040 99374 3080
rect 99742 3068 99748 3120
rect 99800 3068 99806 3120
rect 101582 3068 101588 3120
rect 101640 3108 101646 3120
rect 102045 3111 102103 3117
rect 102045 3108 102057 3111
rect 101640 3080 102057 3108
rect 101640 3068 101646 3080
rect 102045 3077 102057 3080
rect 102091 3077 102103 3111
rect 102045 3071 102103 3077
rect 103698 3068 103704 3120
rect 103756 3068 103762 3120
rect 99561 3043 99619 3049
rect 99561 3040 99573 3043
rect 99346 3012 99573 3040
rect 96893 3003 96951 3009
rect 99561 3009 99573 3012
rect 99607 3009 99619 3043
rect 99561 3003 99619 3009
rect 103606 3000 103612 3052
rect 103664 3040 103670 3052
rect 104636 3049 104664 3148
rect 104986 3136 104992 3188
rect 105044 3176 105050 3188
rect 106182 3176 106188 3188
rect 105044 3148 106188 3176
rect 105044 3136 105050 3148
rect 106182 3136 106188 3148
rect 106240 3136 106246 3188
rect 106274 3136 106280 3188
rect 106332 3136 106338 3188
rect 107381 3111 107439 3117
rect 107381 3108 107393 3111
rect 106200 3080 107393 3108
rect 104437 3043 104495 3049
rect 104437 3040 104449 3043
rect 103664 3012 104449 3040
rect 103664 3000 103670 3012
rect 104437 3009 104449 3012
rect 104483 3009 104495 3043
rect 104437 3003 104495 3009
rect 104621 3043 104679 3049
rect 104621 3009 104633 3043
rect 104667 3009 104679 3043
rect 104621 3003 104679 3009
rect 105354 3000 105360 3052
rect 105412 3000 105418 3052
rect 105630 3000 105636 3052
rect 105688 3000 105694 3052
rect 98733 2975 98791 2981
rect 98733 2941 98745 2975
rect 98779 2972 98791 2975
rect 99006 2972 99012 2984
rect 98779 2944 99012 2972
rect 98779 2941 98791 2944
rect 98733 2935 98791 2941
rect 99006 2932 99012 2944
rect 99064 2932 99070 2984
rect 101401 2975 101459 2981
rect 101401 2941 101413 2975
rect 101447 2941 101459 2975
rect 101401 2935 101459 2941
rect 99374 2904 99380 2916
rect 96540 2876 99380 2904
rect 99374 2864 99380 2876
rect 99432 2864 99438 2916
rect 101416 2904 101444 2935
rect 101490 2932 101496 2984
rect 101548 2972 101554 2984
rect 101861 2975 101919 2981
rect 101861 2972 101873 2975
rect 101548 2944 101873 2972
rect 101548 2932 101554 2944
rect 101861 2941 101873 2944
rect 101907 2941 101919 2975
rect 101861 2935 101919 2941
rect 105446 2932 105452 2984
rect 105504 2981 105510 2984
rect 105504 2975 105532 2981
rect 105520 2941 105532 2975
rect 106200 2972 106228 3080
rect 107381 3077 107393 3080
rect 107427 3077 107439 3111
rect 110156 3109 110368 3137
rect 113358 3136 113364 3188
rect 113416 3176 113422 3188
rect 147214 3176 147220 3188
rect 113416 3148 147220 3176
rect 113416 3136 113422 3148
rect 147214 3136 147220 3148
rect 147272 3136 147278 3188
rect 148045 3179 148103 3185
rect 148045 3145 148057 3179
rect 148091 3176 148103 3179
rect 148091 3148 150204 3176
rect 148091 3145 148103 3148
rect 148045 3139 148103 3145
rect 110156 3108 110184 3109
rect 107381 3071 107439 3077
rect 109512 3080 110184 3108
rect 110340 3108 110368 3109
rect 110340 3080 138014 3108
rect 105504 2935 105532 2941
rect 106016 2944 106228 2972
rect 105504 2932 105510 2935
rect 104986 2904 104992 2916
rect 101416 2876 104992 2904
rect 104986 2864 104992 2876
rect 105044 2864 105050 2916
rect 105081 2907 105139 2913
rect 105081 2873 105093 2907
rect 105127 2904 105139 2907
rect 105170 2904 105176 2916
rect 105127 2876 105176 2904
rect 105127 2873 105139 2876
rect 105081 2867 105139 2873
rect 105170 2864 105176 2876
rect 105228 2864 105234 2916
rect 22094 2796 22100 2848
rect 22152 2836 22158 2848
rect 23017 2839 23075 2845
rect 23017 2836 23029 2839
rect 22152 2808 23029 2836
rect 22152 2796 22158 2808
rect 23017 2805 23029 2808
rect 23063 2805 23075 2839
rect 23017 2799 23075 2805
rect 23842 2796 23848 2848
rect 23900 2796 23906 2848
rect 24394 2796 24400 2848
rect 24452 2836 24458 2848
rect 24765 2839 24823 2845
rect 24765 2836 24777 2839
rect 24452 2808 24777 2836
rect 24452 2796 24458 2808
rect 24765 2805 24777 2808
rect 24811 2805 24823 2839
rect 24765 2799 24823 2805
rect 25774 2796 25780 2848
rect 25832 2796 25838 2848
rect 26510 2796 26516 2848
rect 26568 2796 26574 2848
rect 54478 2796 54484 2848
rect 54536 2796 54542 2848
rect 89530 2796 89536 2848
rect 89588 2796 89594 2848
rect 90818 2796 90824 2848
rect 90876 2796 90882 2848
rect 92014 2796 92020 2848
rect 92072 2796 92078 2848
rect 92750 2796 92756 2848
rect 92808 2796 92814 2848
rect 94317 2839 94375 2845
rect 94317 2805 94329 2839
rect 94363 2836 94375 2839
rect 96982 2836 96988 2848
rect 94363 2808 96988 2836
rect 94363 2805 94375 2808
rect 94317 2799 94375 2805
rect 96982 2796 96988 2808
rect 97040 2796 97046 2848
rect 97350 2796 97356 2848
rect 97408 2836 97414 2848
rect 104342 2836 104348 2848
rect 97408 2808 104348 2836
rect 97408 2796 97414 2808
rect 104342 2796 104348 2808
rect 104400 2796 104406 2848
rect 104710 2796 104716 2848
rect 104768 2836 104774 2848
rect 106016 2836 106044 2944
rect 106458 2932 106464 2984
rect 106516 2972 106522 2984
rect 107197 2975 107255 2981
rect 107197 2972 107209 2975
rect 106516 2944 107209 2972
rect 106516 2932 106522 2944
rect 107197 2941 107209 2944
rect 107243 2941 107255 2975
rect 107197 2935 107255 2941
rect 108942 2932 108948 2984
rect 109000 2932 109006 2984
rect 106366 2864 106372 2916
rect 106424 2904 106430 2916
rect 108960 2904 108988 2932
rect 106424 2876 108988 2904
rect 106424 2864 106430 2876
rect 104768 2808 106044 2836
rect 104768 2796 104774 2808
rect 106182 2796 106188 2848
rect 106240 2836 106246 2848
rect 109512 2836 109540 3080
rect 109773 3043 109831 3049
rect 109773 3009 109785 3043
rect 109819 3009 109831 3043
rect 109773 3003 109831 3009
rect 109788 2972 109816 3003
rect 110230 3000 110236 3052
rect 110288 3000 110294 3052
rect 110340 3012 110828 3040
rect 110340 2972 110368 3012
rect 109788 2944 110368 2972
rect 110506 2932 110512 2984
rect 110564 2932 110570 2984
rect 110414 2864 110420 2916
rect 110472 2904 110478 2916
rect 110800 2913 110828 3012
rect 115014 3000 115020 3052
rect 115072 3000 115078 3052
rect 119246 3000 119252 3052
rect 119304 3040 119310 3052
rect 119341 3043 119399 3049
rect 119341 3040 119353 3043
rect 119304 3012 119353 3040
rect 119304 3000 119310 3012
rect 119341 3009 119353 3012
rect 119387 3009 119399 3043
rect 119341 3003 119399 3009
rect 119982 3000 119988 3052
rect 120040 3000 120046 3052
rect 111610 2932 111616 2984
rect 111668 2972 111674 2984
rect 111797 2975 111855 2981
rect 111797 2972 111809 2975
rect 111668 2944 111809 2972
rect 111668 2932 111674 2944
rect 111797 2941 111809 2944
rect 111843 2941 111855 2975
rect 111797 2935 111855 2941
rect 111981 2975 112039 2981
rect 111981 2941 111993 2975
rect 112027 2941 112039 2975
rect 111981 2935 112039 2941
rect 110785 2907 110843 2913
rect 110472 2876 110552 2904
rect 110472 2864 110478 2876
rect 106240 2808 109540 2836
rect 106240 2796 106246 2808
rect 109586 2796 109592 2848
rect 109644 2796 109650 2848
rect 110524 2845 110552 2876
rect 110785 2873 110797 2907
rect 110831 2873 110843 2907
rect 110785 2867 110843 2873
rect 111702 2864 111708 2916
rect 111760 2904 111766 2916
rect 111996 2904 112024 2935
rect 113450 2932 113456 2984
rect 113508 2932 113514 2984
rect 115198 2932 115204 2984
rect 115256 2932 115262 2984
rect 116857 2975 116915 2981
rect 116857 2941 116869 2975
rect 116903 2941 116915 2975
rect 116857 2935 116915 2941
rect 111760 2876 112024 2904
rect 116872 2904 116900 2935
rect 117498 2932 117504 2984
rect 117556 2932 117562 2984
rect 117685 2975 117743 2981
rect 117685 2941 117697 2975
rect 117731 2972 117743 2975
rect 118602 2972 118608 2984
rect 117731 2944 118608 2972
rect 117731 2941 117743 2944
rect 117685 2935 117743 2941
rect 118602 2932 118608 2944
rect 118660 2932 118666 2984
rect 118970 2932 118976 2984
rect 119028 2972 119034 2984
rect 120169 2975 120227 2981
rect 120169 2972 120181 2975
rect 119028 2944 120181 2972
rect 119028 2932 119034 2944
rect 120169 2941 120181 2944
rect 120215 2941 120227 2975
rect 120169 2935 120227 2941
rect 120718 2932 120724 2984
rect 120776 2932 120782 2984
rect 120905 2975 120963 2981
rect 120905 2941 120917 2975
rect 120951 2972 120963 2975
rect 121638 2972 121644 2984
rect 120951 2944 121644 2972
rect 120951 2941 120963 2944
rect 120905 2935 120963 2941
rect 121638 2932 121644 2944
rect 121696 2932 121702 2984
rect 121825 2975 121883 2981
rect 121825 2941 121837 2975
rect 121871 2941 121883 2975
rect 121825 2935 121883 2941
rect 121730 2904 121736 2916
rect 116872 2876 121736 2904
rect 111760 2864 111766 2876
rect 121730 2864 121736 2876
rect 121788 2904 121794 2916
rect 121840 2904 121868 2935
rect 135346 2932 135352 2984
rect 135404 2932 135410 2984
rect 137986 2972 138014 3080
rect 138290 3068 138296 3120
rect 138348 3108 138354 3120
rect 140685 3111 140743 3117
rect 140685 3108 140697 3111
rect 138348 3080 140697 3108
rect 138348 3068 138354 3080
rect 140685 3077 140697 3080
rect 140731 3077 140743 3111
rect 140685 3071 140743 3077
rect 140866 3068 140872 3120
rect 140924 3108 140930 3120
rect 143077 3111 143135 3117
rect 143077 3108 143089 3111
rect 140924 3080 143089 3108
rect 140924 3068 140930 3080
rect 143077 3077 143089 3080
rect 143123 3077 143135 3111
rect 143077 3071 143135 3077
rect 145650 3068 145656 3120
rect 145708 3108 145714 3120
rect 145837 3111 145895 3117
rect 145837 3108 145849 3111
rect 145708 3080 145849 3108
rect 145708 3068 145714 3080
rect 145837 3077 145849 3080
rect 145883 3077 145895 3111
rect 145837 3071 145895 3077
rect 138385 3043 138443 3049
rect 138385 3009 138397 3043
rect 138431 3040 138443 3043
rect 138934 3040 138940 3052
rect 138431 3012 138940 3040
rect 138431 3009 138443 3012
rect 138385 3003 138443 3009
rect 138934 3000 138940 3012
rect 138992 3000 138998 3052
rect 139026 3000 139032 3052
rect 139084 3000 139090 3052
rect 139670 3000 139676 3052
rect 139728 3000 139734 3052
rect 148226 3000 148232 3052
rect 148284 3040 148290 3052
rect 148413 3043 148471 3049
rect 148413 3040 148425 3043
rect 148284 3012 148425 3040
rect 148284 3000 148290 3012
rect 148413 3009 148425 3012
rect 148459 3009 148471 3043
rect 148413 3003 148471 3009
rect 149330 3000 149336 3052
rect 149388 3000 149394 3052
rect 149606 3000 149612 3052
rect 149664 3000 149670 3052
rect 139946 2972 139952 2984
rect 137986 2944 139952 2972
rect 139946 2932 139952 2944
rect 140004 2932 140010 2984
rect 140501 2975 140559 2981
rect 140501 2941 140513 2975
rect 140547 2972 140559 2975
rect 141142 2972 141148 2984
rect 140547 2944 141148 2972
rect 140547 2941 140559 2944
rect 140501 2935 140559 2941
rect 141142 2932 141148 2944
rect 141200 2932 141206 2984
rect 142062 2932 142068 2984
rect 142120 2932 142126 2984
rect 142893 2975 142951 2981
rect 142893 2941 142905 2975
rect 142939 2941 142951 2975
rect 142893 2935 142951 2941
rect 121788 2876 121868 2904
rect 121788 2864 121794 2876
rect 139486 2864 139492 2916
rect 139544 2864 139550 2916
rect 142908 2904 142936 2935
rect 143534 2932 143540 2984
rect 143592 2972 143598 2984
rect 144546 2972 144552 2984
rect 143592 2944 144552 2972
rect 143592 2932 143598 2944
rect 144546 2932 144552 2944
rect 144604 2932 144610 2984
rect 145653 2975 145711 2981
rect 145653 2941 145665 2975
rect 145699 2941 145711 2975
rect 145653 2935 145711 2941
rect 144638 2904 144644 2916
rect 142908 2876 144644 2904
rect 144638 2864 144644 2876
rect 144696 2864 144702 2916
rect 145668 2904 145696 2935
rect 146478 2932 146484 2984
rect 146536 2932 146542 2984
rect 148597 2975 148655 2981
rect 148597 2941 148609 2975
rect 148643 2972 148655 2975
rect 149146 2972 149152 2984
rect 148643 2944 149152 2972
rect 148643 2941 148655 2944
rect 148597 2935 148655 2941
rect 149146 2932 149152 2944
rect 149204 2932 149210 2984
rect 149471 2975 149529 2981
rect 149471 2941 149483 2975
rect 149517 2972 149529 2975
rect 150176 2972 150204 3148
rect 150434 3136 150440 3188
rect 150492 3176 150498 3188
rect 153749 3179 153807 3185
rect 153749 3176 153761 3179
rect 150492 3148 153761 3176
rect 150492 3136 150498 3148
rect 153749 3145 153761 3148
rect 153795 3145 153807 3179
rect 153749 3139 153807 3145
rect 154393 3179 154451 3185
rect 154393 3145 154405 3179
rect 154439 3176 154451 3179
rect 156230 3176 156236 3188
rect 154439 3148 156236 3176
rect 154439 3145 154451 3148
rect 154393 3139 154451 3145
rect 156230 3136 156236 3148
rect 156288 3136 156294 3188
rect 160278 3136 160284 3188
rect 160336 3176 160342 3188
rect 171778 3176 171784 3188
rect 160336 3148 171784 3176
rect 160336 3136 160342 3148
rect 171778 3136 171784 3148
rect 171836 3136 171842 3188
rect 209682 3176 209688 3188
rect 195946 3148 209688 3176
rect 152458 3068 152464 3120
rect 152516 3108 152522 3120
rect 152516 3080 153976 3108
rect 152516 3068 152522 3080
rect 152550 3000 152556 3052
rect 152608 3040 152614 3052
rect 153948 3049 153976 3080
rect 155034 3068 155040 3120
rect 155092 3108 155098 3120
rect 159358 3108 159364 3120
rect 155092 3080 159364 3108
rect 155092 3068 155098 3080
rect 159358 3068 159364 3080
rect 159416 3068 159422 3120
rect 195946 3108 195974 3148
rect 209682 3136 209688 3148
rect 209740 3136 209746 3188
rect 209774 3136 209780 3188
rect 209832 3176 209838 3188
rect 210789 3179 210847 3185
rect 210789 3176 210801 3179
rect 209832 3148 210801 3176
rect 209832 3136 209838 3148
rect 210789 3145 210801 3148
rect 210835 3145 210847 3179
rect 210789 3139 210847 3145
rect 210970 3136 210976 3188
rect 211028 3176 211034 3188
rect 211614 3176 211620 3188
rect 211028 3148 211620 3176
rect 211028 3136 211034 3148
rect 211614 3136 211620 3148
rect 211672 3176 211678 3188
rect 212994 3176 213000 3188
rect 211672 3148 213000 3176
rect 211672 3136 211678 3148
rect 212994 3136 213000 3148
rect 213052 3136 213058 3188
rect 213454 3136 213460 3188
rect 213512 3176 213518 3188
rect 213822 3176 213828 3188
rect 213512 3148 213828 3176
rect 213512 3136 213518 3148
rect 213822 3136 213828 3148
rect 213880 3136 213886 3188
rect 218790 3136 218796 3188
rect 218848 3176 218854 3188
rect 218848 3148 220860 3176
rect 218848 3136 218854 3148
rect 162136 3080 195974 3108
rect 153289 3043 153347 3049
rect 153289 3040 153301 3043
rect 152608 3012 153301 3040
rect 152608 3000 152614 3012
rect 153289 3009 153301 3012
rect 153335 3009 153347 3043
rect 153289 3003 153347 3009
rect 153933 3043 153991 3049
rect 153933 3009 153945 3043
rect 153979 3009 153991 3043
rect 153933 3003 153991 3009
rect 154577 3043 154635 3049
rect 154577 3009 154589 3043
rect 154623 3040 154635 3043
rect 154666 3040 154672 3052
rect 154623 3012 154672 3040
rect 154623 3009 154635 3012
rect 154577 3003 154635 3009
rect 154666 3000 154672 3012
rect 154724 3000 154730 3052
rect 155221 3043 155279 3049
rect 155221 3009 155233 3043
rect 155267 3009 155279 3043
rect 155221 3003 155279 3009
rect 149517 2944 150204 2972
rect 149517 2941 149529 2944
rect 149471 2935 149529 2941
rect 147398 2904 147404 2916
rect 145668 2876 147404 2904
rect 147398 2864 147404 2876
rect 147456 2864 147462 2916
rect 148502 2864 148508 2916
rect 148560 2904 148566 2916
rect 149057 2907 149115 2913
rect 149057 2904 149069 2907
rect 148560 2876 149069 2904
rect 148560 2864 148566 2876
rect 149057 2873 149069 2876
rect 149103 2873 149115 2907
rect 150176 2904 150204 2944
rect 150253 2975 150311 2981
rect 150253 2941 150265 2975
rect 150299 2972 150311 2975
rect 150805 2975 150863 2981
rect 150805 2972 150817 2975
rect 150299 2944 150817 2972
rect 150299 2941 150311 2944
rect 150253 2935 150311 2941
rect 150805 2941 150817 2944
rect 150851 2941 150863 2975
rect 150805 2935 150863 2941
rect 150989 2975 151047 2981
rect 150989 2941 151001 2975
rect 151035 2941 151047 2975
rect 150989 2935 151047 2941
rect 151004 2904 151032 2935
rect 151262 2932 151268 2984
rect 151320 2972 151326 2984
rect 152645 2975 152703 2981
rect 152645 2972 152657 2975
rect 151320 2944 152657 2972
rect 151320 2932 151326 2944
rect 152645 2941 152657 2944
rect 152691 2972 152703 2975
rect 152826 2972 152832 2984
rect 152691 2944 152832 2972
rect 152691 2941 152703 2944
rect 152645 2935 152703 2941
rect 152826 2932 152832 2944
rect 152884 2932 152890 2984
rect 153654 2932 153660 2984
rect 153712 2972 153718 2984
rect 155236 2972 155264 3003
rect 156138 3000 156144 3052
rect 156196 3000 156202 3052
rect 158441 3043 158499 3049
rect 158441 3009 158453 3043
rect 158487 3040 158499 3043
rect 159082 3040 159088 3052
rect 158487 3012 159088 3040
rect 158487 3009 158499 3012
rect 158441 3003 158499 3009
rect 159082 3000 159088 3012
rect 159140 3000 159146 3052
rect 159177 3043 159235 3049
rect 159177 3009 159189 3043
rect 159223 3040 159235 3043
rect 160278 3040 160284 3052
rect 159223 3012 160284 3040
rect 159223 3009 159235 3012
rect 159177 3003 159235 3009
rect 160278 3000 160284 3012
rect 160336 3000 160342 3052
rect 153712 2944 155264 2972
rect 153712 2932 153718 2944
rect 155770 2932 155776 2984
rect 155828 2972 155834 2984
rect 156325 2975 156383 2981
rect 156325 2972 156337 2975
rect 155828 2944 156337 2972
rect 155828 2932 155834 2944
rect 156325 2941 156337 2944
rect 156371 2941 156383 2975
rect 156325 2935 156383 2941
rect 156414 2932 156420 2984
rect 156472 2972 156478 2984
rect 156601 2975 156659 2981
rect 156601 2972 156613 2975
rect 156472 2944 156613 2972
rect 156472 2932 156478 2944
rect 156601 2941 156613 2944
rect 156647 2972 156659 2975
rect 162136 2972 162164 3080
rect 206646 3068 206652 3120
rect 206704 3108 206710 3120
rect 208854 3108 208860 3120
rect 206704 3080 208860 3108
rect 206704 3068 206710 3080
rect 165706 3000 165712 3052
rect 165764 3040 165770 3052
rect 170306 3040 170312 3052
rect 165764 3012 170312 3040
rect 165764 3000 165770 3012
rect 170306 3000 170312 3012
rect 170364 3000 170370 3052
rect 190917 3043 190975 3049
rect 190917 3009 190929 3043
rect 190963 3040 190975 3043
rect 191282 3040 191288 3052
rect 190963 3012 191288 3040
rect 190963 3009 190975 3012
rect 190917 3003 190975 3009
rect 191282 3000 191288 3012
rect 191340 3000 191346 3052
rect 206554 3000 206560 3052
rect 206612 3040 206618 3052
rect 207768 3049 207796 3080
rect 208854 3068 208860 3080
rect 208912 3068 208918 3120
rect 211982 3068 211988 3120
rect 212040 3108 212046 3120
rect 212813 3111 212871 3117
rect 212813 3108 212825 3111
rect 212040 3080 212825 3108
rect 212040 3068 212046 3080
rect 212813 3077 212825 3080
rect 212859 3077 212871 3111
rect 212813 3071 212871 3077
rect 215110 3068 215116 3120
rect 215168 3068 215174 3120
rect 216766 3068 216772 3120
rect 216824 3108 216830 3120
rect 218422 3108 218428 3120
rect 216824 3080 218428 3108
rect 216824 3068 216830 3080
rect 218422 3068 218428 3080
rect 218480 3068 218486 3120
rect 220832 3108 220860 3148
rect 220906 3136 220912 3188
rect 220964 3136 220970 3188
rect 221016 3148 225644 3176
rect 221016 3108 221044 3148
rect 220832 3080 221044 3108
rect 222166 3080 223620 3108
rect 207661 3043 207719 3049
rect 207661 3040 207673 3043
rect 206612 3012 207673 3040
rect 206612 3000 206618 3012
rect 207661 3009 207673 3012
rect 207707 3009 207719 3043
rect 207661 3003 207719 3009
rect 207753 3043 207811 3049
rect 207753 3009 207765 3043
rect 207799 3009 207811 3043
rect 207753 3003 207811 3009
rect 156647 2944 162164 2972
rect 156647 2941 156659 2944
rect 156601 2935 156659 2941
rect 167914 2932 167920 2984
rect 167972 2932 167978 2984
rect 203150 2932 203156 2984
rect 203208 2932 203214 2984
rect 207676 2972 207704 3003
rect 207934 3000 207940 3052
rect 207992 3000 207998 3052
rect 208762 3000 208768 3052
rect 208820 3040 208826 3052
rect 208949 3043 209007 3049
rect 208949 3040 208961 3043
rect 208820 3012 208961 3040
rect 208820 3000 208826 3012
rect 208949 3009 208961 3012
rect 208995 3009 209007 3043
rect 208949 3003 209007 3009
rect 209958 3000 209964 3052
rect 210016 3049 210022 3052
rect 210016 3043 210044 3049
rect 210032 3009 210044 3043
rect 210016 3003 210044 3009
rect 210016 3000 210022 3003
rect 210142 3000 210148 3052
rect 210200 3000 210206 3052
rect 211338 3000 211344 3052
rect 211396 3000 211402 3052
rect 211430 3000 211436 3052
rect 211488 3000 211494 3052
rect 211614 3000 211620 3052
rect 211672 3000 211678 3052
rect 212350 3000 212356 3052
rect 212408 3040 212414 3052
rect 212534 3040 212540 3052
rect 212408 3012 212540 3040
rect 212408 3000 212414 3012
rect 212534 3000 212540 3012
rect 212592 3000 212598 3052
rect 220541 3043 220599 3049
rect 220541 3009 220553 3043
rect 220587 3009 220599 3043
rect 220541 3003 220599 3009
rect 208670 2972 208676 2984
rect 207676 2944 208676 2972
rect 208670 2932 208676 2944
rect 208728 2932 208734 2984
rect 209130 2932 209136 2984
rect 209188 2932 209194 2984
rect 209869 2975 209927 2981
rect 209869 2941 209881 2975
rect 209915 2972 209927 2975
rect 212629 2975 212687 2981
rect 209915 2944 210556 2972
rect 209915 2941 209927 2944
rect 209869 2935 209927 2941
rect 153105 2907 153163 2913
rect 153105 2904 153117 2907
rect 150176 2876 150480 2904
rect 151004 2876 153117 2904
rect 149057 2867 149115 2873
rect 110509 2839 110567 2845
rect 110509 2805 110521 2839
rect 110555 2805 110567 2839
rect 110509 2799 110567 2805
rect 116118 2796 116124 2848
rect 116176 2836 116182 2848
rect 120074 2836 120080 2848
rect 116176 2808 120080 2836
rect 116176 2796 116182 2808
rect 120074 2796 120080 2808
rect 120132 2796 120138 2848
rect 138198 2796 138204 2848
rect 138256 2796 138262 2848
rect 138845 2839 138903 2845
rect 138845 2805 138857 2839
rect 138891 2836 138903 2839
rect 143258 2836 143264 2848
rect 138891 2808 143264 2836
rect 138891 2805 138903 2808
rect 138845 2799 138903 2805
rect 143258 2796 143264 2808
rect 143316 2796 143322 2848
rect 145466 2796 145472 2848
rect 145524 2836 145530 2848
rect 150342 2836 150348 2848
rect 145524 2808 150348 2836
rect 145524 2796 145530 2808
rect 150342 2796 150348 2808
rect 150400 2796 150406 2848
rect 150452 2836 150480 2876
rect 153105 2873 153117 2876
rect 153151 2873 153163 2907
rect 206186 2904 206192 2916
rect 153105 2867 153163 2873
rect 153304 2876 206192 2904
rect 152918 2836 152924 2848
rect 150452 2808 152924 2836
rect 152918 2796 152924 2808
rect 152976 2796 152982 2848
rect 153010 2796 153016 2848
rect 153068 2836 153074 2848
rect 153304 2836 153332 2876
rect 206186 2864 206192 2876
rect 206244 2864 206250 2916
rect 208302 2864 208308 2916
rect 208360 2864 208366 2916
rect 209590 2904 209596 2916
rect 208412 2876 209596 2904
rect 153068 2808 153332 2836
rect 155037 2839 155095 2845
rect 153068 2796 153074 2808
rect 155037 2805 155049 2839
rect 155083 2836 155095 2839
rect 155126 2836 155132 2848
rect 155083 2808 155132 2836
rect 155083 2805 155095 2808
rect 155037 2799 155095 2805
rect 155126 2796 155132 2808
rect 155184 2796 155190 2848
rect 156230 2796 156236 2848
rect 156288 2836 156294 2848
rect 158438 2836 158444 2848
rect 156288 2808 158444 2836
rect 156288 2796 156294 2808
rect 158438 2796 158444 2808
rect 158496 2796 158502 2848
rect 158622 2796 158628 2848
rect 158680 2796 158686 2848
rect 159358 2796 159364 2848
rect 159416 2796 159422 2848
rect 191098 2796 191104 2848
rect 191156 2796 191162 2848
rect 207658 2796 207664 2848
rect 207716 2836 207722 2848
rect 208412 2836 208440 2876
rect 209590 2864 209596 2876
rect 209648 2864 209654 2916
rect 210528 2904 210556 2944
rect 212629 2941 212641 2975
rect 212675 2972 212687 2975
rect 212675 2944 212948 2972
rect 212675 2941 212687 2944
rect 212629 2935 212687 2941
rect 211154 2904 211160 2916
rect 210528 2876 211160 2904
rect 211154 2864 211160 2876
rect 211212 2864 211218 2916
rect 211893 2907 211951 2913
rect 211893 2873 211905 2907
rect 211939 2873 211951 2907
rect 212920 2904 212948 2944
rect 212994 2932 213000 2984
rect 213052 2972 213058 2984
rect 213822 2972 213828 2984
rect 213052 2944 213828 2972
rect 213052 2932 213058 2944
rect 213822 2932 213828 2944
rect 213880 2932 213886 2984
rect 214282 2932 214288 2984
rect 214340 2932 214346 2984
rect 214926 2932 214932 2984
rect 214984 2932 214990 2984
rect 215386 2932 215392 2984
rect 215444 2932 215450 2984
rect 218149 2975 218207 2981
rect 218149 2941 218161 2975
rect 218195 2941 218207 2975
rect 218149 2935 218207 2941
rect 216674 2904 216680 2916
rect 212920 2876 216680 2904
rect 211893 2867 211951 2873
rect 207716 2808 208440 2836
rect 208673 2839 208731 2845
rect 207716 2796 207722 2808
rect 208673 2805 208685 2839
rect 208719 2836 208731 2839
rect 209958 2836 209964 2848
rect 208719 2808 209964 2836
rect 208719 2805 208731 2808
rect 208673 2799 208731 2805
rect 209958 2796 209964 2808
rect 210016 2796 210022 2848
rect 211908 2836 211936 2867
rect 216674 2864 216680 2876
rect 216732 2864 216738 2916
rect 218164 2904 218192 2935
rect 218330 2932 218336 2984
rect 218388 2932 218394 2984
rect 218422 2932 218428 2984
rect 218480 2972 218486 2984
rect 219342 2972 219348 2984
rect 218480 2944 219348 2972
rect 218480 2932 218486 2944
rect 219342 2932 219348 2944
rect 219400 2932 219406 2984
rect 219618 2932 219624 2984
rect 219676 2932 219682 2984
rect 220556 2916 220584 3003
rect 220630 3000 220636 3052
rect 220688 3000 220694 3052
rect 220737 3049 220795 3055
rect 220737 3015 220749 3049
rect 220783 3046 220795 3049
rect 220783 3018 220860 3046
rect 220783 3015 220795 3018
rect 220737 3009 220795 3015
rect 220832 2984 220860 3018
rect 221366 3000 221372 3052
rect 221424 3040 221430 3052
rect 221461 3043 221519 3049
rect 221461 3040 221473 3043
rect 221424 3012 221473 3040
rect 221424 3000 221430 3012
rect 221461 3009 221473 3012
rect 221507 3009 221519 3043
rect 221461 3003 221519 3009
rect 221642 3000 221648 3052
rect 221700 3000 221706 3052
rect 221826 3000 221832 3052
rect 221884 3040 221890 3052
rect 222166 3040 222194 3080
rect 221884 3012 222194 3040
rect 221884 3000 221890 3012
rect 223390 3000 223396 3052
rect 223448 3000 223454 3052
rect 223592 3040 223620 3080
rect 225230 3068 225236 3120
rect 225288 3068 225294 3120
rect 225616 3108 225644 3148
rect 225690 3136 225696 3188
rect 225748 3136 225754 3188
rect 225782 3136 225788 3188
rect 225840 3176 225846 3188
rect 227438 3176 227444 3188
rect 225840 3148 227444 3176
rect 225840 3136 225846 3148
rect 227438 3136 227444 3148
rect 227496 3136 227502 3188
rect 227990 3136 227996 3188
rect 228048 3176 228054 3188
rect 228358 3176 228364 3188
rect 228048 3148 228364 3176
rect 228048 3136 228054 3148
rect 228358 3136 228364 3148
rect 228416 3136 228422 3188
rect 244366 3176 244372 3188
rect 234586 3148 244372 3176
rect 234586 3108 234614 3148
rect 244366 3136 244372 3148
rect 244424 3136 244430 3188
rect 244461 3179 244519 3185
rect 244461 3145 244473 3179
rect 244507 3176 244519 3179
rect 244918 3176 244924 3188
rect 244507 3148 244924 3176
rect 244507 3145 244519 3148
rect 244461 3139 244519 3145
rect 244918 3136 244924 3148
rect 244976 3136 244982 3188
rect 245010 3136 245016 3188
rect 245068 3176 245074 3188
rect 257663 3179 257721 3185
rect 257663 3176 257675 3179
rect 245068 3148 257675 3176
rect 245068 3136 245074 3148
rect 257663 3145 257675 3148
rect 257709 3145 257721 3179
rect 264238 3176 264244 3188
rect 257663 3139 257721 3145
rect 258736 3148 264244 3176
rect 225616 3080 234614 3108
rect 243998 3068 244004 3120
rect 244056 3108 244062 3120
rect 244826 3108 244832 3120
rect 244056 3080 244832 3108
rect 244056 3068 244062 3080
rect 244826 3068 244832 3080
rect 244884 3068 244890 3120
rect 245102 3068 245108 3120
rect 245160 3068 245166 3120
rect 248598 3068 248604 3120
rect 248656 3108 248662 3120
rect 248877 3111 248935 3117
rect 248877 3108 248889 3111
rect 248656 3080 248889 3108
rect 248656 3068 248662 3080
rect 248877 3077 248889 3080
rect 248923 3077 248935 3111
rect 248877 3071 248935 3077
rect 252833 3111 252891 3117
rect 252833 3077 252845 3111
rect 252879 3108 252891 3111
rect 258736 3108 258764 3148
rect 264238 3136 264244 3148
rect 264296 3136 264302 3188
rect 267274 3136 267280 3188
rect 267332 3136 267338 3188
rect 267826 3136 267832 3188
rect 267884 3176 267890 3188
rect 268565 3179 268623 3185
rect 268565 3176 268577 3179
rect 267884 3148 268577 3176
rect 267884 3136 267890 3148
rect 268565 3145 268577 3148
rect 268611 3145 268623 3179
rect 268565 3139 268623 3145
rect 269574 3136 269580 3188
rect 269632 3176 269638 3188
rect 270773 3179 270831 3185
rect 270773 3176 270785 3179
rect 269632 3148 270785 3176
rect 269632 3136 269638 3148
rect 270773 3145 270785 3148
rect 270819 3145 270831 3179
rect 270773 3139 270831 3145
rect 268010 3108 268016 3120
rect 252879 3080 258764 3108
rect 259012 3080 268016 3108
rect 252879 3077 252891 3080
rect 252833 3071 252891 3077
rect 223758 3040 223764 3052
rect 223592 3012 223764 3040
rect 223758 3000 223764 3012
rect 223816 3000 223822 3052
rect 224310 3000 224316 3052
rect 224368 3000 224374 3052
rect 224586 3000 224592 3052
rect 224644 3000 224650 3052
rect 225874 3000 225880 3052
rect 225932 3000 225938 3052
rect 225966 3000 225972 3052
rect 226024 3040 226030 3052
rect 226521 3043 226579 3049
rect 226521 3040 226533 3043
rect 226024 3012 226533 3040
rect 226024 3000 226030 3012
rect 226521 3009 226533 3012
rect 226567 3009 226579 3043
rect 226521 3003 226579 3009
rect 227714 3000 227720 3052
rect 227772 3040 227778 3052
rect 243354 3040 243360 3052
rect 227772 3012 243360 3040
rect 227772 3000 227778 3012
rect 243354 3000 243360 3012
rect 243412 3000 243418 3052
rect 244274 3000 244280 3052
rect 244332 3000 244338 3052
rect 246761 3043 246819 3049
rect 246761 3009 246773 3043
rect 246807 3040 246819 3043
rect 248414 3040 248420 3052
rect 246807 3012 248420 3040
rect 246807 3009 246819 3012
rect 246761 3003 246819 3009
rect 248414 3000 248420 3012
rect 248472 3000 248478 3052
rect 248690 3000 248696 3052
rect 248748 3000 248754 3052
rect 250070 3000 250076 3052
rect 250128 3040 250134 3052
rect 250993 3043 251051 3049
rect 250993 3040 251005 3043
rect 250128 3012 251005 3040
rect 250128 3000 250134 3012
rect 250993 3009 251005 3012
rect 251039 3009 251051 3043
rect 254121 3043 254179 3049
rect 254121 3040 254133 3043
rect 250993 3003 251051 3009
rect 252388 3012 254133 3040
rect 220814 2932 220820 2984
rect 220872 2972 220878 2984
rect 221844 2972 221872 3000
rect 220872 2944 221872 2972
rect 223577 2975 223635 2981
rect 220872 2932 220878 2944
rect 223577 2941 223589 2975
rect 223623 2941 223635 2975
rect 223577 2935 223635 2941
rect 219250 2904 219256 2916
rect 218164 2876 219256 2904
rect 219250 2864 219256 2876
rect 219308 2864 219314 2916
rect 220538 2864 220544 2916
rect 220596 2904 220602 2916
rect 221366 2904 221372 2916
rect 220596 2876 221372 2904
rect 220596 2864 220602 2876
rect 221366 2864 221372 2876
rect 221424 2864 221430 2916
rect 221476 2876 221688 2904
rect 212994 2836 213000 2848
rect 211908 2808 213000 2836
rect 212994 2796 213000 2808
rect 213052 2796 213058 2848
rect 216490 2796 216496 2848
rect 216548 2836 216554 2848
rect 217870 2836 217876 2848
rect 216548 2808 217876 2836
rect 216548 2796 216554 2808
rect 217870 2796 217876 2808
rect 217928 2836 217934 2848
rect 220556 2836 220584 2864
rect 217928 2808 220584 2836
rect 217928 2796 217934 2808
rect 220630 2796 220636 2848
rect 220688 2836 220694 2848
rect 221476 2836 221504 2876
rect 221660 2848 221688 2876
rect 220688 2808 221504 2836
rect 220688 2796 220694 2808
rect 221550 2796 221556 2848
rect 221608 2796 221614 2848
rect 221642 2796 221648 2848
rect 221700 2836 221706 2848
rect 222746 2836 222752 2848
rect 221700 2808 222752 2836
rect 221700 2796 221706 2808
rect 222746 2796 222752 2808
rect 222804 2796 222810 2848
rect 223592 2836 223620 2935
rect 223666 2932 223672 2984
rect 223724 2972 223730 2984
rect 224037 2975 224095 2981
rect 224037 2972 224049 2975
rect 223724 2944 224049 2972
rect 223724 2932 223730 2944
rect 224037 2941 224049 2944
rect 224083 2972 224095 2975
rect 224126 2972 224132 2984
rect 224083 2944 224132 2972
rect 224083 2941 224095 2944
rect 224037 2935 224095 2941
rect 224126 2932 224132 2944
rect 224184 2932 224190 2984
rect 224451 2975 224509 2981
rect 224451 2941 224463 2975
rect 224497 2972 224509 2975
rect 235721 2975 235779 2981
rect 224497 2944 225184 2972
rect 224497 2941 224509 2944
rect 224451 2935 224509 2941
rect 225156 2904 225184 2944
rect 235721 2941 235733 2975
rect 235767 2972 235779 2975
rect 235810 2972 235816 2984
rect 235767 2944 235816 2972
rect 235767 2941 235779 2944
rect 235721 2935 235779 2941
rect 235810 2932 235816 2944
rect 235868 2932 235874 2984
rect 244185 2975 244243 2981
rect 244185 2941 244197 2975
rect 244231 2941 244243 2975
rect 244185 2935 244243 2941
rect 229738 2904 229744 2916
rect 225156 2876 229744 2904
rect 229738 2864 229744 2876
rect 229796 2864 229802 2916
rect 244200 2904 244228 2935
rect 244366 2932 244372 2984
rect 244424 2972 244430 2984
rect 244921 2975 244979 2981
rect 244921 2972 244933 2975
rect 244424 2944 244933 2972
rect 244424 2932 244430 2944
rect 244921 2941 244933 2944
rect 244967 2941 244979 2975
rect 244921 2935 244979 2941
rect 246850 2932 246856 2984
rect 246908 2972 246914 2984
rect 247221 2975 247279 2981
rect 247221 2972 247233 2975
rect 246908 2944 247233 2972
rect 246908 2932 246914 2944
rect 247221 2941 247233 2944
rect 247267 2941 247279 2975
rect 247221 2935 247279 2941
rect 247402 2932 247408 2984
rect 247460 2972 247466 2984
rect 247497 2975 247555 2981
rect 247497 2972 247509 2975
rect 247460 2944 247509 2972
rect 247460 2932 247466 2944
rect 247497 2941 247509 2944
rect 247543 2941 247555 2975
rect 247497 2935 247555 2941
rect 250530 2932 250536 2984
rect 250588 2932 250594 2984
rect 251174 2932 251180 2984
rect 251232 2932 251238 2984
rect 244550 2904 244556 2916
rect 244200 2876 244556 2904
rect 244550 2864 244556 2876
rect 244608 2864 244614 2916
rect 244642 2864 244648 2916
rect 244700 2904 244706 2916
rect 252388 2904 252416 3012
rect 254121 3009 254133 3012
rect 254167 3009 254179 3043
rect 254121 3003 254179 3009
rect 256510 3000 256516 3052
rect 256568 3040 256574 3052
rect 257433 3043 257491 3049
rect 257433 3040 257445 3043
rect 256568 3012 257445 3040
rect 256568 3000 256574 3012
rect 257433 3009 257445 3012
rect 257479 3009 257491 3043
rect 259012 3040 259040 3080
rect 268010 3068 268016 3080
rect 268068 3068 268074 3120
rect 268654 3108 268660 3120
rect 268120 3080 268660 3108
rect 257433 3003 257491 3009
rect 257632 3012 259040 3040
rect 259089 3043 259147 3049
rect 253842 2932 253848 2984
rect 253900 2932 253906 2984
rect 255133 2975 255191 2981
rect 255133 2941 255145 2975
rect 255179 2941 255191 2975
rect 255133 2935 255191 2941
rect 255317 2975 255375 2981
rect 255317 2941 255329 2975
rect 255363 2941 255375 2975
rect 255317 2935 255375 2941
rect 256973 2975 257031 2981
rect 256973 2941 256985 2975
rect 257019 2972 257031 2975
rect 257632 2972 257660 3012
rect 259089 3009 259101 3043
rect 259135 3040 259147 3043
rect 259733 3043 259791 3049
rect 259733 3040 259745 3043
rect 259135 3012 259745 3040
rect 259135 3009 259147 3012
rect 259089 3003 259147 3009
rect 259733 3009 259745 3012
rect 259779 3040 259791 3043
rect 260006 3040 260012 3052
rect 259779 3012 260012 3040
rect 259779 3009 259791 3012
rect 259733 3003 259791 3009
rect 257019 2944 257660 2972
rect 257019 2941 257031 2944
rect 256973 2935 257031 2941
rect 244700 2876 252416 2904
rect 244700 2864 244706 2876
rect 226337 2839 226395 2845
rect 226337 2836 226349 2839
rect 223592 2808 226349 2836
rect 226337 2805 226349 2808
rect 226383 2805 226395 2839
rect 226337 2799 226395 2805
rect 244277 2839 244335 2845
rect 244277 2805 244289 2839
rect 244323 2836 244335 2839
rect 245654 2836 245660 2848
rect 244323 2808 245660 2836
rect 244323 2805 244335 2808
rect 244277 2799 244335 2805
rect 245654 2796 245660 2808
rect 245712 2796 245718 2848
rect 246298 2796 246304 2848
rect 246356 2836 246362 2848
rect 255148 2836 255176 2935
rect 255332 2904 255360 2935
rect 258166 2932 258172 2984
rect 258224 2972 258230 2984
rect 259104 2972 259132 3003
rect 260006 3000 260012 3012
rect 260064 3000 260070 3052
rect 260466 3000 260472 3052
rect 260524 3040 260530 3052
rect 261018 3040 261024 3052
rect 260524 3012 261024 3040
rect 260524 3000 260530 3012
rect 261018 3000 261024 3012
rect 261076 3000 261082 3052
rect 261110 3000 261116 3052
rect 261168 3000 261174 3052
rect 261849 3043 261907 3049
rect 261849 3009 261861 3043
rect 261895 3009 261907 3043
rect 261849 3003 261907 3009
rect 267461 3043 267519 3049
rect 267461 3009 267473 3043
rect 267507 3040 267519 3043
rect 267734 3040 267740 3052
rect 267507 3012 267740 3040
rect 267507 3009 267519 3012
rect 267461 3003 267519 3009
rect 258224 2944 259132 2972
rect 258224 2932 258230 2944
rect 260282 2932 260288 2984
rect 260340 2972 260346 2984
rect 260558 2972 260564 2984
rect 260340 2944 260564 2972
rect 260340 2932 260346 2944
rect 260558 2932 260564 2944
rect 260616 2932 260622 2984
rect 260653 2975 260711 2981
rect 260653 2941 260665 2975
rect 260699 2972 260711 2975
rect 261864 2972 261892 3003
rect 267734 3000 267740 3012
rect 267792 3000 267798 3052
rect 268120 3049 268148 3080
rect 268654 3068 268660 3080
rect 268712 3068 268718 3120
rect 268105 3043 268163 3049
rect 268105 3009 268117 3043
rect 268151 3009 268163 3043
rect 268105 3003 268163 3009
rect 268749 3043 268807 3049
rect 268749 3009 268761 3043
rect 268795 3040 268807 3043
rect 269022 3040 269028 3052
rect 268795 3012 269028 3040
rect 268795 3009 268807 3012
rect 268749 3003 268807 3009
rect 269022 3000 269028 3012
rect 269080 3000 269086 3052
rect 269850 3000 269856 3052
rect 269908 3000 269914 3052
rect 270954 3000 270960 3052
rect 271012 3000 271018 3052
rect 260699 2944 261892 2972
rect 266633 2975 266691 2981
rect 260699 2941 260711 2944
rect 260653 2935 260711 2941
rect 266633 2941 266645 2975
rect 266679 2972 266691 2975
rect 268654 2972 268660 2984
rect 266679 2944 268660 2972
rect 266679 2941 266691 2944
rect 266633 2935 266691 2941
rect 268654 2932 268660 2944
rect 268712 2932 268718 2984
rect 258810 2904 258816 2916
rect 255332 2876 258816 2904
rect 258810 2864 258816 2876
rect 258868 2864 258874 2916
rect 260466 2864 260472 2916
rect 260524 2904 260530 2916
rect 262033 2907 262091 2913
rect 262033 2904 262045 2907
rect 260524 2876 262045 2904
rect 260524 2864 260530 2876
rect 262033 2873 262045 2876
rect 262079 2873 262091 2907
rect 262033 2867 262091 2873
rect 266814 2864 266820 2916
rect 266872 2904 266878 2916
rect 267550 2904 267556 2916
rect 266872 2876 267556 2904
rect 266872 2864 266878 2876
rect 267550 2864 267556 2876
rect 267608 2864 267614 2916
rect 246356 2808 255176 2836
rect 246356 2796 246362 2808
rect 258258 2796 258264 2848
rect 258316 2836 258322 2848
rect 259086 2836 259092 2848
rect 258316 2808 259092 2836
rect 258316 2796 258322 2808
rect 259086 2796 259092 2808
rect 259144 2836 259150 2848
rect 259181 2839 259239 2845
rect 259181 2836 259193 2839
rect 259144 2808 259193 2836
rect 259144 2796 259150 2808
rect 259181 2805 259193 2808
rect 259227 2805 259239 2839
rect 259181 2799 259239 2805
rect 259822 2796 259828 2848
rect 259880 2836 259886 2848
rect 261297 2839 261355 2845
rect 261297 2836 261309 2839
rect 259880 2808 261309 2836
rect 259880 2796 259886 2808
rect 261297 2805 261309 2808
rect 261343 2805 261355 2839
rect 261297 2799 261355 2805
rect 266173 2839 266231 2845
rect 266173 2805 266185 2839
rect 266219 2836 266231 2839
rect 267642 2836 267648 2848
rect 266219 2808 267648 2836
rect 266219 2805 266231 2808
rect 266173 2799 266231 2805
rect 267642 2796 267648 2808
rect 267700 2796 267706 2848
rect 267918 2796 267924 2848
rect 267976 2796 267982 2848
rect 270037 2839 270095 2845
rect 270037 2805 270049 2839
rect 270083 2836 270095 2839
rect 270678 2836 270684 2848
rect 270083 2808 270684 2836
rect 270083 2805 270095 2808
rect 270037 2799 270095 2805
rect 270678 2796 270684 2808
rect 270736 2796 270742 2848
rect 1104 2746 271492 2768
rect 1104 2694 34748 2746
rect 34800 2694 34812 2746
rect 34864 2694 34876 2746
rect 34928 2694 34940 2746
rect 34992 2694 35004 2746
rect 35056 2694 102345 2746
rect 102397 2694 102409 2746
rect 102461 2694 102473 2746
rect 102525 2694 102537 2746
rect 102589 2694 102601 2746
rect 102653 2694 169942 2746
rect 169994 2694 170006 2746
rect 170058 2694 170070 2746
rect 170122 2694 170134 2746
rect 170186 2694 170198 2746
rect 170250 2694 237539 2746
rect 237591 2694 237603 2746
rect 237655 2694 237667 2746
rect 237719 2694 237731 2746
rect 237783 2694 237795 2746
rect 237847 2694 271492 2746
rect 1104 2672 271492 2694
rect 842 2592 848 2644
rect 900 2632 906 2644
rect 1765 2635 1823 2641
rect 1765 2632 1777 2635
rect 900 2604 1777 2632
rect 900 2592 906 2604
rect 1765 2601 1777 2604
rect 1811 2601 1823 2635
rect 1765 2595 1823 2601
rect 22005 2635 22063 2641
rect 22005 2601 22017 2635
rect 22051 2632 22063 2635
rect 22830 2632 22836 2644
rect 22051 2604 22836 2632
rect 22051 2601 22063 2604
rect 22005 2595 22063 2601
rect 22830 2592 22836 2604
rect 22888 2592 22894 2644
rect 23658 2592 23664 2644
rect 23716 2632 23722 2644
rect 23753 2635 23811 2641
rect 23753 2632 23765 2635
rect 23716 2604 23765 2632
rect 23716 2592 23722 2604
rect 23753 2601 23765 2604
rect 23799 2601 23811 2635
rect 23753 2595 23811 2601
rect 24581 2635 24639 2641
rect 24581 2601 24593 2635
rect 24627 2632 24639 2635
rect 25038 2632 25044 2644
rect 24627 2604 25044 2632
rect 24627 2601 24639 2604
rect 24581 2595 24639 2601
rect 25038 2592 25044 2604
rect 25096 2592 25102 2644
rect 27614 2592 27620 2644
rect 27672 2592 27678 2644
rect 43530 2592 43536 2644
rect 43588 2592 43594 2644
rect 47486 2592 47492 2644
rect 47544 2632 47550 2644
rect 51810 2632 51816 2644
rect 47544 2604 51816 2632
rect 47544 2592 47550 2604
rect 51810 2592 51816 2604
rect 51868 2592 51874 2644
rect 55214 2592 55220 2644
rect 55272 2632 55278 2644
rect 55677 2635 55735 2641
rect 55677 2632 55689 2635
rect 55272 2604 55689 2632
rect 55272 2592 55278 2604
rect 55677 2601 55689 2604
rect 55723 2601 55735 2635
rect 55677 2595 55735 2601
rect 76699 2635 76757 2641
rect 76699 2601 76711 2635
rect 76745 2632 76757 2635
rect 76745 2604 82124 2632
rect 76745 2601 76757 2604
rect 76699 2595 76757 2601
rect 1854 2524 1860 2576
rect 1912 2564 1918 2576
rect 21266 2564 21272 2576
rect 1912 2536 21272 2564
rect 1912 2524 1918 2536
rect 21266 2524 21272 2536
rect 21324 2524 21330 2576
rect 23474 2564 23480 2576
rect 21376 2536 23480 2564
rect 4798 2456 4804 2508
rect 4856 2456 4862 2508
rect 5534 2456 5540 2508
rect 5592 2496 5598 2508
rect 21376 2496 21404 2536
rect 23474 2524 23480 2536
rect 23532 2524 23538 2576
rect 24302 2524 24308 2576
rect 24360 2564 24366 2576
rect 24762 2564 24768 2576
rect 24360 2536 24768 2564
rect 24360 2524 24366 2536
rect 24762 2524 24768 2536
rect 24820 2564 24826 2576
rect 24949 2567 25007 2573
rect 24949 2564 24961 2567
rect 24820 2536 24961 2564
rect 24820 2524 24826 2536
rect 24949 2533 24961 2536
rect 24995 2564 25007 2567
rect 54294 2564 54300 2576
rect 24995 2536 25360 2564
rect 24995 2533 25007 2536
rect 24949 2527 25007 2533
rect 5592 2468 21404 2496
rect 5592 2456 5598 2468
rect 22462 2456 22468 2508
rect 22520 2496 22526 2508
rect 22557 2499 22615 2505
rect 22557 2496 22569 2499
rect 22520 2468 22569 2496
rect 22520 2456 22526 2468
rect 22557 2465 22569 2468
rect 22603 2465 22615 2499
rect 22557 2459 22615 2465
rect 23382 2456 23388 2508
rect 23440 2456 23446 2508
rect 25332 2505 25360 2536
rect 54036 2536 54300 2564
rect 25317 2499 25375 2505
rect 23584 2468 24624 2496
rect 4522 2388 4528 2440
rect 4580 2388 4586 2440
rect 6730 2388 6736 2440
rect 6788 2388 6794 2440
rect 7006 2388 7012 2440
rect 7064 2388 7070 2440
rect 14826 2388 14832 2440
rect 14884 2388 14890 2440
rect 15102 2388 15108 2440
rect 15160 2388 15166 2440
rect 21821 2431 21879 2437
rect 21821 2397 21833 2431
rect 21867 2428 21879 2431
rect 22094 2428 22100 2440
rect 21867 2400 22100 2428
rect 21867 2397 21879 2400
rect 21821 2391 21879 2397
rect 22094 2388 22100 2400
rect 22152 2388 22158 2440
rect 22278 2388 22284 2440
rect 22336 2428 22342 2440
rect 22741 2431 22799 2437
rect 22741 2428 22753 2431
rect 22336 2400 22753 2428
rect 22336 2388 22342 2400
rect 22741 2397 22753 2400
rect 22787 2428 22799 2431
rect 23290 2428 23296 2440
rect 22787 2400 23296 2428
rect 22787 2397 22799 2400
rect 22741 2391 22799 2397
rect 23290 2388 23296 2400
rect 23348 2428 23354 2440
rect 23584 2437 23612 2468
rect 24596 2440 24624 2468
rect 25317 2465 25329 2499
rect 25363 2465 25375 2499
rect 26050 2496 26056 2508
rect 25317 2459 25375 2465
rect 25424 2468 26056 2496
rect 23569 2431 23627 2437
rect 23569 2428 23581 2431
rect 23348 2400 23581 2428
rect 23348 2388 23354 2400
rect 23569 2397 23581 2400
rect 23615 2397 23627 2431
rect 23569 2391 23627 2397
rect 24394 2388 24400 2440
rect 24452 2388 24458 2440
rect 24578 2388 24584 2440
rect 24636 2428 24642 2440
rect 25424 2428 25452 2468
rect 26050 2456 26056 2468
rect 26108 2496 26114 2508
rect 26421 2499 26479 2505
rect 26421 2496 26433 2499
rect 26108 2468 26433 2496
rect 26108 2456 26114 2468
rect 26421 2465 26433 2468
rect 26467 2465 26479 2499
rect 26421 2459 26479 2465
rect 38470 2456 38476 2508
rect 38528 2456 38534 2508
rect 41322 2496 41328 2508
rect 41262 2482 41328 2496
rect 24636 2400 25452 2428
rect 25501 2431 25559 2437
rect 24636 2388 24642 2400
rect 25501 2397 25513 2431
rect 25547 2428 25559 2431
rect 26145 2431 26203 2437
rect 26145 2428 26157 2431
rect 25547 2400 26157 2428
rect 25547 2397 25559 2400
rect 25501 2391 25559 2397
rect 26145 2397 26157 2400
rect 26191 2428 26203 2431
rect 26326 2428 26332 2440
rect 26191 2400 26332 2428
rect 26191 2397 26203 2400
rect 26145 2391 26203 2397
rect 26326 2388 26332 2400
rect 26384 2388 26390 2440
rect 27430 2388 27436 2440
rect 27488 2388 27494 2440
rect 29730 2388 29736 2440
rect 29788 2388 29794 2440
rect 31938 2388 31944 2440
rect 31996 2388 32002 2440
rect 32033 2431 32091 2437
rect 32033 2397 32045 2431
rect 32079 2397 32091 2431
rect 32033 2391 32091 2397
rect 32048 2360 32076 2391
rect 32766 2388 32772 2440
rect 32824 2388 32830 2440
rect 38194 2388 38200 2440
rect 38252 2428 38258 2440
rect 38381 2431 38439 2437
rect 38381 2428 38393 2431
rect 38252 2400 38393 2428
rect 38252 2388 38258 2400
rect 38381 2397 38393 2400
rect 38427 2397 38439 2431
rect 38488 2428 38516 2456
rect 38841 2431 38899 2437
rect 38488 2400 38792 2428
rect 38381 2391 38439 2397
rect 32490 2360 32496 2372
rect 32048 2332 32496 2360
rect 32490 2320 32496 2332
rect 32548 2360 32554 2372
rect 32953 2363 33011 2369
rect 32953 2360 32965 2363
rect 32548 2332 32965 2360
rect 32548 2320 32554 2332
rect 32953 2329 32965 2332
rect 32999 2329 33011 2363
rect 32953 2323 33011 2329
rect 38010 2320 38016 2372
rect 38068 2360 38074 2372
rect 38470 2360 38476 2372
rect 38068 2332 38476 2360
rect 38068 2320 38074 2332
rect 38470 2320 38476 2332
rect 38528 2320 38534 2372
rect 38764 2360 38792 2400
rect 38841 2397 38853 2431
rect 38887 2428 38899 2431
rect 38930 2428 38936 2440
rect 38887 2400 38936 2428
rect 38887 2397 38899 2400
rect 38841 2391 38899 2397
rect 38930 2388 38936 2400
rect 38988 2388 38994 2440
rect 39132 2428 39160 2482
rect 41248 2468 41328 2482
rect 40126 2428 40132 2440
rect 39132 2400 40132 2428
rect 39132 2360 39160 2400
rect 40126 2388 40132 2400
rect 40184 2388 40190 2440
rect 40494 2388 40500 2440
rect 40552 2388 40558 2440
rect 40954 2388 40960 2440
rect 41012 2388 41018 2440
rect 41046 2388 41052 2440
rect 41104 2428 41110 2440
rect 41248 2428 41276 2468
rect 41322 2456 41328 2468
rect 41380 2456 41386 2508
rect 43990 2496 43996 2508
rect 43286 2468 43996 2496
rect 43990 2456 43996 2468
rect 44048 2456 44054 2508
rect 41104 2400 41276 2428
rect 42521 2431 42579 2437
rect 41104 2388 41110 2400
rect 42521 2397 42533 2431
rect 42567 2428 42579 2431
rect 42886 2428 42892 2440
rect 42567 2400 42892 2428
rect 42567 2397 42579 2400
rect 42521 2391 42579 2397
rect 42886 2388 42892 2400
rect 42944 2388 42950 2440
rect 42978 2388 42984 2440
rect 43036 2388 43042 2440
rect 43346 2428 43352 2440
rect 43272 2400 43352 2428
rect 38764 2332 39160 2360
rect 40586 2320 40592 2372
rect 40644 2320 40650 2372
rect 42613 2363 42671 2369
rect 42613 2329 42625 2363
rect 42659 2360 42671 2363
rect 43272 2360 43300 2400
rect 43346 2388 43352 2400
rect 43404 2388 43410 2440
rect 53745 2431 53803 2437
rect 53745 2397 53757 2431
rect 53791 2428 53803 2431
rect 53834 2428 53840 2440
rect 53791 2400 53840 2428
rect 53791 2397 53803 2400
rect 53745 2391 53803 2397
rect 53834 2388 53840 2400
rect 53892 2428 53898 2440
rect 54036 2437 54064 2536
rect 54294 2524 54300 2536
rect 54352 2564 54358 2576
rect 82096 2564 82124 2604
rect 84930 2592 84936 2644
rect 84988 2632 84994 2644
rect 104250 2632 104256 2644
rect 84988 2604 104256 2632
rect 84988 2592 84994 2604
rect 104250 2592 104256 2604
rect 104308 2592 104314 2644
rect 104342 2592 104348 2644
rect 104400 2632 104406 2644
rect 107562 2632 107568 2644
rect 104400 2604 107568 2632
rect 104400 2592 104406 2604
rect 107562 2592 107568 2604
rect 107620 2592 107626 2644
rect 107654 2592 107660 2644
rect 107712 2632 107718 2644
rect 108666 2632 108672 2644
rect 107712 2604 108672 2632
rect 107712 2592 107718 2604
rect 108666 2592 108672 2604
rect 108724 2592 108730 2644
rect 108758 2592 108764 2644
rect 108816 2632 108822 2644
rect 114738 2632 114744 2644
rect 108816 2604 114744 2632
rect 108816 2592 108822 2604
rect 114738 2592 114744 2604
rect 114796 2592 114802 2644
rect 114848 2604 118280 2632
rect 94682 2564 94688 2576
rect 54352 2536 80054 2564
rect 82096 2536 86954 2564
rect 54352 2524 54358 2536
rect 66162 2456 66168 2508
rect 66220 2496 66226 2508
rect 66809 2499 66867 2505
rect 66809 2496 66821 2499
rect 66220 2468 66821 2496
rect 66220 2456 66226 2468
rect 66809 2465 66821 2468
rect 66855 2465 66867 2499
rect 66809 2459 66867 2465
rect 54021 2431 54079 2437
rect 54021 2428 54033 2431
rect 53892 2400 54033 2428
rect 53892 2388 53898 2400
rect 54021 2397 54033 2400
rect 54067 2397 54079 2431
rect 54021 2391 54079 2397
rect 54202 2388 54208 2440
rect 54260 2388 54266 2440
rect 55490 2388 55496 2440
rect 55548 2388 55554 2440
rect 57514 2388 57520 2440
rect 57572 2428 57578 2440
rect 57793 2431 57851 2437
rect 57793 2428 57805 2431
rect 57572 2400 57805 2428
rect 57572 2388 57578 2400
rect 57793 2397 57805 2400
rect 57839 2397 57851 2431
rect 57793 2391 57851 2397
rect 59170 2388 59176 2440
rect 59228 2428 59234 2440
rect 59265 2431 59323 2437
rect 59265 2428 59277 2431
rect 59228 2400 59277 2428
rect 59228 2388 59234 2400
rect 59265 2397 59277 2400
rect 59311 2397 59323 2431
rect 59265 2391 59323 2397
rect 61473 2431 61531 2437
rect 61473 2397 61485 2431
rect 61519 2428 61531 2431
rect 61654 2428 61660 2440
rect 61519 2400 61660 2428
rect 61519 2397 61531 2400
rect 61473 2391 61531 2397
rect 61654 2388 61660 2400
rect 61712 2388 61718 2440
rect 62206 2388 62212 2440
rect 62264 2388 62270 2440
rect 62666 2388 62672 2440
rect 62724 2428 62730 2440
rect 62945 2431 63003 2437
rect 62945 2428 62957 2431
rect 62724 2400 62957 2428
rect 62724 2388 62730 2400
rect 62945 2397 62957 2400
rect 62991 2397 63003 2431
rect 62945 2391 63003 2397
rect 65426 2388 65432 2440
rect 65484 2428 65490 2440
rect 65797 2431 65855 2437
rect 65797 2428 65809 2431
rect 65484 2400 65809 2428
rect 65484 2388 65490 2400
rect 65797 2397 65809 2400
rect 65843 2397 65855 2431
rect 65797 2391 65855 2397
rect 66533 2431 66591 2437
rect 66533 2397 66545 2431
rect 66579 2428 66591 2431
rect 66714 2428 66720 2440
rect 66579 2400 66720 2428
rect 66579 2397 66591 2400
rect 66533 2391 66591 2397
rect 42659 2332 43300 2360
rect 60737 2363 60795 2369
rect 42659 2329 42671 2332
rect 42613 2323 42671 2329
rect 60737 2329 60749 2363
rect 60783 2360 60795 2363
rect 66548 2360 66576 2391
rect 66714 2388 66720 2400
rect 66772 2388 66778 2440
rect 76466 2388 76472 2440
rect 76524 2388 76530 2440
rect 78674 2388 78680 2440
rect 78732 2388 78738 2440
rect 78950 2388 78956 2440
rect 79008 2388 79014 2440
rect 60783 2332 66576 2360
rect 60783 2329 60795 2332
rect 60737 2323 60795 2329
rect 22186 2252 22192 2304
rect 22244 2292 22250 2304
rect 22925 2295 22983 2301
rect 22925 2292 22937 2295
rect 22244 2264 22937 2292
rect 22244 2252 22250 2264
rect 22925 2261 22937 2264
rect 22971 2261 22983 2295
rect 22925 2255 22983 2261
rect 25685 2295 25743 2301
rect 25685 2261 25697 2295
rect 25731 2292 25743 2295
rect 25866 2292 25872 2304
rect 25731 2264 25872 2292
rect 25731 2261 25743 2264
rect 25685 2255 25743 2261
rect 25866 2252 25872 2264
rect 25924 2252 25930 2304
rect 29914 2252 29920 2304
rect 29972 2252 29978 2304
rect 32217 2295 32275 2301
rect 32217 2261 32229 2295
rect 32263 2292 32275 2295
rect 32674 2292 32680 2304
rect 32263 2264 32680 2292
rect 32263 2261 32275 2264
rect 32217 2255 32275 2261
rect 32674 2252 32680 2264
rect 32732 2252 32738 2304
rect 38105 2295 38163 2301
rect 38105 2261 38117 2295
rect 38151 2292 38163 2295
rect 38286 2292 38292 2304
rect 38151 2264 38292 2292
rect 38151 2261 38163 2264
rect 38105 2255 38163 2261
rect 38286 2252 38292 2264
rect 38344 2252 38350 2304
rect 38378 2252 38384 2304
rect 38436 2292 38442 2304
rect 39209 2295 39267 2301
rect 39209 2292 39221 2295
rect 38436 2264 39221 2292
rect 38436 2252 38442 2264
rect 39209 2261 39221 2264
rect 39255 2261 39267 2295
rect 39209 2255 39267 2261
rect 39393 2295 39451 2301
rect 39393 2261 39405 2295
rect 39439 2292 39451 2295
rect 39850 2292 39856 2304
rect 39439 2264 39856 2292
rect 39439 2261 39451 2264
rect 39393 2255 39451 2261
rect 39850 2252 39856 2264
rect 39908 2252 39914 2304
rect 40218 2252 40224 2304
rect 40276 2252 40282 2304
rect 41322 2252 41328 2304
rect 41380 2252 41386 2304
rect 41506 2252 41512 2304
rect 41564 2252 41570 2304
rect 42242 2252 42248 2304
rect 42300 2252 42306 2304
rect 43346 2252 43352 2304
rect 43404 2252 43410 2304
rect 53742 2252 53748 2304
rect 53800 2292 53806 2304
rect 54389 2295 54447 2301
rect 54389 2292 54401 2295
rect 53800 2264 54401 2292
rect 53800 2252 53806 2264
rect 54389 2261 54401 2264
rect 54435 2261 54447 2295
rect 54389 2255 54447 2261
rect 57974 2252 57980 2304
rect 58032 2252 58038 2304
rect 59354 2252 59360 2304
rect 59412 2292 59418 2304
rect 59449 2295 59507 2301
rect 59449 2292 59461 2295
rect 59412 2264 59461 2292
rect 59412 2252 59418 2264
rect 59449 2261 59461 2264
rect 59495 2261 59507 2295
rect 59449 2255 59507 2261
rect 59814 2252 59820 2304
rect 59872 2292 59878 2304
rect 60829 2295 60887 2301
rect 60829 2292 60841 2295
rect 59872 2264 60841 2292
rect 59872 2252 59878 2264
rect 60829 2261 60841 2264
rect 60875 2261 60887 2295
rect 60829 2255 60887 2261
rect 61470 2252 61476 2304
rect 61528 2292 61534 2304
rect 61657 2295 61715 2301
rect 61657 2292 61669 2295
rect 61528 2264 61669 2292
rect 61528 2252 61534 2264
rect 61657 2261 61669 2264
rect 61703 2261 61715 2295
rect 61657 2255 61715 2261
rect 62390 2252 62396 2304
rect 62448 2252 62454 2304
rect 63126 2252 63132 2304
rect 63184 2252 63190 2304
rect 65978 2252 65984 2304
rect 66036 2252 66042 2304
rect 80026 2292 80054 2536
rect 81897 2499 81955 2505
rect 81897 2465 81909 2499
rect 81943 2496 81955 2499
rect 81943 2468 84056 2496
rect 81943 2465 81955 2468
rect 81897 2459 81955 2465
rect 81618 2388 81624 2440
rect 81676 2388 81682 2440
rect 83826 2388 83832 2440
rect 83884 2388 83890 2440
rect 84028 2428 84056 2468
rect 84102 2456 84108 2508
rect 84160 2456 84166 2508
rect 86926 2496 86954 2536
rect 89824 2536 94688 2564
rect 89824 2496 89852 2536
rect 94682 2524 94688 2536
rect 94740 2524 94746 2576
rect 94774 2524 94780 2576
rect 94832 2564 94838 2576
rect 94961 2567 95019 2573
rect 94961 2564 94973 2567
rect 94832 2536 94973 2564
rect 94832 2524 94838 2536
rect 94961 2533 94973 2536
rect 95007 2533 95019 2567
rect 97626 2564 97632 2576
rect 94961 2527 95019 2533
rect 96632 2536 97632 2564
rect 86926 2468 89852 2496
rect 93854 2456 93860 2508
rect 93912 2496 93918 2508
rect 94317 2499 94375 2505
rect 94317 2496 94329 2499
rect 93912 2468 94329 2496
rect 93912 2456 93918 2468
rect 94317 2465 94329 2468
rect 94363 2465 94375 2499
rect 94317 2459 94375 2465
rect 94501 2499 94559 2505
rect 94501 2465 94513 2499
rect 94547 2496 94559 2499
rect 94590 2496 94596 2508
rect 94547 2468 94596 2496
rect 94547 2465 94559 2468
rect 94501 2459 94559 2465
rect 94590 2456 94596 2468
rect 94648 2456 94654 2508
rect 95234 2456 95240 2508
rect 95292 2456 95298 2508
rect 95375 2499 95433 2505
rect 95375 2465 95387 2499
rect 95421 2496 95433 2499
rect 96632 2496 96660 2536
rect 97626 2524 97632 2536
rect 97684 2524 97690 2576
rect 97718 2524 97724 2576
rect 97776 2564 97782 2576
rect 97776 2536 113588 2564
rect 97776 2524 97782 2536
rect 95421 2468 96660 2496
rect 95421 2465 95433 2468
rect 95375 2459 95433 2465
rect 96706 2456 96712 2508
rect 96764 2496 96770 2508
rect 97353 2499 97411 2505
rect 97353 2496 97365 2499
rect 96764 2468 97365 2496
rect 96764 2456 96770 2468
rect 97353 2465 97365 2468
rect 97399 2465 97411 2499
rect 97353 2459 97411 2465
rect 99650 2456 99656 2508
rect 99708 2456 99714 2508
rect 100018 2456 100024 2508
rect 100076 2496 100082 2508
rect 101953 2499 102011 2505
rect 101953 2496 101965 2499
rect 100076 2468 101965 2496
rect 100076 2456 100082 2468
rect 101953 2465 101965 2468
rect 101999 2465 102011 2499
rect 101953 2459 102011 2465
rect 102134 2456 102140 2508
rect 102192 2456 102198 2508
rect 104802 2456 104808 2508
rect 104860 2456 104866 2508
rect 106182 2456 106188 2508
rect 106240 2456 106246 2508
rect 107194 2456 107200 2508
rect 107252 2456 107258 2508
rect 107654 2456 107660 2508
rect 107712 2456 107718 2508
rect 109034 2496 109040 2508
rect 108408 2468 109040 2496
rect 84930 2428 84936 2440
rect 84028 2400 84936 2428
rect 84930 2388 84936 2400
rect 84988 2388 84994 2440
rect 88518 2388 88524 2440
rect 88576 2428 88582 2440
rect 88889 2431 88947 2437
rect 88889 2428 88901 2431
rect 88576 2400 88901 2428
rect 88576 2388 88582 2400
rect 88889 2397 88901 2400
rect 88935 2428 88947 2431
rect 88978 2428 88984 2440
rect 88935 2400 88984 2428
rect 88935 2397 88947 2400
rect 88889 2391 88947 2397
rect 88978 2388 88984 2400
rect 89036 2388 89042 2440
rect 89070 2388 89076 2440
rect 89128 2388 89134 2440
rect 89993 2431 90051 2437
rect 89993 2397 90005 2431
rect 90039 2428 90051 2431
rect 90266 2428 90272 2440
rect 90039 2400 90272 2428
rect 90039 2397 90051 2400
rect 89993 2391 90051 2397
rect 90266 2388 90272 2400
rect 90324 2388 90330 2440
rect 90729 2431 90787 2437
rect 90729 2397 90741 2431
rect 90775 2428 90787 2431
rect 91094 2428 91100 2440
rect 90775 2400 91100 2428
rect 90775 2397 90787 2400
rect 90729 2391 90787 2397
rect 91094 2388 91100 2400
rect 91152 2388 91158 2440
rect 92198 2388 92204 2440
rect 92256 2388 92262 2440
rect 92842 2388 92848 2440
rect 92900 2388 92906 2440
rect 93581 2431 93639 2437
rect 93581 2397 93593 2431
rect 93627 2428 93639 2431
rect 94406 2428 94412 2440
rect 93627 2400 94412 2428
rect 93627 2397 93639 2400
rect 93581 2391 93639 2397
rect 94406 2388 94412 2400
rect 94464 2388 94470 2440
rect 95510 2388 95516 2440
rect 95568 2388 95574 2440
rect 96157 2431 96215 2437
rect 96157 2397 96169 2431
rect 96203 2428 96215 2431
rect 97169 2431 97227 2437
rect 97169 2428 97181 2431
rect 96203 2400 97181 2428
rect 96203 2397 96215 2400
rect 96157 2391 96215 2397
rect 97169 2397 97181 2400
rect 97215 2397 97227 2431
rect 97169 2391 97227 2397
rect 98730 2388 98736 2440
rect 98788 2428 98794 2440
rect 99469 2431 99527 2437
rect 99469 2428 99481 2431
rect 98788 2400 99481 2428
rect 98788 2388 98794 2400
rect 99469 2397 99481 2400
rect 99515 2397 99527 2431
rect 99469 2391 99527 2397
rect 100938 2388 100944 2440
rect 100996 2428 101002 2440
rect 101306 2428 101312 2440
rect 100996 2400 101312 2428
rect 100996 2388 101002 2400
rect 101306 2388 101312 2400
rect 101364 2388 101370 2440
rect 104621 2431 104679 2437
rect 104621 2428 104633 2431
rect 103348 2400 104633 2428
rect 81158 2320 81164 2372
rect 81216 2360 81222 2372
rect 92290 2360 92296 2372
rect 81216 2332 92296 2360
rect 81216 2320 81222 2332
rect 92290 2320 92296 2332
rect 92348 2320 92354 2372
rect 92385 2363 92443 2369
rect 92385 2329 92397 2363
rect 92431 2360 92443 2363
rect 92566 2360 92572 2372
rect 92431 2332 92572 2360
rect 92431 2329 92443 2332
rect 92385 2323 92443 2329
rect 92566 2320 92572 2332
rect 92624 2320 92630 2372
rect 93044 2332 94544 2360
rect 88518 2292 88524 2304
rect 80026 2264 88524 2292
rect 88518 2252 88524 2264
rect 88576 2252 88582 2304
rect 88794 2252 88800 2304
rect 88852 2292 88858 2304
rect 89257 2295 89315 2301
rect 89257 2292 89269 2295
rect 88852 2264 89269 2292
rect 88852 2252 88858 2264
rect 89257 2261 89269 2264
rect 89303 2261 89315 2295
rect 89257 2255 89315 2261
rect 90174 2252 90180 2304
rect 90232 2252 90238 2304
rect 90913 2295 90971 2301
rect 90913 2261 90925 2295
rect 90959 2292 90971 2295
rect 91186 2292 91192 2304
rect 90959 2264 91192 2292
rect 90959 2261 90971 2264
rect 90913 2255 90971 2261
rect 91186 2252 91192 2264
rect 91244 2252 91250 2304
rect 93044 2301 93072 2332
rect 93029 2295 93087 2301
rect 93029 2261 93041 2295
rect 93075 2261 93087 2295
rect 93029 2255 93087 2261
rect 93762 2252 93768 2304
rect 93820 2252 93826 2304
rect 94516 2292 94544 2332
rect 96062 2320 96068 2372
rect 96120 2360 96126 2372
rect 97902 2360 97908 2372
rect 96120 2332 97908 2360
rect 96120 2320 96126 2332
rect 97902 2320 97908 2332
rect 97960 2320 97966 2372
rect 99006 2320 99012 2372
rect 99064 2360 99070 2372
rect 100478 2360 100484 2372
rect 99064 2332 100484 2360
rect 99064 2320 99070 2332
rect 100478 2320 100484 2332
rect 100536 2320 100542 2372
rect 101490 2320 101496 2372
rect 101548 2360 101554 2372
rect 103348 2360 103376 2400
rect 104621 2397 104633 2400
rect 104667 2397 104679 2431
rect 104621 2391 104679 2397
rect 107013 2431 107071 2437
rect 107013 2397 107025 2431
rect 107059 2397 107071 2431
rect 107013 2391 107071 2397
rect 101548 2332 103376 2360
rect 103793 2363 103851 2369
rect 101548 2320 101554 2332
rect 103793 2329 103805 2363
rect 103839 2360 103851 2363
rect 106366 2360 106372 2372
rect 103839 2332 106372 2360
rect 103839 2329 103851 2332
rect 103793 2323 103851 2329
rect 106366 2320 106372 2332
rect 106424 2320 106430 2372
rect 107028 2360 107056 2391
rect 108408 2360 108436 2468
rect 109034 2456 109040 2468
rect 109092 2456 109098 2508
rect 109494 2456 109500 2508
rect 109552 2456 109558 2508
rect 111153 2499 111211 2505
rect 111153 2465 111165 2499
rect 111199 2496 111211 2499
rect 112625 2499 112683 2505
rect 112625 2496 112637 2499
rect 111199 2468 112637 2496
rect 111199 2465 111211 2468
rect 111153 2459 111211 2465
rect 112625 2465 112637 2468
rect 112671 2496 112683 2499
rect 113358 2496 113364 2508
rect 112671 2468 113364 2496
rect 112671 2465 112683 2468
rect 112625 2459 112683 2465
rect 113358 2456 113364 2468
rect 113416 2456 113422 2508
rect 108482 2388 108488 2440
rect 108540 2428 108546 2440
rect 109313 2431 109371 2437
rect 109313 2428 109325 2431
rect 108540 2400 109325 2428
rect 108540 2388 108546 2400
rect 109313 2397 109325 2400
rect 109359 2397 109371 2431
rect 109313 2391 109371 2397
rect 110690 2388 110696 2440
rect 110748 2428 110754 2440
rect 112070 2428 112076 2440
rect 110748 2400 112076 2428
rect 110748 2388 110754 2400
rect 112070 2388 112076 2400
rect 112128 2388 112134 2440
rect 112162 2388 112168 2440
rect 112220 2388 112226 2440
rect 113560 2428 113588 2536
rect 114554 2524 114560 2576
rect 114612 2564 114618 2576
rect 114848 2564 114876 2604
rect 114612 2536 114876 2564
rect 114612 2524 114618 2536
rect 117314 2524 117320 2576
rect 117372 2564 117378 2576
rect 117372 2536 118188 2564
rect 117372 2524 117378 2536
rect 113818 2456 113824 2508
rect 113876 2496 113882 2508
rect 115017 2499 115075 2505
rect 115017 2496 115029 2499
rect 113876 2468 115029 2496
rect 113876 2456 113882 2468
rect 115017 2465 115029 2468
rect 115063 2465 115075 2499
rect 115017 2459 115075 2465
rect 114833 2431 114891 2437
rect 114833 2428 114845 2431
rect 113560 2400 114845 2428
rect 114833 2397 114845 2400
rect 114879 2397 114891 2431
rect 117222 2428 117228 2440
rect 114833 2391 114891 2397
rect 116596 2400 117228 2428
rect 107028 2332 108436 2360
rect 108500 2332 111104 2360
rect 96246 2292 96252 2304
rect 94516 2264 96252 2292
rect 96246 2252 96252 2264
rect 96304 2252 96310 2304
rect 96430 2252 96436 2304
rect 96488 2292 96494 2304
rect 98822 2292 98828 2304
rect 96488 2264 98828 2292
rect 96488 2252 96494 2264
rect 98822 2252 98828 2264
rect 98880 2252 98886 2304
rect 99098 2252 99104 2304
rect 99156 2292 99162 2304
rect 104894 2292 104900 2304
rect 99156 2264 104900 2292
rect 99156 2252 99162 2264
rect 104894 2252 104900 2264
rect 104952 2252 104958 2304
rect 107838 2252 107844 2304
rect 107896 2292 107902 2304
rect 108500 2292 108528 2332
rect 107896 2264 108528 2292
rect 107896 2252 107902 2264
rect 108574 2252 108580 2304
rect 108632 2292 108638 2304
rect 110230 2292 110236 2304
rect 108632 2264 110236 2292
rect 108632 2252 108638 2264
rect 110230 2252 110236 2264
rect 110288 2252 110294 2304
rect 111076 2292 111104 2332
rect 112346 2320 112352 2372
rect 112404 2320 112410 2372
rect 116596 2360 116624 2400
rect 117222 2388 117228 2400
rect 117280 2388 117286 2440
rect 117314 2388 117320 2440
rect 117372 2428 117378 2440
rect 118160 2437 118188 2536
rect 117501 2431 117559 2437
rect 117501 2428 117513 2431
rect 117372 2400 117513 2428
rect 117372 2388 117378 2400
rect 117501 2397 117513 2400
rect 117547 2397 117559 2431
rect 117501 2391 117559 2397
rect 118145 2431 118203 2437
rect 118145 2397 118157 2431
rect 118191 2397 118203 2431
rect 118252 2428 118280 2604
rect 124214 2592 124220 2644
rect 124272 2592 124278 2644
rect 133874 2592 133880 2644
rect 133932 2632 133938 2644
rect 133969 2635 134027 2641
rect 133969 2632 133981 2635
rect 133932 2604 133981 2632
rect 133932 2592 133938 2604
rect 133969 2601 133981 2604
rect 134015 2601 134027 2635
rect 133969 2595 134027 2601
rect 138661 2635 138719 2641
rect 138661 2601 138673 2635
rect 138707 2632 138719 2635
rect 139946 2632 139952 2644
rect 138707 2604 139952 2632
rect 138707 2601 138719 2604
rect 138661 2595 138719 2601
rect 139946 2592 139952 2604
rect 140004 2592 140010 2644
rect 140958 2632 140964 2644
rect 140056 2604 140964 2632
rect 138934 2524 138940 2576
rect 138992 2564 138998 2576
rect 140056 2564 140084 2604
rect 140958 2592 140964 2604
rect 141016 2592 141022 2644
rect 141142 2592 141148 2644
rect 141200 2592 141206 2644
rect 141973 2635 142031 2641
rect 141973 2601 141985 2635
rect 142019 2632 142031 2635
rect 142246 2632 142252 2644
rect 142019 2604 142252 2632
rect 142019 2601 142031 2604
rect 141973 2595 142031 2601
rect 142246 2592 142252 2604
rect 142304 2592 142310 2644
rect 142430 2592 142436 2644
rect 142488 2632 142494 2644
rect 146662 2632 146668 2644
rect 142488 2604 146668 2632
rect 142488 2592 142494 2604
rect 146662 2592 146668 2604
rect 146720 2592 146726 2644
rect 153010 2632 153016 2644
rect 147646 2604 153016 2632
rect 138992 2536 140084 2564
rect 138992 2524 138998 2536
rect 141786 2524 141792 2576
rect 141844 2564 141850 2576
rect 147646 2564 147674 2604
rect 153010 2592 153016 2604
rect 153068 2592 153074 2644
rect 153381 2635 153439 2641
rect 153381 2601 153393 2635
rect 153427 2632 153439 2635
rect 153746 2632 153752 2644
rect 153427 2604 153752 2632
rect 153427 2601 153439 2604
rect 153381 2595 153439 2601
rect 153746 2592 153752 2604
rect 153804 2592 153810 2644
rect 154669 2635 154727 2641
rect 154669 2601 154681 2635
rect 154715 2632 154727 2635
rect 155218 2632 155224 2644
rect 154715 2604 155224 2632
rect 154715 2601 154727 2604
rect 154669 2595 154727 2601
rect 155218 2592 155224 2604
rect 155276 2592 155282 2644
rect 155773 2635 155831 2641
rect 155773 2601 155785 2635
rect 155819 2632 155831 2635
rect 156414 2632 156420 2644
rect 155819 2604 156420 2632
rect 155819 2601 155831 2604
rect 155773 2595 155831 2601
rect 156414 2592 156420 2604
rect 156472 2592 156478 2644
rect 157306 2604 185072 2632
rect 141844 2536 147674 2564
rect 141844 2524 141850 2536
rect 149054 2524 149060 2576
rect 149112 2564 149118 2576
rect 152734 2564 152740 2576
rect 149112 2536 152740 2564
rect 149112 2524 149118 2536
rect 152734 2524 152740 2536
rect 152792 2524 152798 2576
rect 152918 2524 152924 2576
rect 152976 2564 152982 2576
rect 152976 2536 153608 2564
rect 152976 2524 152982 2536
rect 118694 2456 118700 2508
rect 118752 2496 118758 2508
rect 119709 2499 119767 2505
rect 119709 2496 119721 2499
rect 118752 2468 119721 2496
rect 118752 2456 118758 2468
rect 119709 2465 119721 2468
rect 119755 2465 119767 2499
rect 119709 2459 119767 2465
rect 120258 2456 120264 2508
rect 120316 2456 120322 2508
rect 121914 2496 121920 2508
rect 121104 2468 121920 2496
rect 118789 2431 118847 2437
rect 118789 2428 118801 2431
rect 118252 2400 118801 2428
rect 118145 2391 118203 2397
rect 118789 2397 118801 2400
rect 118835 2397 118847 2431
rect 118789 2391 118847 2397
rect 118970 2388 118976 2440
rect 119028 2428 119034 2440
rect 119525 2431 119583 2437
rect 119525 2428 119537 2431
rect 119028 2400 119537 2428
rect 119028 2388 119034 2400
rect 119525 2397 119537 2400
rect 119571 2397 119583 2431
rect 119525 2391 119583 2397
rect 115032 2332 116624 2360
rect 116673 2363 116731 2369
rect 115032 2304 115060 2332
rect 116673 2329 116685 2363
rect 116719 2360 116731 2363
rect 121104 2360 121132 2468
rect 121914 2456 121920 2468
rect 121972 2456 121978 2508
rect 124766 2456 124772 2508
rect 124824 2456 124830 2508
rect 129737 2499 129795 2505
rect 129737 2465 129749 2499
rect 129783 2496 129795 2499
rect 130194 2496 130200 2508
rect 129783 2468 130200 2496
rect 129783 2465 129795 2468
rect 129737 2459 129795 2465
rect 130194 2456 130200 2468
rect 130252 2456 130258 2508
rect 134613 2499 134671 2505
rect 134613 2465 134625 2499
rect 134659 2496 134671 2499
rect 135346 2496 135352 2508
rect 134659 2468 135352 2496
rect 134659 2465 134671 2468
rect 134613 2459 134671 2465
rect 135346 2456 135352 2468
rect 135404 2456 135410 2508
rect 139302 2456 139308 2508
rect 139360 2456 139366 2508
rect 139946 2456 139952 2508
rect 140004 2456 140010 2508
rect 140682 2496 140688 2508
rect 140516 2468 140688 2496
rect 121178 2388 121184 2440
rect 121236 2428 121242 2440
rect 122561 2431 122619 2437
rect 122561 2428 122573 2431
rect 121236 2400 122573 2428
rect 121236 2388 121242 2400
rect 122561 2397 122573 2400
rect 122607 2428 122619 2431
rect 124033 2431 124091 2437
rect 122607 2400 122834 2428
rect 122607 2397 122619 2400
rect 122561 2391 122619 2397
rect 116719 2332 121132 2360
rect 122806 2360 122834 2400
rect 124033 2397 124045 2431
rect 124079 2428 124091 2431
rect 124306 2428 124312 2440
rect 124079 2400 124312 2428
rect 124079 2397 124091 2400
rect 124033 2391 124091 2397
rect 124306 2388 124312 2400
rect 124364 2388 124370 2440
rect 124950 2388 124956 2440
rect 125008 2388 125014 2440
rect 126054 2388 126060 2440
rect 126112 2388 126118 2440
rect 126698 2388 126704 2440
rect 126756 2428 126762 2440
rect 126793 2431 126851 2437
rect 126793 2428 126805 2431
rect 126756 2400 126805 2428
rect 126756 2388 126762 2400
rect 126793 2397 126805 2400
rect 126839 2397 126851 2431
rect 126793 2391 126851 2397
rect 128265 2431 128323 2437
rect 128265 2397 128277 2431
rect 128311 2428 128323 2431
rect 128354 2428 128360 2440
rect 128311 2400 128360 2428
rect 128311 2397 128323 2400
rect 128265 2391 128323 2397
rect 128354 2388 128360 2400
rect 128412 2388 128418 2440
rect 128998 2388 129004 2440
rect 129056 2388 129062 2440
rect 129642 2388 129648 2440
rect 129700 2428 129706 2440
rect 129921 2431 129979 2437
rect 129921 2428 129933 2431
rect 129700 2400 129933 2428
rect 129700 2388 129706 2400
rect 129921 2397 129933 2400
rect 129967 2397 129979 2431
rect 129921 2391 129979 2397
rect 130105 2431 130163 2437
rect 130105 2397 130117 2431
rect 130151 2428 130163 2431
rect 130565 2431 130623 2437
rect 130565 2428 130577 2431
rect 130151 2400 130577 2428
rect 130151 2397 130163 2400
rect 130105 2391 130163 2397
rect 130565 2397 130577 2400
rect 130611 2397 130623 2431
rect 130565 2391 130623 2397
rect 131485 2431 131543 2437
rect 131485 2397 131497 2431
rect 131531 2428 131543 2431
rect 131758 2428 131764 2440
rect 131531 2400 131764 2428
rect 131531 2397 131543 2400
rect 131485 2391 131543 2397
rect 131758 2388 131764 2400
rect 131816 2388 131822 2440
rect 133049 2431 133107 2437
rect 133049 2397 133061 2431
rect 133095 2428 133107 2431
rect 133506 2428 133512 2440
rect 133095 2400 133512 2428
rect 133095 2397 133107 2400
rect 133049 2391 133107 2397
rect 133506 2388 133512 2400
rect 133564 2388 133570 2440
rect 133690 2388 133696 2440
rect 133748 2428 133754 2440
rect 133785 2431 133843 2437
rect 133785 2428 133797 2431
rect 133748 2400 133797 2428
rect 133748 2388 133754 2400
rect 133785 2397 133797 2400
rect 133831 2397 133843 2431
rect 133785 2391 133843 2397
rect 134334 2388 134340 2440
rect 134392 2428 134398 2440
rect 134797 2431 134855 2437
rect 134797 2428 134809 2431
rect 134392 2400 134809 2428
rect 134392 2388 134398 2400
rect 134797 2397 134809 2400
rect 134843 2397 134855 2431
rect 134797 2391 134855 2397
rect 138845 2431 138903 2437
rect 138845 2397 138857 2431
rect 138891 2397 138903 2431
rect 138845 2391 138903 2397
rect 128814 2360 128820 2372
rect 122806 2332 128820 2360
rect 116719 2329 116731 2332
rect 116673 2323 116731 2329
rect 128814 2320 128820 2332
rect 128872 2320 128878 2372
rect 115014 2292 115020 2304
rect 111076 2264 115020 2292
rect 115014 2252 115020 2264
rect 115072 2252 115078 2304
rect 116026 2252 116032 2304
rect 116084 2292 116090 2304
rect 117317 2295 117375 2301
rect 117317 2292 117329 2295
rect 116084 2264 117329 2292
rect 116084 2252 116090 2264
rect 117317 2261 117329 2264
rect 117363 2261 117375 2295
rect 117317 2255 117375 2261
rect 117590 2252 117596 2304
rect 117648 2292 117654 2304
rect 117961 2295 118019 2301
rect 117961 2292 117973 2295
rect 117648 2264 117973 2292
rect 117648 2252 117654 2264
rect 117961 2261 117973 2264
rect 118007 2261 118019 2295
rect 117961 2255 118019 2261
rect 118050 2252 118056 2304
rect 118108 2292 118114 2304
rect 118605 2295 118663 2301
rect 118605 2292 118617 2295
rect 118108 2264 118617 2292
rect 118108 2252 118114 2264
rect 118605 2261 118617 2264
rect 118651 2261 118663 2295
rect 118605 2255 118663 2261
rect 122650 2252 122656 2304
rect 122708 2252 122714 2304
rect 125134 2252 125140 2304
rect 125192 2252 125198 2304
rect 126238 2252 126244 2304
rect 126296 2252 126302 2304
rect 126974 2252 126980 2304
rect 127032 2252 127038 2304
rect 128446 2252 128452 2304
rect 128504 2252 128510 2304
rect 129182 2252 129188 2304
rect 129240 2252 129246 2304
rect 130746 2252 130752 2304
rect 130804 2252 130810 2304
rect 131666 2252 131672 2304
rect 131724 2252 131730 2304
rect 133230 2252 133236 2304
rect 133288 2252 133294 2304
rect 134981 2295 135039 2301
rect 134981 2261 134993 2295
rect 135027 2292 135039 2295
rect 135346 2292 135352 2304
rect 135027 2264 135352 2292
rect 135027 2261 135039 2264
rect 134981 2255 135039 2261
rect 135346 2252 135352 2264
rect 135404 2252 135410 2304
rect 138860 2292 138888 2391
rect 139486 2388 139492 2440
rect 139544 2388 139550 2440
rect 140222 2388 140228 2440
rect 140280 2388 140286 2440
rect 140314 2388 140320 2440
rect 140372 2437 140378 2440
rect 140516 2437 140544 2468
rect 140682 2456 140688 2468
rect 140740 2456 140746 2508
rect 143350 2456 143356 2508
rect 143408 2496 143414 2508
rect 145561 2499 145619 2505
rect 145561 2496 145573 2499
rect 143408 2468 145573 2496
rect 143408 2456 143414 2468
rect 145561 2465 145573 2468
rect 145607 2465 145619 2499
rect 145561 2459 145619 2465
rect 146294 2456 146300 2508
rect 146352 2456 146358 2508
rect 148594 2456 148600 2508
rect 148652 2456 148658 2508
rect 148778 2456 148784 2508
rect 148836 2456 148842 2508
rect 150250 2456 150256 2508
rect 150308 2456 150314 2508
rect 150802 2456 150808 2508
rect 150860 2496 150866 2508
rect 151081 2499 151139 2505
rect 151081 2496 151093 2499
rect 150860 2468 151093 2496
rect 150860 2456 150866 2468
rect 151081 2465 151093 2468
rect 151127 2465 151139 2499
rect 151081 2459 151139 2465
rect 151354 2456 151360 2508
rect 151412 2456 151418 2508
rect 151814 2456 151820 2508
rect 151872 2496 151878 2508
rect 153580 2496 153608 2536
rect 154482 2524 154488 2576
rect 154540 2564 154546 2576
rect 157306 2564 157334 2604
rect 154540 2536 157334 2564
rect 154540 2524 154546 2536
rect 158438 2524 158444 2576
rect 158496 2564 158502 2576
rect 166534 2564 166540 2576
rect 158496 2536 166540 2564
rect 158496 2524 158502 2536
rect 166534 2524 166540 2536
rect 166592 2524 166598 2576
rect 168374 2524 168380 2576
rect 168432 2564 168438 2576
rect 168432 2536 184888 2564
rect 168432 2524 168438 2536
rect 182085 2499 182143 2505
rect 182085 2496 182097 2499
rect 151872 2468 153516 2496
rect 153580 2468 182097 2496
rect 151872 2456 151878 2468
rect 140372 2431 140400 2437
rect 140388 2397 140400 2431
rect 140372 2391 140400 2397
rect 140501 2431 140559 2437
rect 140501 2397 140513 2431
rect 140547 2397 140559 2431
rect 140501 2391 140559 2397
rect 140372 2388 140378 2391
rect 141602 2388 141608 2440
rect 141660 2388 141666 2440
rect 141970 2388 141976 2440
rect 142028 2388 142034 2440
rect 142154 2388 142160 2440
rect 142212 2428 142218 2440
rect 143077 2431 143135 2437
rect 143077 2428 143089 2431
rect 142212 2400 143089 2428
rect 142212 2388 142218 2400
rect 143077 2397 143089 2400
rect 143123 2397 143135 2431
rect 143077 2391 143135 2397
rect 145374 2388 145380 2440
rect 145432 2388 145438 2440
rect 147646 2400 148364 2428
rect 141234 2320 141240 2372
rect 141292 2360 141298 2372
rect 143261 2363 143319 2369
rect 143261 2360 143273 2363
rect 141292 2332 143273 2360
rect 141292 2320 141298 2332
rect 143261 2329 143273 2332
rect 143307 2329 143319 2363
rect 143261 2323 143319 2329
rect 144730 2320 144736 2372
rect 144788 2360 144794 2372
rect 144917 2363 144975 2369
rect 144917 2360 144929 2363
rect 144788 2332 144929 2360
rect 144788 2320 144794 2332
rect 144917 2329 144929 2332
rect 144963 2329 144975 2363
rect 144917 2323 144975 2329
rect 146386 2320 146392 2372
rect 146444 2360 146450 2372
rect 147646 2360 147674 2400
rect 146444 2332 147674 2360
rect 148336 2360 148364 2400
rect 150894 2388 150900 2440
rect 150952 2388 150958 2440
rect 153378 2428 153384 2440
rect 152292 2400 153384 2428
rect 148502 2360 148508 2372
rect 148336 2332 148508 2360
rect 146444 2320 146450 2332
rect 148502 2320 148508 2332
rect 148560 2320 148566 2372
rect 150434 2320 150440 2372
rect 150492 2360 150498 2372
rect 152292 2360 152320 2400
rect 153378 2388 153384 2400
rect 153436 2388 153442 2440
rect 153488 2428 153516 2468
rect 182085 2465 182097 2468
rect 182131 2465 182143 2499
rect 182085 2459 182143 2465
rect 153565 2431 153623 2437
rect 153565 2428 153577 2431
rect 153488 2400 153577 2428
rect 153565 2397 153577 2400
rect 153611 2397 153623 2431
rect 153565 2391 153623 2397
rect 154114 2388 154120 2440
rect 154172 2428 154178 2440
rect 154209 2431 154267 2437
rect 154209 2428 154221 2431
rect 154172 2400 154221 2428
rect 154172 2388 154178 2400
rect 154209 2397 154221 2400
rect 154255 2397 154267 2431
rect 154209 2391 154267 2397
rect 154482 2388 154488 2440
rect 154540 2428 154546 2440
rect 154853 2431 154911 2437
rect 154853 2428 154865 2431
rect 154540 2400 154865 2428
rect 154540 2388 154546 2400
rect 154853 2397 154865 2400
rect 154899 2397 154911 2431
rect 154853 2391 154911 2397
rect 155586 2388 155592 2440
rect 155644 2388 155650 2440
rect 156233 2431 156291 2437
rect 156233 2397 156245 2431
rect 156279 2428 156291 2431
rect 156598 2428 156604 2440
rect 156279 2400 156604 2428
rect 156279 2397 156291 2400
rect 156233 2391 156291 2397
rect 156598 2388 156604 2400
rect 156656 2388 156662 2440
rect 156966 2388 156972 2440
rect 157024 2428 157030 2440
rect 157024 2400 157334 2428
rect 157024 2388 157030 2400
rect 150492 2332 152320 2360
rect 150492 2320 150498 2332
rect 156414 2320 156420 2372
rect 156472 2360 156478 2372
rect 156690 2360 156696 2372
rect 156472 2332 156696 2360
rect 156472 2320 156478 2332
rect 156690 2320 156696 2332
rect 156748 2360 156754 2372
rect 157061 2363 157119 2369
rect 157061 2360 157073 2363
rect 156748 2332 157073 2360
rect 156748 2320 156754 2332
rect 157061 2329 157073 2332
rect 157107 2329 157119 2363
rect 157306 2360 157334 2400
rect 157702 2388 157708 2440
rect 157760 2388 157766 2440
rect 158438 2388 158444 2440
rect 158496 2428 158502 2440
rect 158625 2431 158683 2437
rect 158625 2428 158637 2431
rect 158496 2400 158637 2428
rect 158496 2388 158502 2400
rect 158625 2397 158637 2400
rect 158671 2397 158683 2431
rect 158625 2391 158683 2397
rect 159910 2388 159916 2440
rect 159968 2388 159974 2440
rect 160002 2388 160008 2440
rect 160060 2388 160066 2440
rect 160189 2431 160247 2437
rect 160189 2397 160201 2431
rect 160235 2428 160247 2431
rect 160649 2431 160707 2437
rect 160649 2428 160661 2431
rect 160235 2400 160661 2428
rect 160235 2397 160247 2400
rect 160189 2391 160247 2397
rect 160649 2397 160661 2400
rect 160695 2397 160707 2431
rect 160649 2391 160707 2397
rect 161474 2388 161480 2440
rect 161532 2388 161538 2440
rect 163685 2431 163743 2437
rect 163685 2397 163697 2431
rect 163731 2428 163743 2431
rect 163958 2428 163964 2440
rect 163731 2400 163964 2428
rect 163731 2397 163743 2400
rect 163685 2391 163743 2397
rect 163958 2388 163964 2400
rect 164016 2388 164022 2440
rect 165065 2431 165123 2437
rect 165065 2397 165077 2431
rect 165111 2428 165123 2431
rect 165614 2428 165620 2440
rect 165111 2400 165620 2428
rect 165111 2397 165123 2400
rect 165065 2391 165123 2397
rect 165614 2388 165620 2400
rect 165672 2388 165678 2440
rect 165798 2388 165804 2440
rect 165856 2388 165862 2440
rect 166629 2431 166687 2437
rect 166629 2397 166641 2431
rect 166675 2428 166687 2431
rect 167454 2428 167460 2440
rect 166675 2400 167460 2428
rect 166675 2397 166687 2400
rect 166629 2391 166687 2397
rect 167454 2388 167460 2400
rect 167512 2388 167518 2440
rect 167914 2388 167920 2440
rect 167972 2388 167978 2440
rect 168006 2388 168012 2440
rect 168064 2428 168070 2440
rect 168282 2428 168288 2440
rect 168064 2400 168288 2428
rect 168064 2388 168070 2400
rect 168282 2388 168288 2400
rect 168340 2388 168346 2440
rect 168837 2431 168895 2437
rect 168837 2430 168849 2431
rect 168760 2428 168849 2430
rect 168392 2402 168849 2428
rect 168392 2400 168788 2402
rect 158990 2360 158996 2372
rect 157306 2332 158996 2360
rect 157061 2323 157119 2329
rect 158990 2320 158996 2332
rect 159048 2320 159054 2372
rect 162305 2363 162363 2369
rect 162305 2329 162317 2363
rect 162351 2360 162363 2363
rect 167730 2360 167736 2372
rect 162351 2332 167736 2360
rect 162351 2329 162363 2332
rect 162305 2323 162363 2329
rect 167730 2320 167736 2332
rect 167788 2360 167794 2372
rect 168392 2360 168420 2400
rect 168837 2397 168849 2402
rect 168883 2397 168895 2431
rect 169113 2431 169171 2437
rect 169113 2428 169125 2431
rect 168837 2391 168895 2397
rect 168944 2400 169125 2428
rect 167788 2332 168420 2360
rect 167788 2320 167794 2332
rect 140774 2292 140780 2304
rect 138860 2264 140780 2292
rect 140774 2252 140780 2264
rect 140832 2252 140838 2304
rect 140958 2252 140964 2304
rect 141016 2292 141022 2304
rect 142157 2295 142215 2301
rect 142157 2292 142169 2295
rect 141016 2264 142169 2292
rect 141016 2252 141022 2264
rect 142157 2261 142169 2264
rect 142203 2261 142215 2295
rect 142157 2255 142215 2261
rect 144270 2252 144276 2304
rect 144328 2292 144334 2304
rect 146846 2292 146852 2304
rect 144328 2264 146852 2292
rect 144328 2252 144334 2264
rect 146846 2252 146852 2264
rect 146904 2252 146910 2304
rect 148318 2252 148324 2304
rect 148376 2292 148382 2304
rect 151078 2292 151084 2304
rect 148376 2264 151084 2292
rect 148376 2252 148382 2264
rect 151078 2252 151084 2264
rect 151136 2292 151142 2304
rect 151446 2292 151452 2304
rect 151136 2264 151452 2292
rect 151136 2252 151142 2264
rect 151446 2252 151452 2264
rect 151504 2252 151510 2304
rect 153470 2252 153476 2304
rect 153528 2292 153534 2304
rect 154025 2295 154083 2301
rect 154025 2292 154037 2295
rect 153528 2264 154037 2292
rect 153528 2252 153534 2264
rect 154025 2261 154037 2264
rect 154071 2261 154083 2295
rect 154025 2255 154083 2261
rect 157242 2252 157248 2304
rect 157300 2292 157306 2304
rect 157889 2295 157947 2301
rect 157889 2292 157901 2295
rect 157300 2264 157901 2292
rect 157300 2252 157306 2264
rect 157889 2261 157901 2264
rect 157935 2261 157947 2295
rect 157889 2255 157947 2261
rect 160830 2252 160836 2304
rect 160888 2252 160894 2304
rect 161658 2252 161664 2304
rect 161716 2252 161722 2304
rect 162394 2252 162400 2304
rect 162452 2252 162458 2304
rect 163866 2252 163872 2304
rect 163924 2252 163930 2304
rect 165246 2252 165252 2304
rect 165304 2252 165310 2304
rect 165982 2252 165988 2304
rect 166040 2252 166046 2304
rect 166810 2252 166816 2304
rect 166868 2252 166874 2304
rect 168190 2252 168196 2304
rect 168248 2252 168254 2304
rect 168282 2252 168288 2304
rect 168340 2292 168346 2304
rect 168944 2292 168972 2400
rect 169113 2397 169125 2400
rect 169159 2397 169171 2431
rect 169113 2391 169171 2397
rect 176654 2388 176660 2440
rect 176712 2388 176718 2440
rect 176930 2388 176936 2440
rect 176988 2388 176994 2440
rect 179598 2388 179604 2440
rect 179656 2388 179662 2440
rect 179877 2431 179935 2437
rect 179877 2397 179889 2431
rect 179923 2397 179935 2431
rect 179877 2391 179935 2397
rect 172422 2320 172428 2372
rect 172480 2360 172486 2372
rect 179892 2360 179920 2391
rect 181806 2388 181812 2440
rect 181864 2388 181870 2440
rect 184750 2388 184756 2440
rect 184808 2388 184814 2440
rect 184860 2428 184888 2536
rect 185044 2505 185072 2604
rect 190454 2592 190460 2644
rect 190512 2632 190518 2644
rect 190549 2635 190607 2641
rect 190549 2632 190561 2635
rect 190512 2604 190561 2632
rect 190512 2592 190518 2604
rect 190549 2601 190561 2604
rect 190595 2601 190607 2635
rect 190549 2595 190607 2601
rect 191834 2592 191840 2644
rect 191892 2632 191898 2644
rect 192021 2635 192079 2641
rect 192021 2632 192033 2635
rect 191892 2604 192033 2632
rect 191892 2592 191898 2604
rect 192021 2601 192033 2604
rect 192067 2601 192079 2635
rect 192021 2595 192079 2601
rect 198734 2592 198740 2644
rect 198792 2592 198798 2644
rect 217594 2632 217600 2644
rect 200086 2604 217600 2632
rect 192386 2524 192392 2576
rect 192444 2564 192450 2576
rect 192846 2564 192852 2576
rect 192444 2536 192852 2564
rect 192444 2524 192450 2536
rect 192846 2524 192852 2536
rect 192904 2564 192910 2576
rect 200086 2564 200114 2604
rect 217594 2592 217600 2604
rect 217652 2592 217658 2644
rect 217796 2604 219112 2632
rect 192904 2536 200114 2564
rect 192904 2524 192910 2536
rect 200206 2524 200212 2576
rect 200264 2564 200270 2576
rect 200393 2567 200451 2573
rect 200393 2564 200405 2567
rect 200264 2536 200405 2564
rect 200264 2524 200270 2536
rect 200393 2533 200405 2536
rect 200439 2533 200451 2567
rect 200393 2527 200451 2533
rect 201494 2524 201500 2576
rect 201552 2564 201558 2576
rect 201957 2567 202015 2573
rect 201957 2564 201969 2567
rect 201552 2536 201969 2564
rect 201552 2524 201558 2536
rect 201957 2533 201969 2536
rect 202003 2533 202015 2567
rect 217796 2564 217824 2604
rect 201957 2527 202015 2533
rect 207584 2536 217824 2564
rect 185029 2499 185087 2505
rect 185029 2465 185041 2499
rect 185075 2465 185087 2499
rect 187237 2499 187295 2505
rect 187237 2496 187249 2499
rect 185029 2459 185087 2465
rect 185136 2468 187249 2496
rect 185136 2428 185164 2468
rect 187237 2465 187249 2468
rect 187283 2465 187295 2499
rect 187237 2459 187295 2465
rect 202782 2456 202788 2508
rect 202840 2496 202846 2508
rect 202840 2468 203288 2496
rect 202840 2456 202846 2468
rect 184860 2400 185164 2428
rect 186958 2388 186964 2440
rect 187016 2388 187022 2440
rect 190365 2431 190423 2437
rect 190365 2397 190377 2431
rect 190411 2428 190423 2431
rect 190914 2428 190920 2440
rect 190411 2400 190920 2428
rect 190411 2397 190423 2400
rect 190365 2391 190423 2397
rect 190914 2388 190920 2400
rect 190972 2388 190978 2440
rect 191006 2388 191012 2440
rect 191064 2428 191070 2440
rect 191837 2431 191895 2437
rect 191064 2400 191420 2428
rect 191064 2388 191070 2400
rect 191392 2372 191420 2400
rect 191837 2397 191849 2431
rect 191883 2428 191895 2431
rect 192202 2428 192208 2440
rect 191883 2400 192208 2428
rect 191883 2397 191895 2400
rect 191837 2391 191895 2397
rect 192202 2388 192208 2400
rect 192260 2388 192266 2440
rect 194689 2431 194747 2437
rect 194689 2397 194701 2431
rect 194735 2428 194747 2431
rect 195698 2428 195704 2440
rect 194735 2400 195704 2428
rect 194735 2397 194747 2400
rect 194689 2391 194747 2397
rect 195698 2388 195704 2400
rect 195756 2388 195762 2440
rect 196158 2388 196164 2440
rect 196216 2388 196222 2440
rect 196989 2431 197047 2437
rect 196989 2397 197001 2431
rect 197035 2428 197047 2431
rect 197538 2428 197544 2440
rect 197035 2400 197544 2428
rect 197035 2397 197047 2400
rect 196989 2391 197047 2397
rect 197538 2388 197544 2400
rect 197596 2388 197602 2440
rect 197817 2431 197875 2437
rect 197817 2397 197829 2431
rect 197863 2428 197875 2431
rect 198274 2428 198280 2440
rect 197863 2400 198280 2428
rect 197863 2397 197875 2400
rect 197817 2391 197875 2397
rect 198274 2388 198280 2400
rect 198332 2388 198338 2440
rect 198553 2431 198611 2437
rect 198553 2397 198565 2431
rect 198599 2428 198611 2431
rect 199746 2428 199752 2440
rect 198599 2400 199752 2428
rect 198599 2397 198611 2400
rect 198553 2391 198611 2397
rect 199746 2388 199752 2400
rect 199804 2388 199810 2440
rect 200206 2388 200212 2440
rect 200264 2388 200270 2440
rect 201034 2388 201040 2440
rect 201092 2388 201098 2440
rect 201773 2431 201831 2437
rect 201773 2397 201785 2431
rect 201819 2428 201831 2431
rect 202690 2428 202696 2440
rect 201819 2400 202696 2428
rect 201819 2397 201831 2400
rect 201773 2391 201831 2397
rect 202690 2388 202696 2400
rect 202748 2388 202754 2440
rect 203150 2388 203156 2440
rect 203208 2388 203214 2440
rect 203260 2437 203288 2468
rect 203245 2431 203303 2437
rect 203245 2397 203257 2431
rect 203291 2397 203303 2431
rect 203245 2391 203303 2397
rect 203429 2431 203487 2437
rect 203429 2397 203441 2431
rect 203475 2428 203487 2431
rect 203889 2431 203947 2437
rect 203889 2428 203901 2431
rect 203475 2400 203901 2428
rect 203475 2397 203487 2400
rect 203429 2391 203487 2397
rect 203889 2397 203901 2400
rect 203935 2397 203947 2431
rect 203889 2391 203947 2397
rect 172480 2332 179920 2360
rect 172480 2320 172486 2332
rect 191190 2320 191196 2372
rect 191248 2320 191254 2372
rect 191374 2320 191380 2372
rect 191432 2360 191438 2372
rect 207584 2360 207612 2536
rect 218146 2524 218152 2576
rect 218204 2524 218210 2576
rect 219084 2564 219112 2604
rect 219250 2592 219256 2644
rect 219308 2632 219314 2644
rect 219345 2635 219403 2641
rect 219345 2632 219357 2635
rect 219308 2604 219357 2632
rect 219308 2592 219314 2604
rect 219345 2601 219357 2604
rect 219391 2601 219403 2635
rect 224494 2632 224500 2644
rect 219345 2595 219403 2601
rect 219452 2604 224500 2632
rect 219452 2564 219480 2604
rect 224494 2592 224500 2604
rect 224552 2632 224558 2644
rect 224552 2604 226932 2632
rect 224552 2592 224558 2604
rect 219084 2536 219480 2564
rect 222010 2524 222016 2576
rect 222068 2564 222074 2576
rect 225782 2564 225788 2576
rect 222068 2536 225788 2564
rect 222068 2524 222074 2536
rect 225782 2524 225788 2536
rect 225840 2524 225846 2576
rect 226904 2564 226932 2604
rect 226978 2592 226984 2644
rect 227036 2592 227042 2644
rect 227070 2592 227076 2644
rect 227128 2632 227134 2644
rect 228266 2632 228272 2644
rect 227128 2604 228272 2632
rect 227128 2592 227134 2604
rect 228266 2592 228272 2604
rect 228324 2592 228330 2644
rect 243906 2632 243912 2644
rect 228376 2604 243912 2632
rect 228376 2564 228404 2604
rect 243906 2592 243912 2604
rect 243964 2592 243970 2644
rect 245470 2592 245476 2644
rect 245528 2632 245534 2644
rect 248874 2632 248880 2644
rect 245528 2604 248880 2632
rect 245528 2592 245534 2604
rect 248874 2592 248880 2604
rect 248932 2592 248938 2644
rect 250640 2604 263594 2632
rect 226904 2536 228404 2564
rect 228450 2524 228456 2576
rect 228508 2564 228514 2576
rect 230566 2564 230572 2576
rect 228508 2536 230572 2564
rect 228508 2524 228514 2536
rect 230566 2524 230572 2536
rect 230624 2524 230630 2576
rect 230750 2524 230756 2576
rect 230808 2564 230814 2576
rect 230937 2567 230995 2573
rect 230937 2564 230949 2567
rect 230808 2536 230949 2564
rect 230808 2524 230814 2536
rect 230937 2533 230949 2536
rect 230983 2533 230995 2567
rect 230937 2527 230995 2533
rect 233050 2524 233056 2576
rect 233108 2564 233114 2576
rect 246850 2564 246856 2576
rect 233108 2536 246856 2564
rect 233108 2524 233114 2536
rect 246850 2524 246856 2536
rect 246908 2524 246914 2576
rect 248506 2524 248512 2576
rect 248564 2564 248570 2576
rect 248564 2536 250208 2564
rect 248564 2524 248570 2536
rect 209682 2496 209688 2508
rect 208320 2468 209688 2496
rect 208320 2437 208348 2468
rect 209682 2456 209688 2468
rect 209740 2456 209746 2508
rect 210053 2499 210111 2505
rect 210053 2465 210065 2499
rect 210099 2496 210111 2499
rect 210099 2468 212304 2496
rect 210099 2465 210111 2468
rect 210053 2459 210111 2465
rect 208305 2431 208363 2437
rect 208305 2397 208317 2431
rect 208351 2397 208363 2431
rect 208305 2391 208363 2397
rect 208670 2388 208676 2440
rect 208728 2428 208734 2440
rect 208857 2431 208915 2437
rect 208857 2428 208869 2431
rect 208728 2400 208869 2428
rect 208728 2388 208734 2400
rect 208857 2397 208869 2400
rect 208903 2397 208915 2431
rect 208857 2391 208915 2397
rect 208946 2388 208952 2440
rect 209004 2388 209010 2440
rect 209038 2388 209044 2440
rect 209096 2428 209102 2440
rect 209133 2431 209191 2437
rect 209133 2428 209145 2431
rect 209096 2400 209145 2428
rect 209096 2388 209102 2400
rect 209133 2397 209145 2400
rect 209179 2397 209191 2431
rect 209133 2391 209191 2397
rect 209501 2431 209559 2437
rect 209501 2397 209513 2431
rect 209547 2428 209559 2431
rect 209547 2400 210096 2428
rect 209547 2397 209559 2400
rect 209501 2391 209559 2397
rect 191432 2332 207612 2360
rect 210068 2360 210096 2400
rect 210237 2363 210295 2369
rect 210237 2360 210249 2363
rect 210068 2332 210249 2360
rect 191432 2320 191438 2332
rect 210237 2329 210249 2332
rect 210283 2329 210295 2363
rect 210237 2323 210295 2329
rect 211890 2320 211896 2372
rect 211948 2320 211954 2372
rect 168340 2264 168972 2292
rect 168340 2252 168346 2264
rect 191006 2252 191012 2304
rect 191064 2292 191070 2304
rect 191285 2295 191343 2301
rect 191285 2292 191297 2295
rect 191064 2264 191297 2292
rect 191064 2252 191070 2264
rect 191285 2261 191297 2264
rect 191331 2261 191343 2295
rect 191285 2255 191343 2261
rect 194594 2252 194600 2304
rect 194652 2292 194658 2304
rect 194873 2295 194931 2301
rect 194873 2292 194885 2295
rect 194652 2264 194885 2292
rect 194652 2252 194658 2264
rect 194873 2261 194885 2264
rect 194919 2261 194931 2295
rect 194873 2255 194931 2261
rect 196066 2252 196072 2304
rect 196124 2292 196130 2304
rect 196345 2295 196403 2301
rect 196345 2292 196357 2295
rect 196124 2264 196357 2292
rect 196124 2252 196130 2264
rect 196345 2261 196357 2264
rect 196391 2261 196403 2295
rect 196345 2255 196403 2261
rect 196618 2252 196624 2304
rect 196676 2292 196682 2304
rect 197173 2295 197231 2301
rect 197173 2292 197185 2295
rect 196676 2264 197185 2292
rect 196676 2252 196682 2264
rect 197173 2261 197185 2264
rect 197219 2261 197231 2295
rect 197173 2255 197231 2261
rect 197354 2252 197360 2304
rect 197412 2292 197418 2304
rect 198001 2295 198059 2301
rect 198001 2292 198013 2295
rect 197412 2264 198013 2292
rect 197412 2252 197418 2264
rect 198001 2261 198013 2264
rect 198047 2261 198059 2295
rect 198001 2255 198059 2261
rect 201218 2252 201224 2304
rect 201276 2252 201282 2304
rect 204070 2252 204076 2304
rect 204128 2252 204134 2304
rect 208118 2252 208124 2304
rect 208176 2252 208182 2304
rect 212276 2292 212304 2468
rect 212534 2456 212540 2508
rect 212592 2456 212598 2508
rect 213822 2456 213828 2508
rect 213880 2496 213886 2508
rect 215389 2499 215447 2505
rect 215389 2496 215401 2499
rect 213880 2468 215401 2496
rect 213880 2456 213886 2468
rect 215389 2465 215401 2468
rect 215435 2465 215447 2499
rect 215389 2459 215447 2465
rect 216766 2456 216772 2508
rect 216824 2456 216830 2508
rect 217502 2456 217508 2508
rect 217560 2456 217566 2508
rect 217594 2456 217600 2508
rect 217652 2496 217658 2508
rect 221826 2496 221832 2508
rect 217652 2468 221832 2496
rect 217652 2456 217658 2468
rect 221826 2456 221832 2468
rect 221884 2456 221890 2508
rect 223114 2456 223120 2508
rect 223172 2456 223178 2508
rect 240042 2496 240048 2508
rect 223224 2468 227208 2496
rect 212350 2388 212356 2440
rect 212408 2388 212414 2440
rect 214193 2431 214251 2437
rect 214193 2397 214205 2431
rect 214239 2428 214251 2431
rect 214374 2428 214380 2440
rect 214239 2400 214380 2428
rect 214239 2397 214251 2400
rect 214193 2391 214251 2397
rect 214374 2388 214380 2400
rect 214432 2388 214438 2440
rect 215205 2431 215263 2437
rect 215205 2428 215217 2431
rect 215128 2400 215217 2428
rect 214466 2292 214472 2304
rect 212276 2264 214472 2292
rect 214466 2252 214472 2264
rect 214524 2252 214530 2304
rect 215128 2292 215156 2400
rect 215205 2397 215217 2400
rect 215251 2397 215263 2431
rect 215205 2391 215263 2397
rect 217686 2388 217692 2440
rect 217744 2388 217750 2440
rect 218422 2388 218428 2440
rect 218480 2388 218486 2440
rect 218606 2437 218612 2440
rect 218563 2431 218612 2437
rect 218563 2397 218575 2431
rect 218609 2397 218612 2431
rect 218563 2391 218612 2397
rect 218606 2388 218612 2391
rect 218664 2388 218670 2440
rect 218698 2388 218704 2440
rect 218756 2388 218762 2440
rect 220538 2388 220544 2440
rect 220596 2388 220602 2440
rect 220630 2388 220636 2440
rect 220688 2388 220694 2440
rect 220725 2431 220783 2437
rect 220725 2397 220737 2431
rect 220771 2428 220783 2431
rect 220814 2428 220820 2440
rect 220771 2400 220820 2428
rect 220771 2397 220783 2400
rect 220725 2391 220783 2397
rect 220814 2388 220820 2400
rect 220872 2388 220878 2440
rect 221366 2388 221372 2440
rect 221424 2388 221430 2440
rect 220909 2363 220967 2369
rect 220909 2329 220921 2363
rect 220955 2360 220967 2363
rect 221553 2363 221611 2369
rect 221553 2360 221565 2363
rect 220955 2332 221565 2360
rect 220955 2329 220967 2332
rect 220909 2323 220967 2329
rect 221553 2329 221565 2332
rect 221599 2329 221611 2363
rect 221553 2323 221611 2329
rect 222562 2320 222568 2372
rect 222620 2360 222626 2372
rect 223224 2360 223252 2468
rect 224037 2431 224095 2437
rect 224037 2397 224049 2431
rect 224083 2428 224095 2431
rect 224126 2428 224132 2440
rect 224083 2400 224132 2428
rect 224083 2397 224095 2400
rect 224037 2391 224095 2397
rect 224126 2388 224132 2400
rect 224184 2388 224190 2440
rect 224957 2431 225015 2437
rect 224957 2397 224969 2431
rect 225003 2397 225015 2431
rect 224957 2391 225015 2397
rect 225509 2431 225567 2437
rect 225509 2397 225521 2431
rect 225555 2428 225567 2431
rect 225782 2428 225788 2440
rect 225555 2400 225788 2428
rect 225555 2397 225567 2400
rect 225509 2391 225567 2397
rect 224972 2360 225000 2391
rect 225782 2388 225788 2400
rect 225840 2388 225846 2440
rect 226245 2431 226303 2437
rect 226245 2397 226257 2431
rect 226291 2428 226303 2431
rect 226794 2428 226800 2440
rect 226291 2400 226800 2428
rect 226291 2397 226303 2400
rect 226245 2391 226303 2397
rect 226794 2388 226800 2400
rect 226852 2388 226858 2440
rect 227180 2437 227208 2468
rect 229066 2468 240048 2496
rect 227165 2431 227223 2437
rect 227165 2397 227177 2431
rect 227211 2397 227223 2431
rect 227165 2391 227223 2397
rect 227809 2431 227867 2437
rect 227809 2397 227821 2431
rect 227855 2428 227867 2431
rect 228450 2428 228456 2440
rect 227855 2400 228456 2428
rect 227855 2397 227867 2400
rect 227809 2391 227867 2397
rect 228450 2388 228456 2400
rect 228508 2388 228514 2440
rect 222620 2332 223252 2360
rect 223316 2332 225000 2360
rect 222620 2320 222626 2332
rect 219618 2292 219624 2304
rect 215128 2264 219624 2292
rect 219618 2252 219624 2264
rect 219676 2252 219682 2304
rect 219710 2252 219716 2304
rect 219768 2292 219774 2304
rect 223316 2292 223344 2332
rect 225414 2320 225420 2372
rect 225472 2360 225478 2372
rect 229066 2360 229094 2468
rect 240042 2456 240048 2468
rect 240100 2456 240106 2508
rect 242894 2456 242900 2508
rect 242952 2496 242958 2508
rect 246117 2499 246175 2505
rect 246117 2496 246129 2499
rect 242952 2468 246129 2496
rect 242952 2456 242958 2468
rect 246117 2465 246129 2468
rect 246163 2465 246175 2499
rect 246117 2459 246175 2465
rect 248598 2456 248604 2508
rect 248656 2496 248662 2508
rect 248969 2499 249027 2505
rect 248969 2496 248981 2499
rect 248656 2468 248981 2496
rect 248656 2456 248662 2468
rect 248969 2465 248981 2468
rect 249015 2465 249027 2499
rect 248969 2459 249027 2465
rect 229833 2431 229891 2437
rect 229833 2397 229845 2431
rect 229879 2428 229891 2431
rect 230934 2428 230940 2440
rect 229879 2400 230940 2428
rect 229879 2397 229891 2400
rect 229833 2391 229891 2397
rect 230934 2388 230940 2400
rect 230992 2388 230998 2440
rect 231397 2431 231455 2437
rect 231397 2397 231409 2431
rect 231443 2428 231455 2431
rect 231762 2428 231768 2440
rect 231443 2400 231768 2428
rect 231443 2397 231455 2400
rect 231397 2391 231455 2397
rect 231762 2388 231768 2400
rect 231820 2388 231826 2440
rect 232225 2431 232283 2437
rect 232225 2397 232237 2431
rect 232271 2428 232283 2431
rect 232590 2428 232596 2440
rect 232271 2400 232596 2428
rect 232271 2397 232283 2400
rect 232225 2391 232283 2397
rect 232590 2388 232596 2400
rect 232648 2388 232654 2440
rect 232958 2388 232964 2440
rect 233016 2388 233022 2440
rect 234982 2388 234988 2440
rect 235040 2388 235046 2440
rect 235810 2388 235816 2440
rect 235868 2388 235874 2440
rect 235997 2431 236055 2437
rect 235997 2397 236009 2431
rect 236043 2397 236055 2431
rect 235997 2391 236055 2397
rect 236641 2431 236699 2437
rect 236641 2397 236653 2431
rect 236687 2428 236699 2431
rect 236914 2428 236920 2440
rect 236687 2400 236920 2428
rect 236687 2397 236699 2400
rect 236641 2391 236699 2397
rect 225472 2332 229094 2360
rect 225472 2320 225478 2332
rect 229922 2320 229928 2372
rect 229980 2360 229986 2372
rect 230753 2363 230811 2369
rect 230753 2360 230765 2363
rect 229980 2332 230765 2360
rect 229980 2320 229986 2332
rect 230753 2329 230765 2332
rect 230799 2360 230811 2363
rect 236012 2360 236040 2391
rect 236914 2388 236920 2400
rect 236972 2388 236978 2440
rect 243446 2388 243452 2440
rect 243504 2388 243510 2440
rect 243722 2388 243728 2440
rect 243780 2388 243786 2440
rect 244182 2388 244188 2440
rect 244240 2428 244246 2440
rect 244737 2431 244795 2437
rect 244737 2428 244749 2431
rect 244240 2400 244749 2428
rect 244240 2388 244246 2400
rect 244737 2397 244749 2400
rect 244783 2397 244795 2431
rect 244737 2391 244795 2397
rect 245010 2388 245016 2440
rect 245068 2388 245074 2440
rect 248782 2388 248788 2440
rect 248840 2388 248846 2440
rect 250180 2428 250208 2536
rect 250640 2505 250668 2604
rect 256510 2524 256516 2576
rect 256568 2524 256574 2576
rect 259730 2524 259736 2576
rect 259788 2564 259794 2576
rect 259788 2536 261708 2564
rect 259788 2524 259794 2536
rect 250625 2499 250683 2505
rect 250625 2465 250637 2499
rect 250671 2465 250683 2499
rect 250625 2459 250683 2465
rect 251450 2456 251456 2508
rect 251508 2456 251514 2508
rect 253474 2456 253480 2508
rect 253532 2496 253538 2508
rect 253845 2499 253903 2505
rect 253845 2496 253857 2499
rect 253532 2468 253857 2496
rect 253532 2456 253538 2468
rect 253845 2465 253857 2468
rect 253891 2465 253903 2499
rect 256528 2496 256556 2524
rect 256605 2499 256663 2505
rect 256605 2496 256617 2499
rect 256528 2468 256617 2496
rect 253845 2459 253903 2465
rect 256605 2465 256617 2468
rect 256651 2465 256663 2499
rect 256605 2459 256663 2465
rect 258261 2499 258319 2505
rect 258261 2465 258273 2499
rect 258307 2496 258319 2499
rect 258307 2468 260972 2496
rect 258307 2465 258319 2468
rect 258261 2459 258319 2465
rect 251269 2431 251327 2437
rect 251269 2428 251281 2431
rect 250180 2400 251281 2428
rect 251269 2397 251281 2400
rect 251315 2397 251327 2431
rect 251269 2391 251327 2397
rect 252646 2388 252652 2440
rect 252704 2428 252710 2440
rect 253569 2431 253627 2437
rect 253569 2428 253581 2431
rect 252704 2400 253581 2428
rect 252704 2388 252710 2400
rect 253569 2397 253581 2400
rect 253615 2397 253627 2431
rect 253569 2391 253627 2397
rect 254854 2388 254860 2440
rect 254912 2388 254918 2440
rect 255133 2431 255191 2437
rect 255133 2397 255145 2431
rect 255179 2397 255191 2431
rect 255133 2391 255191 2397
rect 230799 2332 236040 2360
rect 230799 2329 230811 2332
rect 230753 2323 230811 2329
rect 246298 2320 246304 2372
rect 246356 2320 246362 2372
rect 247957 2363 248015 2369
rect 247957 2329 247969 2363
rect 248003 2360 248015 2363
rect 252370 2360 252376 2372
rect 248003 2332 252376 2360
rect 248003 2329 248015 2332
rect 247957 2323 248015 2329
rect 252370 2320 252376 2332
rect 252428 2320 252434 2372
rect 253106 2320 253112 2372
rect 253164 2320 253170 2372
rect 219768 2264 223344 2292
rect 219768 2252 219774 2264
rect 224218 2252 224224 2304
rect 224276 2252 224282 2304
rect 224770 2252 224776 2304
rect 224828 2252 224834 2304
rect 225690 2252 225696 2304
rect 225748 2252 225754 2304
rect 226334 2252 226340 2304
rect 226392 2292 226398 2304
rect 226429 2295 226487 2301
rect 226429 2292 226441 2295
rect 226392 2264 226441 2292
rect 226392 2252 226398 2264
rect 226429 2261 226441 2264
rect 226475 2261 226487 2295
rect 226429 2255 226487 2261
rect 227990 2252 227996 2304
rect 228048 2252 228054 2304
rect 230014 2252 230020 2304
rect 230072 2252 230078 2304
rect 231578 2252 231584 2304
rect 231636 2252 231642 2304
rect 232406 2252 232412 2304
rect 232464 2252 232470 2304
rect 233142 2252 233148 2304
rect 233200 2252 233206 2304
rect 235166 2252 235172 2304
rect 235224 2252 235230 2304
rect 236178 2252 236184 2304
rect 236236 2252 236242 2304
rect 236822 2252 236828 2304
rect 236880 2252 236886 2304
rect 243630 2252 243636 2304
rect 243688 2292 243694 2304
rect 255148 2292 255176 2391
rect 256418 2388 256424 2440
rect 256476 2388 256482 2440
rect 258721 2431 258779 2437
rect 258721 2428 258733 2431
rect 257816 2400 258733 2428
rect 257522 2320 257528 2372
rect 257580 2360 257586 2372
rect 257816 2360 257844 2400
rect 258721 2397 258733 2400
rect 258767 2397 258779 2431
rect 258721 2391 258779 2397
rect 258997 2431 259055 2437
rect 258997 2397 259009 2431
rect 259043 2397 259055 2431
rect 258997 2391 259055 2397
rect 257580 2332 257844 2360
rect 257580 2320 257586 2332
rect 258350 2320 258356 2372
rect 258408 2360 258414 2372
rect 259012 2360 259040 2391
rect 258408 2332 259040 2360
rect 258408 2320 258414 2332
rect 260098 2320 260104 2372
rect 260156 2320 260162 2372
rect 260944 2360 260972 2468
rect 261570 2456 261576 2508
rect 261628 2456 261634 2508
rect 261680 2496 261708 2536
rect 262214 2524 262220 2576
rect 262272 2564 262278 2576
rect 262585 2567 262643 2573
rect 262585 2564 262597 2567
rect 262272 2536 262597 2564
rect 262272 2524 262278 2536
rect 262585 2533 262597 2536
rect 262631 2533 262643 2567
rect 263566 2564 263594 2604
rect 266998 2592 267004 2644
rect 267056 2632 267062 2644
rect 268289 2635 268347 2641
rect 268289 2632 268301 2635
rect 267056 2604 268301 2632
rect 267056 2592 267062 2604
rect 268289 2601 268301 2604
rect 268335 2601 268347 2635
rect 268289 2595 268347 2601
rect 269850 2592 269856 2644
rect 269908 2632 269914 2644
rect 270129 2635 270187 2641
rect 270129 2632 270141 2635
rect 269908 2604 270141 2632
rect 269908 2592 269914 2604
rect 270129 2601 270141 2604
rect 270175 2601 270187 2635
rect 270129 2595 270187 2601
rect 267918 2564 267924 2576
rect 263566 2536 267924 2564
rect 262585 2527 262643 2533
rect 267918 2524 267924 2536
rect 267976 2524 267982 2576
rect 261680 2468 263594 2496
rect 261018 2388 261024 2440
rect 261076 2428 261082 2440
rect 261478 2428 261484 2440
rect 261076 2400 261484 2428
rect 261076 2388 261082 2400
rect 261478 2388 261484 2400
rect 261536 2428 261542 2440
rect 261757 2431 261815 2437
rect 261757 2428 261769 2431
rect 261536 2400 261769 2428
rect 261536 2388 261542 2400
rect 261757 2397 261769 2400
rect 261803 2397 261815 2431
rect 261757 2391 261815 2397
rect 261941 2431 261999 2437
rect 261941 2397 261953 2431
rect 261987 2428 261999 2431
rect 262401 2431 262459 2437
rect 262401 2428 262413 2431
rect 261987 2400 262413 2428
rect 261987 2397 261999 2400
rect 261941 2391 261999 2397
rect 262401 2397 262413 2400
rect 262447 2397 262459 2431
rect 262401 2391 262459 2397
rect 263134 2388 263140 2440
rect 263192 2388 263198 2440
rect 263566 2428 263594 2468
rect 263962 2456 263968 2508
rect 264020 2456 264026 2508
rect 264885 2499 264943 2505
rect 264885 2496 264897 2499
rect 264072 2468 264897 2496
rect 264072 2428 264100 2468
rect 264885 2465 264897 2468
rect 264931 2465 264943 2499
rect 264885 2459 264943 2465
rect 267550 2456 267556 2508
rect 267608 2496 267614 2508
rect 267608 2468 268608 2496
rect 267608 2456 267614 2468
rect 263566 2400 264100 2428
rect 264149 2431 264207 2437
rect 264149 2397 264161 2431
rect 264195 2428 264207 2431
rect 264330 2428 264336 2440
rect 264195 2400 264336 2428
rect 264195 2397 264207 2400
rect 264149 2391 264207 2397
rect 264330 2388 264336 2400
rect 264388 2388 264394 2440
rect 265158 2388 265164 2440
rect 265216 2388 265222 2440
rect 266725 2431 266783 2437
rect 266725 2397 266737 2431
rect 266771 2428 266783 2431
rect 266998 2428 267004 2440
rect 266771 2400 267004 2428
rect 266771 2397 266783 2400
rect 266725 2391 266783 2397
rect 266998 2388 267004 2400
rect 267056 2388 267062 2440
rect 267829 2431 267887 2437
rect 267829 2397 267841 2431
rect 267875 2428 267887 2431
rect 268286 2428 268292 2440
rect 267875 2400 268292 2428
rect 267875 2397 267887 2400
rect 267829 2391 267887 2397
rect 268286 2388 268292 2400
rect 268344 2388 268350 2440
rect 268470 2388 268476 2440
rect 268528 2388 268534 2440
rect 268580 2428 268608 2468
rect 268654 2456 268660 2508
rect 268712 2496 268718 2508
rect 269761 2499 269819 2505
rect 269761 2496 269773 2499
rect 268712 2468 269773 2496
rect 268712 2456 268718 2468
rect 269761 2465 269773 2468
rect 269807 2465 269819 2499
rect 269761 2459 269819 2465
rect 268933 2431 268991 2437
rect 268933 2428 268945 2431
rect 268580 2400 268945 2428
rect 268933 2397 268945 2400
rect 268979 2397 268991 2431
rect 268933 2391 268991 2397
rect 269114 2388 269120 2440
rect 269172 2428 269178 2440
rect 269945 2431 270003 2437
rect 269945 2428 269957 2431
rect 269172 2400 269957 2428
rect 269172 2388 269178 2400
rect 269945 2397 269957 2400
rect 269991 2397 270003 2431
rect 269945 2391 270003 2397
rect 270034 2388 270040 2440
rect 270092 2428 270098 2440
rect 270589 2431 270647 2437
rect 270589 2428 270601 2431
rect 270092 2400 270601 2428
rect 270092 2388 270098 2400
rect 270589 2397 270601 2400
rect 270635 2397 270647 2431
rect 270589 2391 270647 2397
rect 263962 2360 263968 2372
rect 260944 2332 263968 2360
rect 263962 2320 263968 2332
rect 264020 2320 264026 2372
rect 264238 2320 264244 2372
rect 264296 2360 264302 2372
rect 268378 2360 268384 2372
rect 264296 2332 268384 2360
rect 264296 2320 264302 2332
rect 268378 2320 268384 2332
rect 268436 2320 268442 2372
rect 243688 2264 255176 2292
rect 243688 2252 243694 2264
rect 259914 2252 259920 2304
rect 259972 2292 259978 2304
rect 260190 2292 260196 2304
rect 259972 2264 260196 2292
rect 259972 2252 259978 2264
rect 260190 2252 260196 2264
rect 260248 2252 260254 2304
rect 263318 2252 263324 2304
rect 263376 2252 263382 2304
rect 264333 2295 264391 2301
rect 264333 2261 264345 2295
rect 264379 2292 264391 2295
rect 264882 2292 264888 2304
rect 264379 2264 264888 2292
rect 264379 2261 264391 2264
rect 264333 2255 264391 2261
rect 264882 2252 264888 2264
rect 264940 2252 264946 2304
rect 266906 2252 266912 2304
rect 266964 2252 266970 2304
rect 267645 2295 267703 2301
rect 267645 2261 267657 2295
rect 267691 2292 267703 2295
rect 269206 2292 269212 2304
rect 267691 2264 269212 2292
rect 267691 2261 267703 2264
rect 267645 2255 267703 2261
rect 269206 2252 269212 2264
rect 269264 2252 269270 2304
rect 269301 2295 269359 2301
rect 269301 2261 269313 2295
rect 269347 2292 269359 2295
rect 270126 2292 270132 2304
rect 269347 2264 270132 2292
rect 269347 2261 269359 2264
rect 269301 2255 269359 2261
rect 270126 2252 270132 2264
rect 270184 2252 270190 2304
rect 270770 2252 270776 2304
rect 270828 2252 270834 2304
rect 1104 2202 271651 2224
rect 1104 2150 68546 2202
rect 68598 2150 68610 2202
rect 68662 2150 68674 2202
rect 68726 2150 68738 2202
rect 68790 2150 68802 2202
rect 68854 2150 136143 2202
rect 136195 2150 136207 2202
rect 136259 2150 136271 2202
rect 136323 2150 136335 2202
rect 136387 2150 136399 2202
rect 136451 2150 203740 2202
rect 203792 2150 203804 2202
rect 203856 2150 203868 2202
rect 203920 2150 203932 2202
rect 203984 2150 203996 2202
rect 204048 2150 271337 2202
rect 271389 2150 271401 2202
rect 271453 2150 271465 2202
rect 271517 2150 271529 2202
rect 271581 2150 271593 2202
rect 271645 2150 271651 2202
rect 1104 2128 271651 2150
rect 1765 2091 1823 2097
rect 1765 2057 1777 2091
rect 1811 2088 1823 2091
rect 1854 2088 1860 2100
rect 1811 2060 1860 2088
rect 1811 2057 1823 2060
rect 1765 2051 1823 2057
rect 1854 2048 1860 2060
rect 1912 2048 1918 2100
rect 12066 2048 12072 2100
rect 12124 2048 12130 2100
rect 12802 2048 12808 2100
rect 12860 2048 12866 2100
rect 15764 2060 37596 2088
rect 6886 1992 15608 2020
rect 1670 1912 1676 1964
rect 1728 1912 1734 1964
rect 4065 1955 4123 1961
rect 4065 1921 4077 1955
rect 4111 1952 4123 1955
rect 5534 1952 5540 1964
rect 4111 1924 5540 1952
rect 4111 1921 4123 1924
rect 4065 1915 4123 1921
rect 5534 1912 5540 1924
rect 5592 1912 5598 1964
rect 3786 1844 3792 1896
rect 3844 1844 3850 1896
rect 5166 1844 5172 1896
rect 5224 1844 5230 1896
rect 5445 1887 5503 1893
rect 5445 1853 5457 1887
rect 5491 1884 5503 1887
rect 6886 1884 6914 1992
rect 7374 1912 7380 1964
rect 7432 1912 7438 1964
rect 8662 1912 8668 1964
rect 8720 1912 8726 1964
rect 11974 1912 11980 1964
rect 12032 1912 12038 1964
rect 12710 1912 12716 1964
rect 12768 1912 12774 1964
rect 14366 1912 14372 1964
rect 14424 1912 14430 1964
rect 5491 1856 6914 1884
rect 5491 1853 5503 1856
rect 5445 1847 5503 1853
rect 7098 1844 7104 1896
rect 7156 1844 7162 1896
rect 8386 1844 8392 1896
rect 8444 1844 8450 1896
rect 9674 1844 9680 1896
rect 9732 1844 9738 1896
rect 9953 1887 10011 1893
rect 9953 1853 9965 1887
rect 9999 1853 10011 1887
rect 9953 1847 10011 1853
rect 9968 1816 9996 1847
rect 14090 1844 14096 1896
rect 14148 1844 14154 1896
rect 15470 1844 15476 1896
rect 15528 1844 15534 1896
rect 15580 1884 15608 1992
rect 15764 1961 15792 2060
rect 15838 1980 15844 2032
rect 15896 2020 15902 2032
rect 15896 1992 25084 2020
rect 15896 1980 15902 1992
rect 15749 1955 15807 1961
rect 15749 1921 15761 1955
rect 15795 1921 15807 1955
rect 15749 1915 15807 1921
rect 17862 1912 17868 1964
rect 17920 1912 17926 1964
rect 18046 1912 18052 1964
rect 18104 1912 18110 1964
rect 21177 1955 21235 1961
rect 21177 1921 21189 1955
rect 21223 1952 21235 1955
rect 22186 1952 22192 1964
rect 21223 1924 22192 1952
rect 21223 1921 21235 1924
rect 21177 1915 21235 1921
rect 22186 1912 22192 1924
rect 22244 1912 22250 1964
rect 22278 1912 22284 1964
rect 22336 1912 22342 1964
rect 22370 1912 22376 1964
rect 22428 1952 22434 1964
rect 22428 1924 23244 1952
rect 22428 1912 22434 1924
rect 22097 1887 22155 1893
rect 15580 1856 15976 1884
rect 15838 1816 15844 1828
rect 9968 1788 15844 1816
rect 15838 1776 15844 1788
rect 15896 1776 15902 1828
rect 15948 1816 15976 1856
rect 22097 1853 22109 1887
rect 22143 1884 22155 1887
rect 22462 1884 22468 1896
rect 22143 1856 22468 1884
rect 22143 1853 22155 1856
rect 22097 1847 22155 1853
rect 22462 1844 22468 1856
rect 22520 1844 22526 1896
rect 22833 1887 22891 1893
rect 22833 1853 22845 1887
rect 22879 1884 22891 1887
rect 23106 1884 23112 1896
rect 22879 1856 23112 1884
rect 22879 1853 22891 1856
rect 22833 1847 22891 1853
rect 23106 1844 23112 1856
rect 23164 1844 23170 1896
rect 23216 1884 23244 1924
rect 23290 1912 23296 1964
rect 23348 1912 23354 1964
rect 23477 1955 23535 1961
rect 23477 1921 23489 1955
rect 23523 1952 23535 1955
rect 24029 1955 24087 1961
rect 24029 1952 24041 1955
rect 23523 1924 24041 1952
rect 23523 1921 23535 1924
rect 23477 1915 23535 1921
rect 24029 1921 24041 1924
rect 24075 1921 24087 1955
rect 24029 1915 24087 1921
rect 24118 1912 24124 1964
rect 24176 1952 24182 1964
rect 24176 1924 24440 1952
rect 24176 1912 24182 1924
rect 24305 1887 24363 1893
rect 24305 1884 24317 1887
rect 23216 1856 24317 1884
rect 24305 1853 24317 1856
rect 24351 1853 24363 1887
rect 24412 1884 24440 1924
rect 24946 1912 24952 1964
rect 25004 1912 25010 1964
rect 25056 1952 25084 1992
rect 25866 1980 25872 2032
rect 25924 1980 25930 2032
rect 37568 2020 37596 2060
rect 37642 2048 37648 2100
rect 37700 2088 37706 2100
rect 37921 2091 37979 2097
rect 37921 2088 37933 2091
rect 37700 2060 37933 2088
rect 37700 2048 37706 2060
rect 37921 2057 37933 2060
rect 37967 2057 37979 2091
rect 37921 2051 37979 2057
rect 38470 2048 38476 2100
rect 38528 2088 38534 2100
rect 40586 2088 40592 2100
rect 38528 2060 40592 2088
rect 38528 2048 38534 2060
rect 38562 2020 38568 2032
rect 26206 1992 35894 2020
rect 37568 1992 38568 2020
rect 26206 1952 26234 1992
rect 25056 1924 26234 1952
rect 26326 1912 26332 1964
rect 26384 1952 26390 1964
rect 27338 1952 27344 1964
rect 26384 1924 27344 1952
rect 26384 1912 26390 1924
rect 27338 1912 27344 1924
rect 27396 1952 27402 1964
rect 27893 1955 27951 1961
rect 27893 1952 27905 1955
rect 27396 1924 27905 1952
rect 27396 1912 27402 1924
rect 27893 1921 27905 1924
rect 27939 1952 27951 1955
rect 28721 1955 28779 1961
rect 28721 1952 28733 1955
rect 27939 1924 28733 1952
rect 27939 1921 27951 1924
rect 27893 1915 27951 1921
rect 28721 1921 28733 1924
rect 28767 1952 28779 1955
rect 29549 1955 29607 1961
rect 29549 1952 29561 1955
rect 28767 1924 29561 1952
rect 28767 1921 28779 1924
rect 28721 1915 28779 1921
rect 29549 1921 29561 1924
rect 29595 1952 29607 1955
rect 30193 1955 30251 1961
rect 30193 1952 30205 1955
rect 29595 1924 30205 1952
rect 29595 1921 29607 1924
rect 29549 1915 29607 1921
rect 30193 1921 30205 1924
rect 30239 1952 30251 1955
rect 31205 1955 31263 1961
rect 31205 1952 31217 1955
rect 30239 1924 31217 1952
rect 30239 1921 30251 1924
rect 30193 1915 30251 1921
rect 31205 1921 31217 1924
rect 31251 1952 31263 1955
rect 32490 1952 32496 1964
rect 31251 1924 32496 1952
rect 31251 1921 31263 1924
rect 31205 1915 31263 1921
rect 32490 1912 32496 1924
rect 32548 1912 32554 1964
rect 32674 1912 32680 1964
rect 32732 1952 32738 1964
rect 33137 1955 33195 1961
rect 33137 1952 33149 1955
rect 32732 1924 33149 1952
rect 32732 1912 32738 1924
rect 33137 1921 33149 1924
rect 33183 1921 33195 1955
rect 33137 1915 33195 1921
rect 27614 1884 27620 1896
rect 24412 1856 27620 1884
rect 24305 1847 24363 1853
rect 27614 1844 27620 1856
rect 27672 1844 27678 1896
rect 27706 1844 27712 1896
rect 27764 1844 27770 1896
rect 28534 1844 28540 1896
rect 28592 1844 28598 1896
rect 29365 1887 29423 1893
rect 29365 1853 29377 1887
rect 29411 1884 29423 1887
rect 29454 1884 29460 1896
rect 29411 1856 29460 1884
rect 29411 1853 29423 1856
rect 29365 1847 29423 1853
rect 29454 1844 29460 1856
rect 29512 1844 29518 1896
rect 29730 1844 29736 1896
rect 29788 1844 29794 1896
rect 30009 1887 30067 1893
rect 30009 1853 30021 1887
rect 30055 1884 30067 1887
rect 30098 1884 30104 1896
rect 30055 1856 30104 1884
rect 30055 1853 30067 1856
rect 30009 1847 30067 1853
rect 30098 1844 30104 1856
rect 30156 1844 30162 1896
rect 30742 1844 30748 1896
rect 30800 1884 30806 1896
rect 31021 1887 31079 1893
rect 31021 1884 31033 1887
rect 30800 1856 31033 1884
rect 30800 1844 30806 1856
rect 31021 1853 31033 1856
rect 31067 1884 31079 1887
rect 31294 1884 31300 1896
rect 31067 1856 31300 1884
rect 31067 1853 31079 1856
rect 31021 1847 31079 1853
rect 31294 1844 31300 1856
rect 31352 1844 31358 1896
rect 31846 1844 31852 1896
rect 31904 1884 31910 1896
rect 32309 1887 32367 1893
rect 32309 1884 32321 1887
rect 31904 1856 32321 1884
rect 31904 1844 31910 1856
rect 32309 1853 32321 1856
rect 32355 1853 32367 1887
rect 35866 1884 35894 1992
rect 38562 1980 38568 1992
rect 38620 1980 38626 2032
rect 39022 2020 39028 2032
rect 38856 1992 39028 2020
rect 38102 1912 38108 1964
rect 38160 1912 38166 1964
rect 38856 1884 38884 1992
rect 39022 1980 39028 1992
rect 39080 1980 39086 2032
rect 39117 2023 39175 2029
rect 39117 1989 39129 2023
rect 39163 2020 39175 2023
rect 39298 2020 39304 2032
rect 39163 1992 39304 2020
rect 39163 1989 39175 1992
rect 39117 1983 39175 1989
rect 39298 1980 39304 1992
rect 39356 1980 39362 2032
rect 39390 1980 39396 2032
rect 39448 1980 39454 2032
rect 39500 2029 39528 2060
rect 40586 2048 40592 2060
rect 40644 2048 40650 2100
rect 41506 2048 41512 2100
rect 41564 2088 41570 2100
rect 73430 2088 73436 2100
rect 41564 2060 73436 2088
rect 41564 2048 41570 2060
rect 73430 2048 73436 2060
rect 73488 2048 73494 2100
rect 73614 2048 73620 2100
rect 73672 2088 73678 2100
rect 80054 2088 80060 2100
rect 73672 2060 80060 2088
rect 73672 2048 73678 2060
rect 80054 2048 80060 2060
rect 80112 2048 80118 2100
rect 89257 2091 89315 2097
rect 89257 2057 89269 2091
rect 89303 2088 89315 2091
rect 89346 2088 89352 2100
rect 89303 2060 89352 2088
rect 89303 2057 89315 2060
rect 89257 2051 89315 2057
rect 89346 2048 89352 2060
rect 89404 2048 89410 2100
rect 90266 2048 90272 2100
rect 90324 2048 90330 2100
rect 91094 2048 91100 2100
rect 91152 2048 91158 2100
rect 91830 2048 91836 2100
rect 91888 2088 91894 2100
rect 91925 2091 91983 2097
rect 91925 2088 91937 2091
rect 91888 2060 91937 2088
rect 91888 2048 91894 2060
rect 91925 2057 91937 2060
rect 91971 2057 91983 2091
rect 91925 2051 91983 2057
rect 93210 2048 93216 2100
rect 93268 2088 93274 2100
rect 93581 2091 93639 2097
rect 93581 2088 93593 2091
rect 93268 2060 93593 2088
rect 93268 2048 93274 2060
rect 93581 2057 93593 2060
rect 93627 2057 93639 2091
rect 93581 2051 93639 2057
rect 94130 2048 94136 2100
rect 94188 2088 94194 2100
rect 94593 2091 94651 2097
rect 94593 2088 94605 2091
rect 94188 2060 94605 2088
rect 94188 2048 94194 2060
rect 94593 2057 94605 2060
rect 94639 2057 94651 2091
rect 94593 2051 94651 2057
rect 94682 2048 94688 2100
rect 94740 2088 94746 2100
rect 96062 2088 96068 2100
rect 94740 2060 96068 2088
rect 94740 2048 94746 2060
rect 96062 2048 96068 2060
rect 96120 2048 96126 2100
rect 96430 2048 96436 2100
rect 96488 2048 96494 2100
rect 97902 2088 97908 2100
rect 97092 2060 97908 2088
rect 39485 2023 39543 2029
rect 39485 1989 39497 2023
rect 39531 1989 39543 2023
rect 39485 1983 39543 1989
rect 39574 1980 39580 2032
rect 39632 2020 39638 2032
rect 39853 2023 39911 2029
rect 39853 2020 39865 2023
rect 39632 1992 39865 2020
rect 39632 1980 39638 1992
rect 39853 1989 39865 1992
rect 39899 1989 39911 2023
rect 39853 1983 39911 1989
rect 40034 1980 40040 2032
rect 40092 2020 40098 2032
rect 40221 2023 40279 2029
rect 40221 2020 40233 2023
rect 40092 1992 40233 2020
rect 40092 1980 40098 1992
rect 40221 1989 40233 1992
rect 40267 1989 40279 2023
rect 40221 1983 40279 1989
rect 53282 1980 53288 2032
rect 53340 1980 53346 2032
rect 54021 2023 54079 2029
rect 54021 1989 54033 2023
rect 54067 2020 54079 2023
rect 55490 2020 55496 2032
rect 54067 1992 55496 2020
rect 54067 1989 54079 1992
rect 54021 1983 54079 1989
rect 55490 1980 55496 1992
rect 55548 1980 55554 2032
rect 56226 2020 56232 2032
rect 55600 1992 56232 2020
rect 45462 1912 45468 1964
rect 45520 1912 45526 1964
rect 52733 1955 52791 1961
rect 52733 1921 52745 1955
rect 52779 1952 52791 1955
rect 53742 1952 53748 1964
rect 52779 1924 53748 1952
rect 52779 1921 52791 1924
rect 52733 1915 52791 1921
rect 53742 1912 53748 1924
rect 53800 1912 53806 1964
rect 53837 1955 53895 1961
rect 53837 1921 53849 1955
rect 53883 1952 53895 1955
rect 54202 1952 54208 1964
rect 53883 1924 54208 1952
rect 53883 1921 53895 1924
rect 53837 1915 53895 1921
rect 54202 1912 54208 1924
rect 54260 1952 54266 1964
rect 54570 1952 54576 1964
rect 54260 1924 54576 1952
rect 54260 1912 54266 1924
rect 54570 1912 54576 1924
rect 54628 1952 54634 1964
rect 55600 1961 55628 1992
rect 56226 1980 56232 1992
rect 56284 1980 56290 2032
rect 57514 1980 57520 2032
rect 57572 1980 57578 2032
rect 59170 1980 59176 2032
rect 59228 1980 59234 2032
rect 61654 1980 61660 2032
rect 61712 1980 61718 2032
rect 62666 1980 62672 2032
rect 62724 1980 62730 2032
rect 63144 1992 64276 2020
rect 54849 1955 54907 1961
rect 54849 1952 54861 1955
rect 54628 1924 54861 1952
rect 54628 1912 54634 1924
rect 54849 1921 54861 1924
rect 54895 1952 54907 1955
rect 55585 1955 55643 1961
rect 54895 1924 55214 1952
rect 54895 1921 54907 1924
rect 54849 1915 54907 1921
rect 35866 1856 38884 1884
rect 40132 1896 40184 1902
rect 32309 1847 32367 1853
rect 41046 1884 41052 1896
rect 40184 1856 41052 1884
rect 41046 1844 41052 1856
rect 41104 1844 41110 1896
rect 53282 1844 53288 1896
rect 53340 1884 53346 1896
rect 53653 1887 53711 1893
rect 53653 1884 53665 1887
rect 53340 1856 53665 1884
rect 53340 1844 53346 1856
rect 53653 1853 53665 1856
rect 53699 1884 53711 1887
rect 54110 1884 54116 1896
rect 53699 1856 54116 1884
rect 53699 1853 53711 1856
rect 53653 1847 53711 1853
rect 54110 1844 54116 1856
rect 54168 1844 54174 1896
rect 54665 1887 54723 1893
rect 54665 1884 54677 1887
rect 54312 1856 54677 1884
rect 40132 1838 40184 1844
rect 38378 1816 38384 1828
rect 15948 1788 38384 1816
rect 38378 1776 38384 1788
rect 38436 1776 38442 1828
rect 45278 1776 45284 1828
rect 45336 1776 45342 1828
rect 54312 1760 54340 1856
rect 54665 1853 54677 1856
rect 54711 1853 54723 1887
rect 55186 1884 55214 1924
rect 55585 1921 55597 1955
rect 55631 1921 55643 1955
rect 55585 1915 55643 1921
rect 55677 1955 55735 1961
rect 55677 1921 55689 1955
rect 55723 1921 55735 1955
rect 55677 1915 55735 1921
rect 55692 1884 55720 1915
rect 56410 1912 56416 1964
rect 56468 1912 56474 1964
rect 56505 1955 56563 1961
rect 56505 1921 56517 1955
rect 56551 1921 56563 1955
rect 56505 1915 56563 1921
rect 56520 1884 56548 1915
rect 56870 1912 56876 1964
rect 56928 1952 56934 1964
rect 57149 1955 57207 1961
rect 57149 1952 57161 1955
rect 56928 1924 57161 1952
rect 56928 1912 56934 1924
rect 57149 1921 57161 1924
rect 57195 1921 57207 1955
rect 57149 1915 57207 1921
rect 57333 1955 57391 1961
rect 57333 1921 57345 1955
rect 57379 1921 57391 1955
rect 57333 1915 57391 1921
rect 57348 1884 57376 1915
rect 58066 1912 58072 1964
rect 58124 1912 58130 1964
rect 58618 1912 58624 1964
rect 58676 1952 58682 1964
rect 58805 1955 58863 1961
rect 58805 1952 58817 1955
rect 58676 1924 58817 1952
rect 58676 1912 58682 1924
rect 58805 1921 58817 1924
rect 58851 1921 58863 1955
rect 58805 1915 58863 1921
rect 58989 1955 59047 1961
rect 58989 1921 59001 1955
rect 59035 1921 59047 1955
rect 58989 1915 59047 1921
rect 58526 1884 58532 1896
rect 55186 1856 58532 1884
rect 54665 1847 54723 1853
rect 54680 1816 54708 1847
rect 58526 1844 58532 1856
rect 58584 1884 58590 1896
rect 59004 1884 59032 1915
rect 59722 1912 59728 1964
rect 59780 1912 59786 1964
rect 59814 1912 59820 1964
rect 59872 1912 59878 1964
rect 60550 1912 60556 1964
rect 60608 1912 60614 1964
rect 60645 1955 60703 1961
rect 60645 1921 60657 1955
rect 60691 1921 60703 1955
rect 60645 1915 60703 1921
rect 59832 1884 59860 1912
rect 58584 1856 59860 1884
rect 60660 1884 60688 1915
rect 61286 1912 61292 1964
rect 61344 1912 61350 1964
rect 61473 1955 61531 1961
rect 61473 1921 61485 1955
rect 61519 1921 61531 1955
rect 61473 1915 61531 1921
rect 61488 1884 61516 1915
rect 62298 1912 62304 1964
rect 62356 1912 62362 1964
rect 62482 1912 62488 1964
rect 62540 1952 62546 1964
rect 63144 1952 63172 1992
rect 62540 1924 63172 1952
rect 62540 1912 62546 1924
rect 63218 1912 63224 1964
rect 63276 1952 63282 1964
rect 63604 1961 63632 1992
rect 63405 1955 63463 1961
rect 63405 1952 63417 1955
rect 63276 1924 63417 1952
rect 63276 1912 63282 1924
rect 63405 1921 63417 1924
rect 63451 1921 63463 1955
rect 63405 1915 63463 1921
rect 63589 1955 63647 1961
rect 63589 1921 63601 1955
rect 63635 1921 63647 1955
rect 63589 1915 63647 1921
rect 64046 1912 64052 1964
rect 64104 1912 64110 1964
rect 64248 1961 64276 1992
rect 65426 1980 65432 2032
rect 65484 1980 65490 2032
rect 66162 1980 66168 2032
rect 66220 2020 66226 2032
rect 89533 2023 89591 2029
rect 89533 2020 89545 2023
rect 66220 1992 66484 2020
rect 66220 1980 66226 1992
rect 64233 1955 64291 1961
rect 64233 1921 64245 1955
rect 64279 1952 64291 1955
rect 65245 1955 65303 1961
rect 65245 1952 65257 1955
rect 64279 1924 65257 1952
rect 64279 1921 64291 1924
rect 64233 1915 64291 1921
rect 65245 1921 65257 1924
rect 65291 1952 65303 1955
rect 66180 1952 66208 1980
rect 65291 1924 66208 1952
rect 65291 1921 65303 1924
rect 65245 1915 65303 1921
rect 66346 1912 66352 1964
rect 66404 1912 66410 1964
rect 66456 1961 66484 1992
rect 73632 1992 89545 2020
rect 73632 1964 73660 1992
rect 89533 1989 89545 1992
rect 89579 2020 89591 2023
rect 89898 2020 89904 2032
rect 89579 1992 89904 2020
rect 89579 1989 89591 1992
rect 89533 1983 89591 1989
rect 89898 1980 89904 1992
rect 89956 1980 89962 2032
rect 91002 2020 91008 2032
rect 90836 1992 91008 2020
rect 66441 1955 66499 1961
rect 66441 1921 66453 1955
rect 66487 1921 66499 1955
rect 66441 1915 66499 1921
rect 66625 1955 66683 1961
rect 66625 1921 66637 1955
rect 66671 1952 66683 1955
rect 67085 1955 67143 1961
rect 67085 1952 67097 1955
rect 66671 1924 67097 1952
rect 66671 1921 66683 1924
rect 66625 1915 66683 1921
rect 67085 1921 67097 1924
rect 67131 1921 67143 1955
rect 67085 1915 67143 1921
rect 71498 1912 71504 1964
rect 71556 1912 71562 1964
rect 72234 1912 72240 1964
rect 72292 1912 72298 1964
rect 73614 1912 73620 1964
rect 73672 1912 73678 1964
rect 73706 1912 73712 1964
rect 73764 1912 73770 1964
rect 78582 1952 78588 1964
rect 76024 1924 78588 1952
rect 62500 1884 62528 1912
rect 60660 1856 62528 1884
rect 64785 1887 64843 1893
rect 58584 1844 58590 1856
rect 64785 1853 64797 1887
rect 64831 1884 64843 1887
rect 65058 1884 65064 1896
rect 64831 1856 65064 1884
rect 64831 1853 64843 1856
rect 64785 1847 64843 1853
rect 65058 1844 65064 1856
rect 65116 1844 65122 1896
rect 71332 1856 74304 1884
rect 55582 1816 55588 1828
rect 54680 1788 55588 1816
rect 55582 1776 55588 1788
rect 55640 1816 55646 1828
rect 71332 1825 71360 1856
rect 71317 1819 71375 1825
rect 55640 1788 67634 1816
rect 55640 1776 55646 1788
rect 21361 1751 21419 1757
rect 21361 1717 21373 1751
rect 21407 1748 21419 1751
rect 22002 1748 22008 1760
rect 21407 1720 22008 1748
rect 21407 1717 21419 1720
rect 21361 1711 21419 1717
rect 22002 1708 22008 1720
rect 22060 1708 22066 1760
rect 22094 1708 22100 1760
rect 22152 1748 22158 1760
rect 22465 1751 22523 1757
rect 22465 1748 22477 1751
rect 22152 1720 22477 1748
rect 22152 1708 22158 1720
rect 22465 1717 22477 1720
rect 22511 1717 22523 1751
rect 22465 1711 22523 1717
rect 22554 1708 22560 1760
rect 22612 1748 22618 1760
rect 23753 1751 23811 1757
rect 23753 1748 23765 1751
rect 22612 1720 23765 1748
rect 22612 1708 22618 1720
rect 23753 1717 23765 1720
rect 23799 1748 23811 1751
rect 24118 1748 24124 1760
rect 23799 1720 24124 1748
rect 23799 1717 23811 1720
rect 23753 1711 23811 1717
rect 24118 1708 24124 1720
rect 24176 1708 24182 1760
rect 25038 1708 25044 1760
rect 25096 1708 25102 1760
rect 25958 1708 25964 1760
rect 26016 1708 26022 1760
rect 27982 1708 27988 1760
rect 28040 1748 28046 1760
rect 28077 1751 28135 1757
rect 28077 1748 28089 1751
rect 28040 1720 28089 1748
rect 28040 1708 28046 1720
rect 28077 1717 28089 1720
rect 28123 1717 28135 1751
rect 28077 1711 28135 1717
rect 28810 1708 28816 1760
rect 28868 1748 28874 1760
rect 28905 1751 28963 1757
rect 28905 1748 28917 1751
rect 28868 1720 28917 1748
rect 28868 1708 28874 1720
rect 28905 1717 28917 1720
rect 28951 1717 28963 1751
rect 28905 1711 28963 1717
rect 30374 1708 30380 1760
rect 30432 1708 30438 1760
rect 31018 1708 31024 1760
rect 31076 1748 31082 1760
rect 31389 1751 31447 1757
rect 31389 1748 31401 1751
rect 31076 1720 31401 1748
rect 31076 1708 31082 1720
rect 31389 1717 31401 1720
rect 31435 1717 31447 1751
rect 31389 1711 31447 1717
rect 32306 1708 32312 1760
rect 32364 1748 32370 1760
rect 32677 1751 32735 1757
rect 32677 1748 32689 1751
rect 32364 1720 32689 1748
rect 32364 1708 32370 1720
rect 32677 1717 32689 1720
rect 32723 1717 32735 1751
rect 32677 1711 32735 1717
rect 33134 1708 33140 1760
rect 33192 1748 33198 1760
rect 33321 1751 33379 1757
rect 33321 1748 33333 1751
rect 33192 1720 33333 1748
rect 33192 1708 33198 1720
rect 33321 1717 33333 1720
rect 33367 1717 33379 1751
rect 33321 1711 33379 1717
rect 35158 1708 35164 1760
rect 35216 1708 35222 1760
rect 40402 1708 40408 1760
rect 40460 1708 40466 1760
rect 52914 1708 52920 1760
rect 52972 1708 52978 1760
rect 54294 1708 54300 1760
rect 54352 1708 54358 1760
rect 55030 1708 55036 1760
rect 55088 1708 55094 1760
rect 55861 1751 55919 1757
rect 55861 1717 55873 1751
rect 55907 1748 55919 1751
rect 56226 1748 56232 1760
rect 55907 1720 56232 1748
rect 55907 1717 55919 1720
rect 55861 1711 55919 1717
rect 56226 1708 56232 1720
rect 56284 1708 56290 1760
rect 56689 1751 56747 1757
rect 56689 1717 56701 1751
rect 56735 1748 56747 1751
rect 56962 1748 56968 1760
rect 56735 1720 56968 1748
rect 56735 1717 56747 1720
rect 56689 1711 56747 1717
rect 56962 1708 56968 1720
rect 57020 1708 57026 1760
rect 58250 1708 58256 1760
rect 58308 1708 58314 1760
rect 59814 1708 59820 1760
rect 59872 1748 59878 1760
rect 60001 1751 60059 1757
rect 60001 1748 60013 1751
rect 59872 1720 60013 1748
rect 59872 1708 59878 1720
rect 60001 1717 60013 1720
rect 60047 1717 60059 1751
rect 60001 1711 60059 1717
rect 60734 1708 60740 1760
rect 60792 1748 60798 1760
rect 60829 1751 60887 1757
rect 60829 1748 60841 1751
rect 60792 1720 60841 1748
rect 60792 1708 60798 1720
rect 60829 1717 60841 1720
rect 60875 1717 60887 1751
rect 60829 1711 60887 1717
rect 63678 1708 63684 1760
rect 63736 1748 63742 1760
rect 63773 1751 63831 1757
rect 63773 1748 63785 1751
rect 63736 1720 63785 1748
rect 63736 1708 63742 1720
rect 63773 1717 63785 1720
rect 63819 1717 63831 1751
rect 63773 1711 63831 1717
rect 64414 1708 64420 1760
rect 64472 1708 64478 1760
rect 67266 1708 67272 1760
rect 67324 1708 67330 1760
rect 67606 1748 67634 1788
rect 71317 1785 71329 1819
rect 71363 1785 71375 1819
rect 71317 1779 71375 1785
rect 72050 1776 72056 1828
rect 72108 1776 72114 1828
rect 73430 1776 73436 1828
rect 73488 1816 73494 1828
rect 73525 1819 73583 1825
rect 73525 1816 73537 1819
rect 73488 1788 73537 1816
rect 73488 1776 73494 1788
rect 73525 1785 73537 1788
rect 73571 1785 73583 1819
rect 73525 1779 73583 1785
rect 73338 1748 73344 1760
rect 67606 1720 73344 1748
rect 73338 1708 73344 1720
rect 73396 1708 73402 1760
rect 74276 1748 74304 1856
rect 75730 1844 75736 1896
rect 75788 1844 75794 1896
rect 76024 1893 76052 1924
rect 78582 1912 78588 1924
rect 78640 1912 78646 1964
rect 79689 1955 79747 1961
rect 79689 1921 79701 1955
rect 79735 1952 79747 1955
rect 79735 1924 81112 1952
rect 79735 1921 79747 1924
rect 79689 1915 79747 1921
rect 76009 1887 76067 1893
rect 76009 1853 76021 1887
rect 76055 1853 76067 1887
rect 76009 1847 76067 1853
rect 77202 1844 77208 1896
rect 77260 1844 77266 1896
rect 77478 1844 77484 1896
rect 77536 1844 77542 1896
rect 79410 1844 79416 1896
rect 79468 1844 79474 1896
rect 80882 1844 80888 1896
rect 80940 1844 80946 1896
rect 81084 1884 81112 1924
rect 81158 1912 81164 1964
rect 81216 1912 81222 1964
rect 81268 1924 84792 1952
rect 81268 1884 81296 1924
rect 81084 1856 81296 1884
rect 82354 1844 82360 1896
rect 82412 1844 82418 1896
rect 82630 1844 82636 1896
rect 82688 1844 82694 1896
rect 84562 1844 84568 1896
rect 84620 1844 84626 1896
rect 84764 1884 84792 1924
rect 84838 1912 84844 1964
rect 84896 1912 84902 1964
rect 86313 1955 86371 1961
rect 84948 1924 86172 1952
rect 84948 1884 84976 1924
rect 84764 1856 84976 1884
rect 86034 1844 86040 1896
rect 86092 1844 86098 1896
rect 86144 1884 86172 1924
rect 86313 1921 86325 1955
rect 86359 1952 86371 1955
rect 86862 1952 86868 1964
rect 86359 1924 86868 1952
rect 86359 1921 86371 1924
rect 86313 1915 86371 1921
rect 86862 1912 86868 1924
rect 86920 1912 86926 1964
rect 88153 1955 88211 1961
rect 88153 1921 88165 1955
rect 88199 1952 88211 1955
rect 88242 1952 88248 1964
rect 88199 1924 88248 1952
rect 88199 1921 88211 1924
rect 88153 1915 88211 1921
rect 88242 1912 88248 1924
rect 88300 1912 88306 1964
rect 89070 1912 89076 1964
rect 89128 1952 89134 1964
rect 90836 1961 90864 1992
rect 91002 1980 91008 1992
rect 91060 1980 91066 2032
rect 93762 1980 93768 2032
rect 93820 2020 93826 2032
rect 97092 2020 97120 2060
rect 97902 2048 97908 2060
rect 97960 2048 97966 2100
rect 98730 2048 98736 2100
rect 98788 2048 98794 2100
rect 98822 2048 98828 2100
rect 98880 2088 98886 2100
rect 107654 2088 107660 2100
rect 98880 2060 101904 2088
rect 98880 2048 98886 2060
rect 93820 1992 97120 2020
rect 99469 2023 99527 2029
rect 93820 1980 93826 1992
rect 99469 1989 99481 2023
rect 99515 2020 99527 2023
rect 99926 2020 99932 2032
rect 99515 1992 99932 2020
rect 99515 1989 99527 1992
rect 99469 1983 99527 1989
rect 99926 1980 99932 1992
rect 99984 1980 99990 2032
rect 101030 1980 101036 2032
rect 101088 2020 101094 2032
rect 101125 2023 101183 2029
rect 101125 2020 101137 2023
rect 101088 1992 101137 2020
rect 101088 1980 101094 1992
rect 101125 1989 101137 1992
rect 101171 1989 101183 2023
rect 101125 1983 101183 1989
rect 90085 1955 90143 1961
rect 90085 1952 90097 1955
rect 89128 1924 90097 1952
rect 89128 1912 89134 1924
rect 90085 1921 90097 1924
rect 90131 1921 90143 1955
rect 90085 1915 90143 1921
rect 90821 1955 90879 1961
rect 90821 1921 90833 1955
rect 90867 1921 90879 1955
rect 90821 1915 90879 1921
rect 90913 1955 90971 1961
rect 90913 1921 90925 1955
rect 90959 1921 90971 1955
rect 90913 1915 90971 1921
rect 88518 1884 88524 1896
rect 86144 1856 88524 1884
rect 88518 1844 88524 1856
rect 88576 1844 88582 1896
rect 88889 1887 88947 1893
rect 88889 1853 88901 1887
rect 88935 1884 88947 1887
rect 89622 1884 89628 1896
rect 88935 1856 89628 1884
rect 88935 1853 88947 1856
rect 88889 1847 88947 1853
rect 89622 1844 89628 1856
rect 89680 1844 89686 1896
rect 89898 1844 89904 1896
rect 89956 1844 89962 1896
rect 90100 1884 90128 1915
rect 90726 1884 90732 1896
rect 90100 1856 90732 1884
rect 90726 1844 90732 1856
rect 90784 1884 90790 1896
rect 90928 1884 90956 1915
rect 91646 1912 91652 1964
rect 91704 1912 91710 1964
rect 91741 1955 91799 1961
rect 91741 1921 91753 1955
rect 91787 1952 91799 1955
rect 92566 1952 92572 1964
rect 91787 1924 92572 1952
rect 91787 1921 91799 1924
rect 91741 1915 91799 1921
rect 91756 1884 91784 1915
rect 92566 1912 92572 1924
rect 92624 1912 92630 1964
rect 93118 1912 93124 1964
rect 93176 1952 93182 1964
rect 93213 1955 93271 1961
rect 93213 1952 93225 1955
rect 93176 1924 93225 1952
rect 93176 1912 93182 1924
rect 93213 1921 93225 1924
rect 93259 1921 93271 1955
rect 93213 1915 93271 1921
rect 93397 1955 93455 1961
rect 93397 1921 93409 1955
rect 93443 1952 93455 1955
rect 93443 1924 94176 1952
rect 93443 1921 93455 1924
rect 93397 1915 93455 1921
rect 90784 1856 91784 1884
rect 90784 1844 90790 1856
rect 92382 1844 92388 1896
rect 92440 1844 92446 1896
rect 92584 1884 92612 1912
rect 93486 1884 93492 1896
rect 92584 1856 93492 1884
rect 93486 1844 93492 1856
rect 93544 1844 93550 1896
rect 94148 1884 94176 1924
rect 94222 1912 94228 1964
rect 94280 1912 94286 1964
rect 94409 1955 94467 1961
rect 94409 1921 94421 1955
rect 94455 1952 94467 1955
rect 95421 1955 95479 1961
rect 95421 1952 95433 1955
rect 94455 1924 95433 1952
rect 94455 1921 94467 1924
rect 94409 1915 94467 1921
rect 95421 1921 95433 1924
rect 95467 1921 95479 1955
rect 95421 1915 95479 1921
rect 94424 1884 94452 1915
rect 94148 1856 94452 1884
rect 94961 1887 95019 1893
rect 94961 1853 94973 1887
rect 95007 1884 95019 1887
rect 95050 1884 95056 1896
rect 95007 1856 95056 1884
rect 95007 1853 95019 1856
rect 94961 1847 95019 1853
rect 95050 1844 95056 1856
rect 95108 1884 95114 1896
rect 95237 1887 95295 1893
rect 95237 1884 95249 1887
rect 95108 1856 95249 1884
rect 95108 1844 95114 1856
rect 95237 1853 95249 1856
rect 95283 1853 95295 1887
rect 95436 1884 95464 1915
rect 95878 1912 95884 1964
rect 95936 1952 95942 1964
rect 96065 1955 96123 1961
rect 96065 1952 96077 1955
rect 95936 1924 96077 1952
rect 95936 1912 95942 1924
rect 96065 1921 96077 1924
rect 96111 1921 96123 1955
rect 96065 1915 96123 1921
rect 96249 1955 96307 1961
rect 96249 1921 96261 1955
rect 96295 1952 96307 1955
rect 96338 1952 96344 1964
rect 96295 1924 96344 1952
rect 96295 1921 96307 1924
rect 96249 1915 96307 1921
rect 95602 1884 95608 1896
rect 95436 1856 95608 1884
rect 95237 1847 95295 1853
rect 95602 1844 95608 1856
rect 95660 1884 95666 1896
rect 96264 1884 96292 1915
rect 96338 1912 96344 1924
rect 96396 1912 96402 1964
rect 96890 1912 96896 1964
rect 96948 1912 96954 1964
rect 97828 1912 97834 1964
rect 97886 1912 97892 1964
rect 97930 1955 97988 1961
rect 97930 1921 97942 1955
rect 97976 1952 97988 1955
rect 97976 1921 97994 1952
rect 97930 1918 97994 1921
rect 97930 1915 98040 1918
rect 95660 1856 96292 1884
rect 95660 1844 95666 1856
rect 97074 1844 97080 1896
rect 97132 1844 97138 1896
rect 97966 1890 98040 1915
rect 98086 1912 98092 1964
rect 98144 1912 98150 1964
rect 101876 1961 101904 2060
rect 103716 2060 107660 2088
rect 103716 2029 103744 2060
rect 107654 2048 107660 2060
rect 107712 2048 107718 2100
rect 107746 2048 107752 2100
rect 107804 2088 107810 2100
rect 108758 2088 108764 2100
rect 107804 2060 108764 2088
rect 107804 2048 107810 2060
rect 108758 2048 108764 2060
rect 108816 2048 108822 2100
rect 110874 2048 110880 2100
rect 110932 2088 110938 2100
rect 110932 2060 112484 2088
rect 110932 2048 110938 2060
rect 103701 2023 103759 2029
rect 103701 1989 103713 2023
rect 103747 1989 103759 2023
rect 103701 1983 103759 1989
rect 107381 2023 107439 2029
rect 107381 1989 107393 2023
rect 107427 2020 107439 2023
rect 107930 2020 107936 2032
rect 107427 1992 107936 2020
rect 107427 1989 107439 1992
rect 107381 1983 107439 1989
rect 107930 1980 107936 1992
rect 107988 1980 107994 2032
rect 108298 1980 108304 2032
rect 108356 2020 108362 2032
rect 110322 2020 110328 2032
rect 108356 1992 110328 2020
rect 108356 1980 108362 1992
rect 110322 1980 110328 1992
rect 110380 1980 110386 2032
rect 112456 2020 112484 2060
rect 112530 2048 112536 2100
rect 112588 2048 112594 2100
rect 114005 2091 114063 2097
rect 114005 2057 114017 2091
rect 114051 2057 114063 2091
rect 114005 2051 114063 2057
rect 114020 2020 114048 2051
rect 114554 2048 114560 2100
rect 114612 2088 114618 2100
rect 116857 2091 116915 2097
rect 114612 2060 116716 2088
rect 114612 2048 114618 2060
rect 112456 1992 114048 2020
rect 116688 2020 116716 2060
rect 116857 2057 116869 2091
rect 116903 2088 116915 2091
rect 118970 2088 118976 2100
rect 116903 2060 118976 2088
rect 116903 2057 116915 2060
rect 116857 2051 116915 2057
rect 118970 2048 118976 2060
rect 119028 2048 119034 2100
rect 119341 2091 119399 2097
rect 119341 2057 119353 2091
rect 119387 2088 119399 2091
rect 120718 2088 120724 2100
rect 119387 2060 120724 2088
rect 119387 2057 119399 2060
rect 119341 2051 119399 2057
rect 120718 2048 120724 2060
rect 120776 2048 120782 2100
rect 121086 2048 121092 2100
rect 121144 2048 121150 2100
rect 124306 2048 124312 2100
rect 124364 2048 124370 2100
rect 126698 2048 126704 2100
rect 126756 2048 126762 2100
rect 128354 2048 128360 2100
rect 128412 2048 128418 2100
rect 128464 2060 133644 2088
rect 117130 2020 117136 2032
rect 116688 1992 117136 2020
rect 117130 1980 117136 1992
rect 117188 1980 117194 2032
rect 117222 1980 117228 2032
rect 117280 1980 117286 2032
rect 101861 1955 101919 1961
rect 101861 1921 101873 1955
rect 101907 1921 101919 1955
rect 101861 1915 101919 1921
rect 104894 1912 104900 1964
rect 104952 1912 104958 1964
rect 105814 1912 105820 1964
rect 105872 1912 105878 1964
rect 105998 1961 106004 1964
rect 105955 1955 106004 1961
rect 105955 1921 105967 1955
rect 106001 1921 106004 1955
rect 105955 1915 106004 1921
rect 105998 1912 106004 1915
rect 106056 1912 106062 1964
rect 106090 1912 106096 1964
rect 106148 1912 106154 1964
rect 109589 1955 109647 1961
rect 109589 1921 109601 1955
rect 109635 1952 109647 1955
rect 110230 1952 110236 1964
rect 109635 1924 110236 1952
rect 109635 1921 109647 1924
rect 109589 1915 109647 1921
rect 110230 1912 110236 1924
rect 110288 1912 110294 1964
rect 110506 1912 110512 1964
rect 110564 1952 110570 1964
rect 110693 1955 110751 1961
rect 110693 1952 110705 1955
rect 110564 1924 110705 1952
rect 110564 1912 110570 1924
rect 110693 1921 110705 1924
rect 110739 1921 110751 1955
rect 110693 1915 110751 1921
rect 111886 1912 111892 1964
rect 111944 1912 111950 1964
rect 113545 1955 113603 1961
rect 113545 1921 113557 1955
rect 113591 1921 113603 1955
rect 113545 1915 113603 1921
rect 114189 1955 114247 1961
rect 114189 1921 114201 1955
rect 114235 1952 114247 1955
rect 114235 1924 115428 1952
rect 114235 1921 114247 1924
rect 114189 1915 114247 1921
rect 98012 1884 98040 1890
rect 98012 1856 99236 1884
rect 74626 1776 74632 1828
rect 74684 1816 74690 1828
rect 94038 1816 94044 1828
rect 74684 1788 94044 1816
rect 74684 1776 74690 1788
rect 94038 1776 94044 1788
rect 94096 1776 94102 1828
rect 94774 1776 94780 1828
rect 94832 1816 94838 1828
rect 97442 1816 97448 1828
rect 94832 1788 97448 1816
rect 94832 1776 94838 1788
rect 97442 1776 97448 1788
rect 97500 1816 97506 1828
rect 97537 1819 97595 1825
rect 97537 1816 97549 1819
rect 97500 1788 97549 1816
rect 97500 1776 97506 1788
rect 97537 1785 97549 1788
rect 97583 1785 97595 1819
rect 99208 1816 99236 1856
rect 99282 1844 99288 1896
rect 99340 1844 99346 1896
rect 101122 1844 101128 1896
rect 101180 1884 101186 1896
rect 102045 1887 102103 1893
rect 102045 1884 102057 1887
rect 101180 1856 102057 1884
rect 101180 1844 101186 1856
rect 102045 1853 102057 1856
rect 102091 1853 102103 1887
rect 102045 1847 102103 1853
rect 105078 1844 105084 1896
rect 105136 1844 105142 1896
rect 106737 1887 106795 1893
rect 105188 1856 106596 1884
rect 103238 1816 103244 1828
rect 97537 1779 97595 1785
rect 98656 1788 98868 1816
rect 99208 1788 103244 1816
rect 81434 1748 81440 1760
rect 74276 1720 81440 1748
rect 81434 1708 81440 1720
rect 81492 1708 81498 1760
rect 88334 1708 88340 1760
rect 88392 1708 88398 1760
rect 89898 1708 89904 1760
rect 89956 1748 89962 1760
rect 91370 1748 91376 1760
rect 89956 1720 91376 1748
rect 89956 1708 89962 1720
rect 91370 1708 91376 1720
rect 91428 1708 91434 1760
rect 91646 1708 91652 1760
rect 91704 1748 91710 1760
rect 92753 1751 92811 1757
rect 92753 1748 92765 1751
rect 91704 1720 92765 1748
rect 91704 1708 91710 1720
rect 92753 1717 92765 1720
rect 92799 1717 92811 1751
rect 92753 1711 92811 1717
rect 92934 1708 92940 1760
rect 92992 1748 92998 1760
rect 94590 1748 94596 1760
rect 92992 1720 94596 1748
rect 92992 1708 92998 1720
rect 94590 1708 94596 1720
rect 94648 1708 94654 1760
rect 95605 1751 95663 1757
rect 95605 1717 95617 1751
rect 95651 1748 95663 1751
rect 98656 1748 98684 1788
rect 95651 1720 98684 1748
rect 98840 1748 98868 1788
rect 103238 1776 103244 1788
rect 103296 1776 103302 1828
rect 104158 1776 104164 1828
rect 104216 1816 104222 1828
rect 105188 1816 105216 1856
rect 104216 1788 105216 1816
rect 105541 1819 105599 1825
rect 104216 1776 104222 1788
rect 105541 1785 105553 1819
rect 105587 1785 105599 1819
rect 106568 1816 106596 1856
rect 106737 1853 106749 1887
rect 106783 1884 106795 1887
rect 107197 1887 107255 1893
rect 107197 1884 107209 1887
rect 106783 1856 107209 1884
rect 106783 1853 106795 1856
rect 106737 1847 106795 1853
rect 107197 1853 107209 1856
rect 107243 1853 107255 1887
rect 107197 1847 107255 1853
rect 107654 1844 107660 1896
rect 107712 1884 107718 1896
rect 109126 1884 109132 1896
rect 107712 1856 109132 1884
rect 107712 1844 107718 1856
rect 109126 1844 109132 1856
rect 109184 1844 109190 1896
rect 109773 1887 109831 1893
rect 109773 1853 109785 1887
rect 109819 1853 109831 1887
rect 109773 1847 109831 1853
rect 108574 1816 108580 1828
rect 106568 1788 108580 1816
rect 105541 1779 105599 1785
rect 101674 1748 101680 1760
rect 98840 1720 101680 1748
rect 95651 1717 95663 1720
rect 95605 1711 95663 1717
rect 101674 1708 101680 1720
rect 101732 1708 101738 1760
rect 105556 1748 105584 1779
rect 108574 1776 108580 1788
rect 108632 1776 108638 1828
rect 107838 1748 107844 1760
rect 105556 1720 107844 1748
rect 107838 1708 107844 1720
rect 107896 1708 107902 1760
rect 107930 1708 107936 1760
rect 107988 1748 107994 1760
rect 109788 1748 109816 1847
rect 110874 1844 110880 1896
rect 110932 1844 110938 1896
rect 111613 1887 111671 1893
rect 111613 1884 111625 1887
rect 111444 1856 111625 1884
rect 111334 1776 111340 1828
rect 111392 1776 111398 1828
rect 107988 1720 109816 1748
rect 111444 1748 111472 1856
rect 111613 1853 111625 1856
rect 111659 1853 111671 1887
rect 111613 1847 111671 1853
rect 111751 1887 111809 1893
rect 111751 1853 111763 1887
rect 111797 1884 111809 1887
rect 113560 1884 113588 1915
rect 114830 1884 114836 1896
rect 111797 1856 113404 1884
rect 113560 1856 114836 1884
rect 111797 1853 111809 1856
rect 111751 1847 111809 1853
rect 113376 1825 113404 1856
rect 114830 1844 114836 1856
rect 114888 1844 114894 1896
rect 115014 1844 115020 1896
rect 115072 1844 115078 1896
rect 115198 1844 115204 1896
rect 115256 1844 115262 1896
rect 115400 1884 115428 1924
rect 115934 1912 115940 1964
rect 115992 1912 115998 1964
rect 116026 1912 116032 1964
rect 116084 1961 116090 1964
rect 116084 1955 116112 1961
rect 116100 1921 116112 1955
rect 116084 1915 116112 1921
rect 116084 1912 116090 1915
rect 116210 1912 116216 1964
rect 116268 1912 116274 1964
rect 117406 1912 117412 1964
rect 117464 1952 117470 1964
rect 117501 1955 117559 1961
rect 117501 1952 117513 1955
rect 117464 1924 117513 1952
rect 117464 1912 117470 1924
rect 117501 1921 117513 1924
rect 117547 1921 117559 1955
rect 117501 1915 117559 1921
rect 117682 1912 117688 1964
rect 117740 1912 117746 1964
rect 118421 1955 118479 1961
rect 118421 1921 118433 1955
rect 118467 1921 118479 1955
rect 118421 1915 118479 1921
rect 120077 1955 120135 1961
rect 120077 1921 120089 1955
rect 120123 1952 120135 1955
rect 120166 1952 120172 1964
rect 120123 1924 120172 1952
rect 120123 1921 120135 1924
rect 120077 1915 120135 1921
rect 115566 1884 115572 1896
rect 115400 1856 115572 1884
rect 115566 1844 115572 1856
rect 115624 1844 115630 1896
rect 118142 1884 118148 1896
rect 116596 1856 118148 1884
rect 113361 1819 113419 1825
rect 113361 1785 113373 1819
rect 113407 1785 113419 1819
rect 113361 1779 113419 1785
rect 115658 1776 115664 1828
rect 115716 1776 115722 1828
rect 111978 1748 111984 1760
rect 111444 1720 111984 1748
rect 107988 1708 107994 1720
rect 111978 1708 111984 1720
rect 112036 1708 112042 1760
rect 115676 1748 115704 1776
rect 116596 1748 116624 1856
rect 118142 1844 118148 1856
rect 118200 1844 118206 1896
rect 118436 1884 118464 1915
rect 120166 1912 120172 1924
rect 120224 1912 120230 1964
rect 120718 1912 120724 1964
rect 120776 1912 120782 1964
rect 121104 1952 121132 2048
rect 121730 1980 121736 2032
rect 121788 2020 121794 2032
rect 128464 2020 128492 2060
rect 121788 1992 128492 2020
rect 121788 1980 121794 1992
rect 131758 1980 131764 2032
rect 131816 1980 131822 2032
rect 133616 2020 133644 2060
rect 133690 2048 133696 2100
rect 133748 2048 133754 2100
rect 139486 2048 139492 2100
rect 139544 2088 139550 2100
rect 139581 2091 139639 2097
rect 139581 2088 139593 2091
rect 139544 2060 139593 2088
rect 139544 2048 139550 2060
rect 139581 2057 139593 2060
rect 139627 2057 139639 2091
rect 139581 2051 139639 2057
rect 139946 2048 139952 2100
rect 140004 2088 140010 2100
rect 140004 2060 140728 2088
rect 140004 2048 140010 2060
rect 138934 2020 138940 2032
rect 132512 1992 133460 2020
rect 133616 1992 138940 2020
rect 121454 1952 121460 1964
rect 121104 1924 121460 1952
rect 121454 1912 121460 1924
rect 121512 1912 121518 1964
rect 121641 1955 121699 1961
rect 121641 1921 121653 1955
rect 121687 1952 121699 1955
rect 122285 1955 122343 1961
rect 122285 1952 122297 1955
rect 121687 1924 122297 1952
rect 121687 1921 121699 1924
rect 121641 1915 121699 1921
rect 122285 1921 122297 1924
rect 122331 1952 122343 1955
rect 122650 1952 122656 1964
rect 122331 1924 122656 1952
rect 122331 1921 122343 1924
rect 122285 1915 122343 1921
rect 122650 1912 122656 1924
rect 122708 1952 122714 1964
rect 123297 1955 123355 1961
rect 123297 1952 123309 1955
rect 122708 1924 123309 1952
rect 122708 1912 122714 1924
rect 123297 1921 123309 1924
rect 123343 1952 123355 1955
rect 124125 1955 124183 1961
rect 124125 1952 124137 1955
rect 123343 1924 124137 1952
rect 123343 1921 123355 1924
rect 123297 1915 123355 1921
rect 124125 1921 124137 1924
rect 124171 1952 124183 1955
rect 124950 1952 124956 1964
rect 124171 1924 124956 1952
rect 124171 1921 124183 1924
rect 124125 1915 124183 1921
rect 124950 1912 124956 1924
rect 125008 1912 125014 1964
rect 125042 1912 125048 1964
rect 125100 1952 125106 1964
rect 125413 1955 125471 1961
rect 125413 1952 125425 1955
rect 125100 1924 125425 1952
rect 125100 1912 125106 1924
rect 125413 1921 125425 1924
rect 125459 1921 125471 1955
rect 125413 1915 125471 1921
rect 125597 1955 125655 1961
rect 125597 1921 125609 1955
rect 125643 1921 125655 1955
rect 125597 1915 125655 1921
rect 118252 1856 118464 1884
rect 115676 1720 116624 1748
rect 118142 1708 118148 1760
rect 118200 1748 118206 1760
rect 118252 1748 118280 1856
rect 118510 1844 118516 1896
rect 118568 1893 118574 1896
rect 118568 1887 118596 1893
rect 118584 1853 118596 1887
rect 118568 1847 118596 1853
rect 118697 1887 118755 1893
rect 118697 1853 118709 1887
rect 118743 1884 118755 1887
rect 119062 1884 119068 1896
rect 118743 1856 119068 1884
rect 118743 1853 118755 1856
rect 118697 1847 118755 1853
rect 118568 1844 118574 1847
rect 119062 1844 119068 1856
rect 119120 1844 119126 1896
rect 122098 1844 122104 1896
rect 122156 1844 122162 1896
rect 122834 1844 122840 1896
rect 122892 1884 122898 1896
rect 123110 1884 123116 1896
rect 122892 1856 123116 1884
rect 122892 1844 122898 1856
rect 123110 1844 123116 1856
rect 123168 1844 123174 1896
rect 123941 1887 123999 1893
rect 123941 1853 123953 1887
rect 123987 1884 123999 1887
rect 124030 1884 124036 1896
rect 123987 1856 124036 1884
rect 123987 1853 123999 1856
rect 123941 1847 123999 1853
rect 124030 1844 124036 1856
rect 124088 1844 124094 1896
rect 124968 1884 124996 1912
rect 125612 1884 125640 1915
rect 126330 1912 126336 1964
rect 126388 1912 126394 1964
rect 126517 1955 126575 1961
rect 126517 1921 126529 1955
rect 126563 1952 126575 1955
rect 127345 1955 127403 1961
rect 127345 1952 127357 1955
rect 126563 1924 127357 1952
rect 126563 1921 126575 1924
rect 126517 1915 126575 1921
rect 127345 1921 127357 1924
rect 127391 1952 127403 1955
rect 127391 1924 127848 1952
rect 127391 1921 127403 1924
rect 127345 1915 127403 1921
rect 126422 1884 126428 1896
rect 124968 1856 126428 1884
rect 126422 1844 126428 1856
rect 126480 1884 126486 1896
rect 126532 1884 126560 1915
rect 126480 1856 126560 1884
rect 127161 1887 127219 1893
rect 126480 1844 126486 1856
rect 127161 1853 127173 1887
rect 127207 1884 127219 1887
rect 127434 1884 127440 1896
rect 127207 1856 127440 1884
rect 127207 1853 127219 1856
rect 127161 1847 127219 1853
rect 127434 1844 127440 1856
rect 127492 1844 127498 1896
rect 127820 1884 127848 1924
rect 127986 1912 127992 1964
rect 128044 1912 128050 1964
rect 128173 1955 128231 1961
rect 128173 1921 128185 1955
rect 128219 1921 128231 1955
rect 128173 1915 128231 1921
rect 128188 1884 128216 1915
rect 128814 1912 128820 1964
rect 128872 1912 128878 1964
rect 130102 1912 130108 1964
rect 130160 1952 130166 1964
rect 130473 1955 130531 1961
rect 130473 1952 130485 1955
rect 130160 1924 130485 1952
rect 130160 1912 130166 1924
rect 130473 1921 130485 1924
rect 130519 1921 130531 1955
rect 130473 1915 130531 1921
rect 130657 1955 130715 1961
rect 130657 1921 130669 1955
rect 130703 1921 130715 1955
rect 130657 1915 130715 1921
rect 127820 1856 128216 1884
rect 129090 1844 129096 1896
rect 129148 1884 129154 1896
rect 129642 1884 129648 1896
rect 129148 1856 129648 1884
rect 129148 1844 129154 1856
rect 129642 1844 129648 1856
rect 129700 1884 129706 1896
rect 130672 1884 130700 1915
rect 131114 1912 131120 1964
rect 131172 1952 131178 1964
rect 131393 1955 131451 1961
rect 131393 1952 131405 1955
rect 131172 1924 131405 1952
rect 131172 1912 131178 1924
rect 131393 1921 131405 1924
rect 131439 1921 131451 1955
rect 131393 1915 131451 1921
rect 131577 1955 131635 1961
rect 131577 1921 131589 1955
rect 131623 1921 131635 1955
rect 131577 1915 131635 1921
rect 131592 1884 131620 1915
rect 131850 1912 131856 1964
rect 131908 1952 131914 1964
rect 132512 1961 132540 1992
rect 133432 1964 133460 1992
rect 138934 1980 138940 1992
rect 138992 1980 138998 2032
rect 140222 2020 140228 2032
rect 139136 1992 140228 2020
rect 132313 1955 132371 1961
rect 132313 1952 132325 1955
rect 131908 1924 132325 1952
rect 131908 1912 131914 1924
rect 132313 1921 132325 1924
rect 132359 1921 132371 1955
rect 132497 1955 132555 1961
rect 132497 1952 132509 1955
rect 132313 1915 132371 1921
rect 132420 1924 132509 1952
rect 132420 1884 132448 1924
rect 132497 1921 132509 1924
rect 132543 1921 132555 1955
rect 132497 1915 132555 1921
rect 132586 1912 132592 1964
rect 132644 1952 132650 1964
rect 133325 1955 133383 1961
rect 133325 1952 133337 1955
rect 132644 1924 133337 1952
rect 132644 1912 132650 1924
rect 133325 1921 133337 1924
rect 133371 1921 133383 1955
rect 133325 1915 133383 1921
rect 133414 1912 133420 1964
rect 133472 1952 133478 1964
rect 133509 1955 133567 1961
rect 133509 1952 133521 1955
rect 133472 1924 133521 1952
rect 133472 1912 133478 1924
rect 133509 1921 133521 1924
rect 133555 1952 133567 1955
rect 134334 1952 134340 1964
rect 133555 1924 134340 1952
rect 133555 1921 133567 1924
rect 133509 1915 133567 1921
rect 134334 1912 134340 1924
rect 134392 1912 134398 1964
rect 135346 1912 135352 1964
rect 135404 1912 135410 1964
rect 138477 1955 138535 1961
rect 138477 1921 138489 1955
rect 138523 1952 138535 1955
rect 139026 1952 139032 1964
rect 138523 1924 139032 1952
rect 138523 1921 138535 1924
rect 138477 1915 138535 1921
rect 139026 1912 139032 1924
rect 139084 1912 139090 1964
rect 139136 1961 139164 1992
rect 140222 1980 140228 1992
rect 140280 1980 140286 2032
rect 139121 1955 139179 1961
rect 139121 1921 139133 1955
rect 139167 1921 139179 1955
rect 139121 1915 139179 1921
rect 139762 1912 139768 1964
rect 139820 1912 139826 1964
rect 140498 1912 140504 1964
rect 140556 1912 140562 1964
rect 140700 1952 140728 2060
rect 140866 2048 140872 2100
rect 140924 2088 140930 2100
rect 141694 2088 141700 2100
rect 140924 2060 141700 2088
rect 140924 2048 140930 2060
rect 141694 2048 141700 2060
rect 141752 2048 141758 2100
rect 142338 2048 142344 2100
rect 142396 2048 142402 2100
rect 144638 2048 144644 2100
rect 144696 2048 144702 2100
rect 145742 2048 145748 2100
rect 145800 2088 145806 2100
rect 145800 2060 147352 2088
rect 145800 2048 145806 2060
rect 147324 2020 147352 2060
rect 147398 2048 147404 2100
rect 147456 2088 147462 2100
rect 147493 2091 147551 2097
rect 147493 2088 147505 2091
rect 147456 2060 147505 2088
rect 147456 2048 147462 2060
rect 147493 2057 147505 2060
rect 147539 2057 147551 2091
rect 147493 2051 147551 2057
rect 148594 2048 148600 2100
rect 148652 2088 148658 2100
rect 149793 2091 149851 2097
rect 149793 2088 149805 2091
rect 148652 2060 149805 2088
rect 148652 2048 148658 2060
rect 149793 2057 149805 2060
rect 149839 2057 149851 2091
rect 149793 2051 149851 2057
rect 152090 2048 152096 2100
rect 152148 2088 152154 2100
rect 152148 2060 152504 2088
rect 152148 2048 152154 2060
rect 152476 2020 152504 2060
rect 152550 2048 152556 2100
rect 152608 2088 152614 2100
rect 152645 2091 152703 2097
rect 152645 2088 152657 2091
rect 152608 2060 152657 2088
rect 152608 2048 152614 2060
rect 152645 2057 152657 2060
rect 152691 2057 152703 2091
rect 152645 2051 152703 2057
rect 152734 2048 152740 2100
rect 152792 2088 152798 2100
rect 153105 2091 153163 2097
rect 153105 2088 153117 2091
rect 152792 2060 153117 2088
rect 152792 2048 152798 2060
rect 153105 2057 153117 2060
rect 153151 2057 153163 2091
rect 153105 2051 153163 2057
rect 153749 2091 153807 2097
rect 153749 2057 153761 2091
rect 153795 2088 153807 2091
rect 153838 2088 153844 2100
rect 153795 2060 153844 2088
rect 153795 2057 153807 2060
rect 153749 2051 153807 2057
rect 153838 2048 153844 2060
rect 153896 2048 153902 2100
rect 153930 2048 153936 2100
rect 153988 2088 153994 2100
rect 154393 2091 154451 2097
rect 154393 2088 154405 2091
rect 153988 2060 154405 2088
rect 153988 2048 153994 2060
rect 154393 2057 154405 2060
rect 154439 2057 154451 2091
rect 154393 2051 154451 2057
rect 154942 2048 154948 2100
rect 155000 2088 155006 2100
rect 155037 2091 155095 2097
rect 155037 2088 155049 2091
rect 155000 2060 155049 2088
rect 155000 2048 155006 2060
rect 155037 2057 155049 2060
rect 155083 2057 155095 2091
rect 155037 2051 155095 2057
rect 159082 2048 159088 2100
rect 159140 2088 159146 2100
rect 159453 2091 159511 2097
rect 159453 2088 159465 2091
rect 159140 2060 159465 2088
rect 159140 2048 159146 2060
rect 159453 2057 159465 2060
rect 159499 2057 159511 2091
rect 160186 2088 160192 2100
rect 159453 2051 159511 2057
rect 160020 2060 160192 2088
rect 147324 1992 147674 2020
rect 152476 1992 155264 2020
rect 140700 1924 140820 1952
rect 129700 1856 132448 1884
rect 129700 1844 129706 1856
rect 134150 1844 134156 1896
rect 134208 1844 134214 1896
rect 140685 1887 140743 1893
rect 140685 1884 140697 1887
rect 138952 1856 140697 1884
rect 138952 1825 138980 1856
rect 140685 1853 140697 1856
rect 140731 1853 140743 1887
rect 140792 1884 140820 1924
rect 141418 1912 141424 1964
rect 141476 1912 141482 1964
rect 141694 1912 141700 1964
rect 141752 1912 141758 1964
rect 142798 1912 142804 1964
rect 142856 1912 142862 1964
rect 143718 1912 143724 1964
rect 143776 1912 143782 1964
rect 143902 1961 143908 1964
rect 143859 1955 143908 1961
rect 143859 1921 143871 1955
rect 143905 1921 143908 1955
rect 143859 1915 143908 1921
rect 143902 1912 143908 1915
rect 143960 1912 143966 1964
rect 145190 1912 145196 1964
rect 145248 1952 145254 1964
rect 145653 1955 145711 1961
rect 145653 1952 145665 1955
rect 145248 1924 145665 1952
rect 145248 1912 145254 1924
rect 145653 1921 145665 1924
rect 145699 1921 145711 1955
rect 145653 1915 145711 1921
rect 146570 1912 146576 1964
rect 146628 1912 146634 1964
rect 147646 1952 147674 1992
rect 147953 1955 148011 1961
rect 147953 1952 147965 1955
rect 147646 1924 147965 1952
rect 147953 1921 147965 1924
rect 147999 1921 148011 1955
rect 147953 1915 148011 1921
rect 150618 1912 150624 1964
rect 150676 1952 150682 1964
rect 150805 1955 150863 1961
rect 150805 1952 150817 1955
rect 150676 1924 150817 1952
rect 150676 1912 150682 1924
rect 150805 1921 150817 1924
rect 150851 1921 150863 1955
rect 150805 1915 150863 1921
rect 151722 1912 151728 1964
rect 151780 1912 151786 1964
rect 151998 1912 152004 1964
rect 152056 1912 152062 1964
rect 153286 1912 153292 1964
rect 153344 1912 153350 1964
rect 153378 1912 153384 1964
rect 153436 1952 153442 1964
rect 153933 1955 153991 1961
rect 153933 1952 153945 1955
rect 153436 1924 153945 1952
rect 153436 1912 153442 1924
rect 153933 1921 153945 1924
rect 153979 1921 153991 1955
rect 153933 1915 153991 1921
rect 154574 1912 154580 1964
rect 154632 1912 154638 1964
rect 155236 1961 155264 1992
rect 157334 1980 157340 2032
rect 157392 2020 157398 2032
rect 158349 2023 158407 2029
rect 158349 2020 158361 2023
rect 157392 1992 158361 2020
rect 157392 1980 157398 1992
rect 158349 1989 158361 1992
rect 158395 2020 158407 2023
rect 158530 2020 158536 2032
rect 158395 1992 158536 2020
rect 158395 1989 158407 1992
rect 158349 1983 158407 1989
rect 158530 1980 158536 1992
rect 158588 1980 158594 2032
rect 160020 2020 160048 2060
rect 160186 2048 160192 2060
rect 160244 2048 160250 2100
rect 160278 2048 160284 2100
rect 160336 2048 160342 2100
rect 161474 2048 161480 2100
rect 161532 2088 161538 2100
rect 162305 2091 162363 2097
rect 162305 2088 162317 2091
rect 161532 2060 162317 2088
rect 161532 2048 161538 2060
rect 162305 2057 162317 2060
rect 162351 2057 162363 2091
rect 162305 2051 162363 2057
rect 163958 2048 163964 2100
rect 164016 2048 164022 2100
rect 165614 2048 165620 2100
rect 165672 2048 165678 2100
rect 165798 2048 165804 2100
rect 165856 2088 165862 2100
rect 166629 2091 166687 2097
rect 166629 2088 166641 2091
rect 165856 2060 166641 2088
rect 165856 2048 165862 2060
rect 166629 2057 166641 2060
rect 166675 2057 166687 2091
rect 166629 2051 166687 2057
rect 167454 2048 167460 2100
rect 167512 2048 167518 2100
rect 190914 2048 190920 2100
rect 190972 2048 190978 2100
rect 192202 2048 192208 2100
rect 192260 2048 192266 2100
rect 192312 2060 197492 2088
rect 162394 2020 162400 2032
rect 158916 1992 160048 2020
rect 160112 1992 162400 2020
rect 155221 1955 155279 1961
rect 155221 1921 155233 1955
rect 155267 1921 155279 1955
rect 155221 1915 155279 1921
rect 155773 1955 155831 1961
rect 155773 1921 155785 1955
rect 155819 1952 155831 1955
rect 156322 1952 156328 1964
rect 155819 1924 156328 1952
rect 155819 1921 155831 1924
rect 155773 1915 155831 1921
rect 156322 1912 156328 1924
rect 156380 1912 156386 1964
rect 156417 1955 156475 1961
rect 156417 1921 156429 1955
rect 156463 1952 156475 1955
rect 156782 1952 156788 1964
rect 156463 1924 156788 1952
rect 156463 1921 156475 1924
rect 156417 1915 156475 1921
rect 156782 1912 156788 1924
rect 156840 1912 156846 1964
rect 157981 1955 158039 1961
rect 157981 1921 157993 1955
rect 158027 1952 158039 1955
rect 158916 1952 158944 1992
rect 158027 1924 158944 1952
rect 158027 1921 158039 1924
rect 157981 1915 158039 1921
rect 158990 1912 158996 1964
rect 159048 1952 159054 1964
rect 159085 1955 159143 1961
rect 159085 1952 159097 1955
rect 159048 1924 159097 1952
rect 159048 1912 159054 1924
rect 159085 1921 159097 1924
rect 159131 1921 159143 1955
rect 159085 1915 159143 1921
rect 159266 1912 159272 1964
rect 159324 1952 159330 1964
rect 160002 1952 160008 1964
rect 159324 1924 160008 1952
rect 159324 1912 159330 1924
rect 160002 1912 160008 1924
rect 160060 1952 160066 1964
rect 160112 1961 160140 1992
rect 160097 1955 160155 1961
rect 160097 1952 160109 1955
rect 160060 1924 160109 1952
rect 160060 1912 160066 1924
rect 160097 1921 160109 1924
rect 160143 1921 160155 1955
rect 160097 1915 160155 1921
rect 161106 1912 161112 1964
rect 161164 1912 161170 1964
rect 161308 1961 161336 1992
rect 161293 1955 161351 1961
rect 161293 1921 161305 1955
rect 161339 1921 161351 1955
rect 161293 1915 161351 1921
rect 161566 1912 161572 1964
rect 161624 1952 161630 1964
rect 162136 1961 162164 1992
rect 162394 1980 162400 1992
rect 162452 2020 162458 2032
rect 167178 2020 167184 2032
rect 162452 1992 162992 2020
rect 162452 1980 162458 1992
rect 161937 1955 161995 1961
rect 161937 1952 161949 1955
rect 161624 1924 161949 1952
rect 161624 1912 161630 1924
rect 161937 1921 161949 1924
rect 161983 1921 161995 1955
rect 161937 1915 161995 1921
rect 162121 1955 162179 1961
rect 162121 1921 162133 1955
rect 162167 1921 162179 1955
rect 162121 1915 162179 1921
rect 162670 1912 162676 1964
rect 162728 1952 162734 1964
rect 162964 1961 162992 1992
rect 166966 1992 167184 2020
rect 162765 1955 162823 1961
rect 162765 1952 162777 1955
rect 162728 1924 162777 1952
rect 162728 1912 162734 1924
rect 162765 1921 162777 1924
rect 162811 1921 162823 1955
rect 162765 1915 162823 1921
rect 162949 1955 163007 1961
rect 162949 1921 162961 1955
rect 162995 1921 163007 1955
rect 162949 1915 163007 1921
rect 163590 1912 163596 1964
rect 163648 1912 163654 1964
rect 163777 1955 163835 1961
rect 163777 1921 163789 1955
rect 163823 1921 163835 1955
rect 163777 1915 163835 1921
rect 141050 1884 141056 1896
rect 140792 1856 141056 1884
rect 140685 1847 140743 1853
rect 141050 1844 141056 1856
rect 141108 1884 141114 1896
rect 141602 1893 141608 1896
rect 141145 1887 141203 1893
rect 141145 1884 141157 1887
rect 141108 1856 141157 1884
rect 141108 1844 141114 1856
rect 141145 1853 141157 1856
rect 141191 1853 141203 1887
rect 141145 1847 141203 1853
rect 141559 1887 141608 1893
rect 141559 1853 141571 1887
rect 141605 1853 141608 1887
rect 141559 1847 141608 1853
rect 141602 1844 141608 1847
rect 141660 1844 141666 1896
rect 142985 1887 143043 1893
rect 142985 1853 142997 1887
rect 143031 1853 143043 1887
rect 142985 1847 143043 1853
rect 143997 1887 144055 1893
rect 143997 1853 144009 1887
rect 144043 1884 144055 1887
rect 144178 1884 144184 1896
rect 144043 1856 144184 1884
rect 144043 1853 144055 1856
rect 143997 1847 144055 1853
rect 138937 1819 138995 1825
rect 138937 1785 138949 1819
rect 138983 1785 138995 1819
rect 138937 1779 138995 1785
rect 139026 1776 139032 1828
rect 139084 1816 139090 1828
rect 139084 1788 140728 1816
rect 139084 1776 139090 1788
rect 140700 1760 140728 1788
rect 118200 1720 118280 1748
rect 118200 1708 118206 1720
rect 118602 1708 118608 1760
rect 118660 1748 118666 1760
rect 119893 1751 119951 1757
rect 119893 1748 119905 1751
rect 118660 1720 119905 1748
rect 118660 1708 118666 1720
rect 119893 1717 119905 1720
rect 119939 1717 119951 1751
rect 119893 1711 119951 1717
rect 120534 1708 120540 1760
rect 120592 1708 120598 1760
rect 121638 1708 121644 1760
rect 121696 1748 121702 1760
rect 121825 1751 121883 1757
rect 121825 1748 121837 1751
rect 121696 1720 121837 1748
rect 121696 1708 121702 1720
rect 121825 1717 121837 1720
rect 121871 1717 121883 1751
rect 121825 1711 121883 1717
rect 122466 1708 122472 1760
rect 122524 1708 122530 1760
rect 123202 1708 123208 1760
rect 123260 1748 123266 1760
rect 123481 1751 123539 1757
rect 123481 1748 123493 1751
rect 123260 1720 123493 1748
rect 123260 1708 123266 1720
rect 123481 1717 123493 1720
rect 123527 1717 123539 1751
rect 123481 1711 123539 1717
rect 125778 1708 125784 1760
rect 125836 1708 125842 1760
rect 127529 1751 127587 1757
rect 127529 1717 127541 1751
rect 127575 1748 127587 1751
rect 127618 1748 127624 1760
rect 127575 1720 127624 1748
rect 127575 1717 127587 1720
rect 127529 1711 127587 1717
rect 127618 1708 127624 1720
rect 127676 1708 127682 1760
rect 130654 1708 130660 1760
rect 130712 1748 130718 1760
rect 130841 1751 130899 1757
rect 130841 1748 130853 1751
rect 130712 1720 130853 1748
rect 130712 1708 130718 1720
rect 130841 1717 130853 1720
rect 130887 1717 130899 1751
rect 130841 1711 130899 1717
rect 132678 1708 132684 1760
rect 132736 1708 132742 1760
rect 134334 1708 134340 1760
rect 134392 1748 134398 1760
rect 134521 1751 134579 1757
rect 134521 1748 134533 1751
rect 134392 1720 134533 1748
rect 134392 1708 134398 1720
rect 134521 1717 134533 1720
rect 134567 1717 134579 1751
rect 134521 1711 134579 1717
rect 135254 1708 135260 1760
rect 135312 1748 135318 1760
rect 135533 1751 135591 1757
rect 135533 1748 135545 1751
rect 135312 1720 135545 1748
rect 135312 1708 135318 1720
rect 135533 1717 135545 1720
rect 135579 1717 135591 1751
rect 135533 1711 135591 1717
rect 138293 1751 138351 1757
rect 138293 1717 138305 1751
rect 138339 1748 138351 1751
rect 140222 1748 140228 1760
rect 138339 1720 140228 1748
rect 138339 1717 138351 1720
rect 138293 1711 138351 1717
rect 140222 1708 140228 1720
rect 140280 1708 140286 1760
rect 140682 1708 140688 1760
rect 140740 1708 140746 1760
rect 140866 1708 140872 1760
rect 140924 1748 140930 1760
rect 142430 1748 142436 1760
rect 140924 1720 142436 1748
rect 140924 1708 140930 1720
rect 142430 1708 142436 1720
rect 142488 1708 142494 1760
rect 143000 1748 143028 1847
rect 144178 1844 144184 1856
rect 144236 1844 144242 1896
rect 145837 1887 145895 1893
rect 145837 1853 145849 1887
rect 145883 1884 145895 1887
rect 146386 1884 146392 1896
rect 145883 1856 146392 1884
rect 145883 1853 145895 1856
rect 145837 1847 145895 1853
rect 146386 1844 146392 1856
rect 146444 1844 146450 1896
rect 146662 1844 146668 1896
rect 146720 1893 146726 1896
rect 146720 1887 146769 1893
rect 146720 1853 146723 1887
rect 146757 1853 146769 1887
rect 146720 1847 146769 1853
rect 146720 1844 146726 1847
rect 146846 1844 146852 1896
rect 146904 1844 146910 1896
rect 148137 1887 148195 1893
rect 148137 1853 148149 1887
rect 148183 1853 148195 1887
rect 148137 1847 148195 1853
rect 143442 1776 143448 1828
rect 143500 1776 143506 1828
rect 146294 1776 146300 1828
rect 146352 1776 146358 1828
rect 144822 1748 144828 1760
rect 143000 1720 144828 1748
rect 144822 1708 144828 1720
rect 144880 1708 144886 1760
rect 148152 1748 148180 1847
rect 148502 1844 148508 1896
rect 148560 1884 148566 1896
rect 148597 1887 148655 1893
rect 148597 1884 148609 1887
rect 148560 1856 148609 1884
rect 148560 1844 148566 1856
rect 148597 1853 148609 1856
rect 148643 1853 148655 1887
rect 148597 1847 148655 1853
rect 148686 1844 148692 1896
rect 148744 1884 148750 1896
rect 148873 1887 148931 1893
rect 148873 1884 148885 1887
rect 148744 1856 148885 1884
rect 148744 1844 148750 1856
rect 148873 1853 148885 1856
rect 148919 1853 148931 1887
rect 148873 1847 148931 1853
rect 148962 1844 148968 1896
rect 149020 1893 149026 1896
rect 149020 1887 149048 1893
rect 149036 1853 149048 1887
rect 149020 1847 149048 1853
rect 149149 1887 149207 1893
rect 149149 1853 149161 1887
rect 149195 1884 149207 1887
rect 149330 1884 149336 1896
rect 149195 1856 149336 1884
rect 149195 1853 149207 1856
rect 149149 1847 149207 1853
rect 149020 1844 149026 1847
rect 149330 1844 149336 1856
rect 149388 1884 149394 1896
rect 149698 1884 149704 1896
rect 149388 1856 149704 1884
rect 149388 1844 149394 1856
rect 149698 1844 149704 1856
rect 149756 1844 149762 1896
rect 150989 1887 151047 1893
rect 150989 1853 151001 1887
rect 151035 1884 151047 1887
rect 151538 1884 151544 1896
rect 151035 1856 151544 1884
rect 151035 1853 151047 1856
rect 150989 1847 151047 1853
rect 151538 1844 151544 1856
rect 151596 1844 151602 1896
rect 151863 1887 151921 1893
rect 151863 1853 151875 1887
rect 151909 1884 151921 1887
rect 151909 1856 154436 1884
rect 151909 1853 151921 1856
rect 151863 1847 151921 1853
rect 150618 1776 150624 1828
rect 150676 1816 150682 1828
rect 150676 1788 151400 1816
rect 150676 1776 150682 1788
rect 151262 1748 151268 1760
rect 148152 1720 151268 1748
rect 151262 1708 151268 1720
rect 151320 1708 151326 1760
rect 151372 1748 151400 1788
rect 151446 1776 151452 1828
rect 151504 1776 151510 1828
rect 154408 1816 154436 1856
rect 154592 1856 154804 1884
rect 154592 1816 154620 1856
rect 154408 1788 154620 1816
rect 154776 1816 154804 1856
rect 156598 1844 156604 1896
rect 156656 1884 156662 1896
rect 157061 1887 157119 1893
rect 157061 1884 157073 1887
rect 156656 1856 157073 1884
rect 156656 1844 156662 1856
rect 157061 1853 157073 1856
rect 157107 1884 157119 1887
rect 157150 1884 157156 1896
rect 157107 1856 157156 1884
rect 157107 1853 157119 1856
rect 157061 1847 157119 1853
rect 157150 1844 157156 1856
rect 157208 1844 157214 1896
rect 159174 1844 159180 1896
rect 159232 1884 159238 1896
rect 159913 1887 159971 1893
rect 159913 1884 159925 1887
rect 159232 1856 159925 1884
rect 159232 1844 159238 1856
rect 159913 1853 159925 1856
rect 159959 1853 159971 1887
rect 159913 1847 159971 1853
rect 162854 1844 162860 1896
rect 162912 1884 162918 1896
rect 163792 1884 163820 1915
rect 164510 1912 164516 1964
rect 164568 1912 164574 1964
rect 164605 1955 164663 1961
rect 164605 1921 164617 1955
rect 164651 1921 164663 1955
rect 164605 1915 164663 1921
rect 164620 1884 164648 1915
rect 165154 1912 165160 1964
rect 165212 1952 165218 1964
rect 165249 1955 165307 1961
rect 165249 1952 165261 1955
rect 165212 1924 165261 1952
rect 165212 1912 165218 1924
rect 165249 1921 165261 1924
rect 165295 1921 165307 1955
rect 165249 1915 165307 1921
rect 165433 1955 165491 1961
rect 165433 1921 165445 1955
rect 165479 1921 165491 1955
rect 165433 1915 165491 1921
rect 165448 1884 165476 1915
rect 166258 1912 166264 1964
rect 166316 1912 166322 1964
rect 166445 1955 166503 1961
rect 166445 1921 166457 1955
rect 166491 1952 166503 1955
rect 166966 1952 166994 1992
rect 167178 1980 167184 1992
rect 167236 2020 167242 2032
rect 167236 1992 167316 2020
rect 167236 1980 167242 1992
rect 166491 1924 166994 1952
rect 166491 1921 166503 1924
rect 166445 1915 166503 1921
rect 166460 1884 166488 1915
rect 167086 1912 167092 1964
rect 167144 1912 167150 1964
rect 167288 1961 167316 1992
rect 173802 1980 173808 2032
rect 173860 2020 173866 2032
rect 173860 1992 180794 2020
rect 173860 1980 173866 1992
rect 167273 1955 167331 1961
rect 167273 1921 167285 1955
rect 167319 1952 167331 1955
rect 168006 1952 168012 1964
rect 167319 1924 168012 1952
rect 167319 1921 167331 1924
rect 167273 1915 167331 1921
rect 168006 1912 168012 1924
rect 168064 1952 168070 1964
rect 168101 1955 168159 1961
rect 168101 1952 168113 1955
rect 168064 1924 168113 1952
rect 168064 1912 168070 1924
rect 168101 1921 168113 1924
rect 168147 1921 168159 1955
rect 168101 1915 168159 1921
rect 168285 1955 168343 1961
rect 168285 1921 168297 1955
rect 168331 1952 168343 1955
rect 168745 1955 168803 1961
rect 168745 1952 168757 1955
rect 168331 1924 168757 1952
rect 168331 1921 168343 1924
rect 168285 1915 168343 1921
rect 168745 1921 168757 1924
rect 168791 1921 168803 1955
rect 168745 1915 168803 1921
rect 169754 1912 169760 1964
rect 169812 1952 169818 1964
rect 173253 1955 173311 1961
rect 173253 1952 173265 1955
rect 169812 1924 173265 1952
rect 169812 1912 169818 1924
rect 173253 1921 173265 1924
rect 173299 1921 173311 1955
rect 173253 1915 173311 1921
rect 176838 1912 176844 1964
rect 176896 1912 176902 1964
rect 179414 1912 179420 1964
rect 179472 1912 179478 1964
rect 180766 1952 180794 1992
rect 182082 1980 182088 2032
rect 182140 2020 182146 2032
rect 190638 2020 190644 2032
rect 182140 1992 188476 2020
rect 182140 1980 182146 1992
rect 183281 1955 183339 1961
rect 183281 1952 183293 1955
rect 180766 1924 183293 1952
rect 183281 1921 183293 1924
rect 183327 1921 183339 1955
rect 183281 1915 183339 1921
rect 184566 1912 184572 1964
rect 184624 1912 184630 1964
rect 187142 1912 187148 1964
rect 187200 1912 187206 1964
rect 188448 1961 188476 1992
rect 190426 1992 190644 2020
rect 188433 1955 188491 1961
rect 188433 1921 188445 1955
rect 188479 1921 188491 1955
rect 188433 1915 188491 1921
rect 190273 1955 190331 1961
rect 190273 1921 190285 1955
rect 190319 1952 190331 1955
rect 190426 1952 190454 1992
rect 190638 1980 190644 1992
rect 190696 2020 190702 2032
rect 192312 2020 192340 2060
rect 196434 2020 196440 2032
rect 190696 1992 192340 2020
rect 194704 1992 196440 2020
rect 190696 1980 190702 1992
rect 190549 1955 190607 1961
rect 190549 1952 190561 1955
rect 190319 1924 190561 1952
rect 190319 1921 190331 1924
rect 190273 1915 190331 1921
rect 190549 1921 190561 1924
rect 190595 1921 190607 1955
rect 190549 1915 190607 1921
rect 190733 1955 190791 1961
rect 190733 1921 190745 1955
rect 190779 1952 190791 1955
rect 191006 1952 191012 1964
rect 190779 1924 191012 1952
rect 190779 1921 190791 1924
rect 190733 1915 190791 1921
rect 191006 1912 191012 1924
rect 191064 1952 191070 1964
rect 192021 1955 192079 1961
rect 192021 1952 192033 1955
rect 191064 1924 192033 1952
rect 191064 1912 191070 1924
rect 192021 1921 192033 1924
rect 192067 1952 192079 1955
rect 193033 1955 193091 1961
rect 193033 1952 193045 1955
rect 192067 1924 193045 1952
rect 192067 1921 192079 1924
rect 192021 1915 192079 1921
rect 193033 1921 193045 1924
rect 193079 1921 193091 1955
rect 193033 1915 193091 1921
rect 162912 1856 166488 1884
rect 162912 1844 162918 1856
rect 166534 1844 166540 1896
rect 166592 1884 166598 1896
rect 167822 1884 167828 1896
rect 166592 1856 167828 1884
rect 166592 1844 166598 1856
rect 167822 1844 167828 1856
rect 167880 1884 167886 1896
rect 167917 1887 167975 1893
rect 167917 1884 167929 1887
rect 167880 1856 167929 1884
rect 167880 1844 167886 1856
rect 167917 1853 167929 1856
rect 167963 1853 167975 1887
rect 167917 1847 167975 1853
rect 172974 1844 172980 1896
rect 173032 1844 173038 1896
rect 174446 1844 174452 1896
rect 174504 1844 174510 1896
rect 174722 1844 174728 1896
rect 174780 1844 174786 1896
rect 176562 1844 176568 1896
rect 176620 1844 176626 1896
rect 177850 1844 177856 1896
rect 177908 1844 177914 1896
rect 178126 1844 178132 1896
rect 178184 1844 178190 1896
rect 179138 1844 179144 1896
rect 179196 1844 179202 1896
rect 181714 1844 181720 1896
rect 181772 1844 181778 1896
rect 181993 1887 182051 1893
rect 181993 1853 182005 1887
rect 182039 1853 182051 1887
rect 181993 1847 182051 1853
rect 182008 1816 182036 1847
rect 183002 1844 183008 1896
rect 183060 1844 183066 1896
rect 184290 1844 184296 1896
rect 184348 1844 184354 1896
rect 186314 1844 186320 1896
rect 186372 1884 186378 1896
rect 186869 1887 186927 1893
rect 186869 1884 186881 1887
rect 186372 1856 186881 1884
rect 186372 1844 186378 1856
rect 186869 1853 186881 1856
rect 186915 1853 186927 1887
rect 186869 1847 186927 1853
rect 188154 1844 188160 1896
rect 188212 1844 188218 1896
rect 191834 1844 191840 1896
rect 191892 1844 191898 1896
rect 192573 1887 192631 1893
rect 192573 1853 192585 1887
rect 192619 1884 192631 1887
rect 192846 1884 192852 1896
rect 192619 1856 192852 1884
rect 192619 1853 192631 1856
rect 192573 1847 192631 1853
rect 192846 1844 192852 1856
rect 192904 1844 192910 1896
rect 193048 1884 193076 1915
rect 193490 1912 193496 1964
rect 193548 1952 193554 1964
rect 194704 1961 194732 1992
rect 193677 1955 193735 1961
rect 193677 1952 193689 1955
rect 193548 1924 193689 1952
rect 193548 1912 193554 1924
rect 193677 1921 193689 1924
rect 193723 1921 193735 1955
rect 193677 1915 193735 1921
rect 193861 1955 193919 1961
rect 193861 1921 193873 1955
rect 193907 1952 193919 1955
rect 194689 1955 194747 1961
rect 194689 1952 194701 1955
rect 193907 1924 194701 1952
rect 193907 1921 193919 1924
rect 193861 1915 193919 1921
rect 194689 1921 194701 1924
rect 194735 1921 194747 1955
rect 194689 1915 194747 1921
rect 193876 1884 193904 1915
rect 195330 1912 195336 1964
rect 195388 1912 195394 1964
rect 195532 1961 195560 1992
rect 195517 1955 195575 1961
rect 195517 1921 195529 1955
rect 195563 1921 195575 1955
rect 195517 1915 195575 1921
rect 195698 1912 195704 1964
rect 195756 1912 195762 1964
rect 195974 1912 195980 1964
rect 196032 1952 196038 1964
rect 196360 1961 196388 1992
rect 196434 1980 196440 1992
rect 196492 2020 196498 2032
rect 197464 2020 197492 2060
rect 197538 2048 197544 2100
rect 197596 2048 197602 2100
rect 199746 2048 199752 2100
rect 199804 2048 199810 2100
rect 216582 2088 216588 2100
rect 200086 2060 216588 2088
rect 200086 2020 200114 2060
rect 216582 2048 216588 2060
rect 216640 2048 216646 2100
rect 216674 2048 216680 2100
rect 216732 2088 216738 2100
rect 216769 2091 216827 2097
rect 216769 2088 216781 2091
rect 216732 2060 216781 2088
rect 216732 2048 216738 2060
rect 216769 2057 216781 2060
rect 216815 2057 216827 2091
rect 216769 2051 216827 2057
rect 218422 2048 218428 2100
rect 218480 2088 218486 2100
rect 218480 2060 219572 2088
rect 218480 2048 218486 2060
rect 196492 1992 197400 2020
rect 197464 1992 200114 2020
rect 196492 1980 196498 1992
rect 196161 1955 196219 1961
rect 196161 1952 196173 1955
rect 196032 1924 196173 1952
rect 196032 1912 196038 1924
rect 196161 1921 196173 1924
rect 196207 1921 196219 1955
rect 196161 1915 196219 1921
rect 196345 1955 196403 1961
rect 196345 1921 196357 1955
rect 196391 1921 196403 1955
rect 196345 1915 196403 1921
rect 197170 1912 197176 1964
rect 197228 1912 197234 1964
rect 197372 1961 197400 1992
rect 200206 1980 200212 2032
rect 200264 2020 200270 2032
rect 201405 2023 201463 2029
rect 201405 2020 201417 2023
rect 200264 1992 201417 2020
rect 200264 1980 200270 1992
rect 201405 1989 201417 1992
rect 201451 1989 201463 2023
rect 201405 1983 201463 1989
rect 202690 1980 202696 2032
rect 202748 1980 202754 2032
rect 209682 2020 209688 2032
rect 207860 1992 209688 2020
rect 197357 1955 197415 1961
rect 197357 1921 197369 1955
rect 197403 1921 197415 1955
rect 197357 1915 197415 1921
rect 199378 1912 199384 1964
rect 199436 1912 199442 1964
rect 199565 1955 199623 1961
rect 199565 1921 199577 1955
rect 199611 1952 199623 1955
rect 199611 1924 200114 1952
rect 199611 1921 199623 1924
rect 199565 1915 199623 1921
rect 193048 1856 193904 1884
rect 194505 1887 194563 1893
rect 194505 1853 194517 1887
rect 194551 1884 194563 1887
rect 194778 1884 194784 1896
rect 194551 1856 194784 1884
rect 194551 1853 194563 1856
rect 194505 1847 194563 1853
rect 194778 1844 194784 1856
rect 194836 1844 194842 1896
rect 198093 1887 198151 1893
rect 198093 1853 198105 1887
rect 198139 1853 198151 1887
rect 198093 1847 198151 1853
rect 154776 1788 182036 1816
rect 191190 1776 191196 1828
rect 191248 1816 191254 1828
rect 198108 1816 198136 1847
rect 198366 1844 198372 1896
rect 198424 1884 198430 1896
rect 199580 1884 199608 1915
rect 198424 1856 199608 1884
rect 200086 1884 200114 1924
rect 200298 1912 200304 1964
rect 200356 1912 200362 1964
rect 200393 1955 200451 1961
rect 200393 1921 200405 1955
rect 200439 1921 200451 1955
rect 200393 1915 200451 1921
rect 200408 1884 200436 1915
rect 200666 1912 200672 1964
rect 200724 1952 200730 1964
rect 201037 1955 201095 1961
rect 201037 1952 201049 1955
rect 200724 1924 201049 1952
rect 200724 1912 200730 1924
rect 201037 1921 201049 1924
rect 201083 1921 201095 1955
rect 201037 1915 201095 1921
rect 201221 1955 201279 1961
rect 201221 1921 201233 1955
rect 201267 1921 201279 1955
rect 201221 1915 201279 1921
rect 201236 1884 201264 1915
rect 202322 1912 202328 1964
rect 202380 1912 202386 1964
rect 202509 1955 202567 1961
rect 202509 1921 202521 1955
rect 202555 1921 202567 1955
rect 202509 1915 202567 1921
rect 201494 1884 201500 1896
rect 200086 1856 201500 1884
rect 198424 1844 198430 1856
rect 201494 1844 201500 1856
rect 201552 1884 201558 1896
rect 202524 1884 202552 1915
rect 203242 1912 203248 1964
rect 203300 1912 203306 1964
rect 207860 1961 207888 1992
rect 209682 1980 209688 1992
rect 209740 1980 209746 2032
rect 210694 1980 210700 2032
rect 210752 2020 210758 2032
rect 210752 1992 211752 2020
rect 210752 1980 210758 1992
rect 203337 1955 203395 1961
rect 203337 1921 203349 1955
rect 203383 1921 203395 1955
rect 203337 1915 203395 1921
rect 203521 1955 203579 1961
rect 203521 1921 203533 1955
rect 203567 1952 203579 1955
rect 203981 1955 204039 1961
rect 203981 1952 203993 1955
rect 203567 1924 203993 1952
rect 203567 1921 203579 1924
rect 203521 1915 203579 1921
rect 203981 1921 203993 1924
rect 204027 1921 204039 1955
rect 203981 1915 204039 1921
rect 207845 1955 207903 1961
rect 207845 1921 207857 1955
rect 207891 1921 207903 1955
rect 207845 1915 207903 1921
rect 202782 1884 202788 1896
rect 201552 1856 202788 1884
rect 201552 1844 201558 1856
rect 202782 1844 202788 1856
rect 202840 1884 202846 1896
rect 203352 1884 203380 1915
rect 208486 1912 208492 1964
rect 208544 1912 208550 1964
rect 208946 1912 208952 1964
rect 209004 1912 209010 1964
rect 211338 1912 211344 1964
rect 211396 1912 211402 1964
rect 211430 1912 211436 1964
rect 211488 1912 211494 1964
rect 211614 1912 211620 1964
rect 211672 1912 211678 1964
rect 211724 1952 211752 1992
rect 211982 1980 211988 2032
rect 212040 1980 212046 2032
rect 214466 1980 214472 2032
rect 214524 1980 214530 2032
rect 219544 2020 219572 2060
rect 219618 2048 219624 2100
rect 219676 2048 219682 2100
rect 220722 2088 220728 2100
rect 220280 2060 220728 2088
rect 220280 2020 220308 2060
rect 220722 2048 220728 2060
rect 220780 2048 220786 2100
rect 221366 2048 221372 2100
rect 221424 2088 221430 2100
rect 221921 2091 221979 2097
rect 221921 2088 221933 2091
rect 221424 2060 221933 2088
rect 221424 2048 221430 2060
rect 221921 2057 221933 2060
rect 221967 2057 221979 2091
rect 221921 2051 221979 2057
rect 222654 2048 222660 2100
rect 222712 2088 222718 2100
rect 222933 2091 222991 2097
rect 222933 2088 222945 2091
rect 222712 2060 222945 2088
rect 222712 2048 222718 2060
rect 222933 2057 222945 2060
rect 222979 2057 222991 2091
rect 222933 2051 222991 2057
rect 224126 2048 224132 2100
rect 224184 2048 224190 2100
rect 224494 2048 224500 2100
rect 224552 2048 224558 2100
rect 225782 2048 225788 2100
rect 225840 2048 225846 2100
rect 226794 2048 226800 2100
rect 226852 2048 226858 2100
rect 228450 2048 228456 2100
rect 228508 2048 228514 2100
rect 230934 2048 230940 2100
rect 230992 2048 230998 2100
rect 231762 2048 231768 2100
rect 231820 2048 231826 2100
rect 232590 2048 232596 2100
rect 232648 2048 232654 2100
rect 232958 2048 232964 2100
rect 233016 2088 233022 2100
rect 233605 2091 233663 2097
rect 233605 2088 233617 2091
rect 233016 2060 233617 2088
rect 233016 2048 233022 2060
rect 233605 2057 233617 2060
rect 233651 2057 233663 2091
rect 233605 2051 233663 2057
rect 234982 2048 234988 2100
rect 235040 2088 235046 2100
rect 236089 2091 236147 2097
rect 236089 2088 236101 2091
rect 235040 2060 236101 2088
rect 235040 2048 235046 2060
rect 236089 2057 236101 2060
rect 236135 2057 236147 2091
rect 236089 2051 236147 2057
rect 236914 2048 236920 2100
rect 236972 2048 236978 2100
rect 237006 2048 237012 2100
rect 237064 2088 237070 2100
rect 237064 2060 238754 2088
rect 237064 2048 237070 2060
rect 214576 1992 215064 2020
rect 219544 1992 220308 2020
rect 212629 1955 212687 1961
rect 212629 1952 212641 1955
rect 211724 1924 212641 1952
rect 212629 1921 212641 1924
rect 212675 1921 212687 1955
rect 212629 1915 212687 1921
rect 213638 1912 213644 1964
rect 213696 1961 213702 1964
rect 213696 1955 213724 1961
rect 213712 1921 213724 1955
rect 213696 1915 213724 1921
rect 213696 1912 213702 1915
rect 213822 1912 213828 1964
rect 213880 1912 213886 1964
rect 214576 1952 214604 1992
rect 214392 1924 214604 1952
rect 202840 1856 203380 1884
rect 202840 1844 202846 1856
rect 208302 1844 208308 1896
rect 208360 1884 208366 1896
rect 209133 1887 209191 1893
rect 209133 1884 209145 1887
rect 208360 1856 209145 1884
rect 208360 1844 208366 1856
rect 209133 1853 209145 1856
rect 209179 1853 209191 1887
rect 209133 1847 209191 1853
rect 209774 1844 209780 1896
rect 209832 1844 209838 1896
rect 212813 1887 212871 1893
rect 212813 1853 212825 1887
rect 212859 1853 212871 1887
rect 212813 1847 212871 1853
rect 213273 1887 213331 1893
rect 213273 1853 213285 1887
rect 213319 1884 213331 1887
rect 213362 1884 213368 1896
rect 213319 1856 213368 1884
rect 213319 1853 213331 1856
rect 213273 1847 213331 1853
rect 191248 1788 198136 1816
rect 207661 1819 207719 1825
rect 191248 1776 191254 1788
rect 207661 1785 207673 1819
rect 207707 1816 207719 1819
rect 212828 1816 212856 1847
rect 207707 1788 212856 1816
rect 207707 1785 207719 1788
rect 207661 1779 207719 1785
rect 213086 1776 213092 1828
rect 213144 1816 213150 1828
rect 213288 1816 213316 1847
rect 213362 1844 213368 1856
rect 213420 1844 213426 1896
rect 213549 1887 213607 1893
rect 213549 1853 213561 1887
rect 213595 1884 213607 1887
rect 214392 1884 214420 1924
rect 214650 1912 214656 1964
rect 214708 1952 214714 1964
rect 214929 1955 214987 1961
rect 214929 1952 214941 1955
rect 214708 1924 214941 1952
rect 214708 1912 214714 1924
rect 214929 1921 214941 1924
rect 214975 1921 214987 1955
rect 215036 1952 215064 1992
rect 221826 1980 221832 2032
rect 221884 2020 221890 2032
rect 226061 2023 226119 2029
rect 226061 2020 226073 2023
rect 221884 1992 226073 2020
rect 221884 1980 221890 1992
rect 226061 1989 226073 1992
rect 226107 2020 226119 2023
rect 226426 2020 226432 2032
rect 226107 1992 226432 2020
rect 226107 1989 226119 1992
rect 226061 1983 226119 1989
rect 226426 1980 226432 1992
rect 226484 1980 226490 2032
rect 228358 2020 228364 2032
rect 228192 1992 228364 2020
rect 215036 1924 215248 1952
rect 214929 1915 214987 1921
rect 215113 1887 215171 1893
rect 215113 1884 215125 1887
rect 213595 1856 214420 1884
rect 214484 1856 215125 1884
rect 213595 1853 213607 1856
rect 213549 1847 213607 1853
rect 213144 1788 213316 1816
rect 213144 1776 213150 1788
rect 154574 1748 154580 1760
rect 151372 1720 154580 1748
rect 154574 1708 154580 1720
rect 154632 1708 154638 1760
rect 155954 1708 155960 1760
rect 156012 1708 156018 1760
rect 161474 1708 161480 1760
rect 161532 1708 161538 1760
rect 163130 1708 163136 1760
rect 163188 1708 163194 1760
rect 164418 1708 164424 1760
rect 164476 1748 164482 1760
rect 164789 1751 164847 1757
rect 164789 1748 164801 1751
rect 164476 1720 164801 1748
rect 164476 1708 164482 1720
rect 164789 1717 164801 1720
rect 164835 1717 164847 1751
rect 164789 1711 164847 1717
rect 168374 1708 168380 1760
rect 168432 1748 168438 1760
rect 168929 1751 168987 1757
rect 168929 1748 168941 1751
rect 168432 1720 168941 1748
rect 168432 1708 168438 1720
rect 168929 1717 168941 1720
rect 168975 1717 168987 1751
rect 168929 1711 168987 1717
rect 193214 1708 193220 1760
rect 193272 1708 193278 1760
rect 194042 1708 194048 1760
rect 194100 1708 194106 1760
rect 194594 1708 194600 1760
rect 194652 1748 194658 1760
rect 194873 1751 194931 1757
rect 194873 1748 194885 1751
rect 194652 1720 194885 1748
rect 194652 1708 194658 1720
rect 194873 1717 194885 1720
rect 194919 1717 194931 1751
rect 194873 1711 194931 1717
rect 196066 1708 196072 1760
rect 196124 1748 196130 1760
rect 196529 1751 196587 1757
rect 196529 1748 196541 1751
rect 196124 1720 196541 1748
rect 196124 1708 196130 1720
rect 196529 1717 196541 1720
rect 196575 1717 196587 1751
rect 196529 1711 196587 1717
rect 200574 1708 200580 1760
rect 200632 1708 200638 1760
rect 202874 1708 202880 1760
rect 202932 1748 202938 1760
rect 204165 1751 204223 1757
rect 204165 1748 204177 1751
rect 202932 1720 204177 1748
rect 202932 1708 202938 1720
rect 204165 1717 204177 1720
rect 204211 1717 204223 1751
rect 204165 1711 204223 1717
rect 208305 1751 208363 1757
rect 208305 1717 208317 1751
rect 208351 1748 208363 1751
rect 210234 1748 210240 1760
rect 208351 1720 210240 1748
rect 208351 1717 208363 1720
rect 208305 1711 208363 1717
rect 210234 1708 210240 1720
rect 210292 1708 210298 1760
rect 210694 1708 210700 1760
rect 210752 1748 210758 1760
rect 213104 1748 213132 1776
rect 210752 1720 213132 1748
rect 210752 1708 210758 1720
rect 213730 1708 213736 1760
rect 213788 1748 213794 1760
rect 214484 1748 214512 1856
rect 215113 1853 215125 1856
rect 215159 1853 215171 1887
rect 215220 1884 215248 1924
rect 215846 1912 215852 1964
rect 215904 1912 215910 1964
rect 216030 1961 216036 1964
rect 215987 1955 216036 1961
rect 215987 1921 215999 1955
rect 216033 1921 216036 1955
rect 215987 1915 216036 1921
rect 216030 1912 216036 1915
rect 216088 1912 216094 1964
rect 218698 1912 218704 1964
rect 218756 1912 218762 1964
rect 218974 1912 218980 1964
rect 219032 1912 219038 1964
rect 220170 1912 220176 1964
rect 220228 1952 220234 1964
rect 220265 1955 220323 1961
rect 220265 1952 220277 1955
rect 220228 1924 220277 1952
rect 220228 1912 220234 1924
rect 220265 1921 220277 1924
rect 220311 1921 220323 1955
rect 220265 1915 220323 1921
rect 220998 1910 221004 1962
rect 221056 1961 221062 1962
rect 221056 1955 221077 1961
rect 221065 1921 221077 1955
rect 221056 1915 221077 1921
rect 221056 1910 221062 1915
rect 221274 1912 221280 1964
rect 221332 1912 221338 1964
rect 222010 1912 222016 1964
rect 222068 1952 222074 1964
rect 223117 1955 223175 1961
rect 223117 1952 223129 1955
rect 222068 1924 223129 1952
rect 222068 1912 222074 1924
rect 223117 1921 223129 1924
rect 223163 1921 223175 1955
rect 223117 1915 223175 1921
rect 223945 1955 224003 1961
rect 223945 1921 223957 1955
rect 223991 1952 224003 1955
rect 224402 1952 224408 1964
rect 223991 1924 224408 1952
rect 223991 1921 224003 1924
rect 223945 1915 224003 1921
rect 224402 1912 224408 1924
rect 224460 1952 224466 1964
rect 224957 1955 225015 1961
rect 224957 1952 224969 1955
rect 224460 1924 224969 1952
rect 224460 1912 224466 1924
rect 224957 1921 224969 1924
rect 225003 1952 225015 1955
rect 225601 1955 225659 1961
rect 225601 1952 225613 1955
rect 225003 1924 225613 1952
rect 225003 1921 225015 1924
rect 224957 1915 225015 1921
rect 225601 1921 225613 1924
rect 225647 1952 225659 1955
rect 226613 1955 226671 1961
rect 226613 1952 226625 1955
rect 225647 1924 226625 1952
rect 225647 1921 225659 1924
rect 225601 1915 225659 1921
rect 226613 1921 226625 1924
rect 226659 1921 226671 1955
rect 226613 1915 226671 1921
rect 215478 1884 215484 1896
rect 215220 1856 215484 1884
rect 215113 1847 215171 1853
rect 215478 1844 215484 1856
rect 215536 1844 215542 1896
rect 216122 1844 216128 1896
rect 216180 1844 216186 1896
rect 217781 1887 217839 1893
rect 217781 1853 217793 1887
rect 217827 1853 217839 1887
rect 217781 1847 217839 1853
rect 217965 1887 218023 1893
rect 217965 1853 217977 1887
rect 218011 1853 218023 1887
rect 217965 1847 218023 1853
rect 218839 1887 218897 1893
rect 218839 1853 218851 1887
rect 218885 1884 218897 1887
rect 219342 1884 219348 1896
rect 218885 1856 219348 1884
rect 218885 1853 218897 1856
rect 218839 1847 218897 1853
rect 215570 1776 215576 1828
rect 215628 1776 215634 1828
rect 213788 1720 214512 1748
rect 213788 1708 213794 1720
rect 214834 1708 214840 1760
rect 214892 1748 214898 1760
rect 217796 1748 217824 1847
rect 214892 1720 217824 1748
rect 217980 1748 218008 1847
rect 219342 1844 219348 1856
rect 219400 1844 219406 1896
rect 219526 1844 219532 1896
rect 219584 1884 219590 1896
rect 220081 1887 220139 1893
rect 220081 1884 220093 1887
rect 219584 1856 220093 1884
rect 219584 1844 219590 1856
rect 220081 1853 220093 1856
rect 220127 1853 220139 1887
rect 220081 1847 220139 1853
rect 220354 1844 220360 1896
rect 220412 1884 220418 1896
rect 220725 1887 220783 1893
rect 220725 1884 220737 1887
rect 220412 1856 220737 1884
rect 220412 1844 220418 1856
rect 220725 1853 220737 1856
rect 220771 1853 220783 1887
rect 220725 1847 220783 1853
rect 221118 1887 221176 1893
rect 221118 1853 221130 1887
rect 221164 1884 221176 1887
rect 221164 1856 223068 1884
rect 221164 1853 221176 1856
rect 221118 1847 221176 1853
rect 218146 1776 218152 1828
rect 218204 1816 218210 1828
rect 218425 1819 218483 1825
rect 218425 1816 218437 1819
rect 218204 1788 218437 1816
rect 218204 1776 218210 1788
rect 218425 1785 218437 1788
rect 218471 1785 218483 1819
rect 218425 1779 218483 1785
rect 219434 1776 219440 1828
rect 219492 1816 219498 1828
rect 220446 1816 220452 1828
rect 219492 1788 220452 1816
rect 219492 1776 219498 1788
rect 220446 1776 220452 1788
rect 220504 1776 220510 1828
rect 223040 1816 223068 1856
rect 223390 1844 223396 1896
rect 223448 1884 223454 1896
rect 223761 1887 223819 1893
rect 223761 1884 223773 1887
rect 223448 1856 223773 1884
rect 223448 1844 223454 1856
rect 223761 1853 223773 1856
rect 223807 1853 223819 1887
rect 223761 1847 223819 1853
rect 224494 1844 224500 1896
rect 224552 1884 224558 1896
rect 224773 1887 224831 1893
rect 224773 1884 224785 1887
rect 224552 1856 224785 1884
rect 224552 1844 224558 1856
rect 224773 1853 224785 1856
rect 224819 1853 224831 1887
rect 224773 1847 224831 1853
rect 225414 1844 225420 1896
rect 225472 1844 225478 1896
rect 226426 1844 226432 1896
rect 226484 1844 226490 1896
rect 226628 1884 226656 1915
rect 227254 1912 227260 1964
rect 227312 1912 227318 1964
rect 228192 1961 228220 1992
rect 228358 1980 228364 1992
rect 228416 1980 228422 2032
rect 229830 1980 229836 2032
rect 229888 2020 229894 2032
rect 231486 2020 231492 2032
rect 229888 1992 230060 2020
rect 229888 1980 229894 1992
rect 228177 1955 228235 1961
rect 228177 1921 228189 1955
rect 228223 1921 228235 1955
rect 228177 1915 228235 1921
rect 228269 1955 228327 1961
rect 228269 1921 228281 1955
rect 228315 1921 228327 1955
rect 228269 1915 228327 1921
rect 227070 1884 227076 1896
rect 226628 1856 227076 1884
rect 227070 1844 227076 1856
rect 227128 1884 227134 1896
rect 228284 1884 228312 1915
rect 228910 1912 228916 1964
rect 228968 1912 228974 1964
rect 229097 1955 229155 1961
rect 229097 1952 229109 1955
rect 229020 1924 229109 1952
rect 229020 1884 229048 1924
rect 229097 1921 229109 1924
rect 229143 1921 229155 1955
rect 229097 1915 229155 1921
rect 227128 1856 229048 1884
rect 229112 1884 229140 1915
rect 229738 1912 229744 1964
rect 229796 1912 229802 1964
rect 229922 1912 229928 1964
rect 229980 1912 229986 1964
rect 229940 1884 229968 1912
rect 229112 1856 229968 1884
rect 230032 1884 230060 1992
rect 230768 1992 231492 2020
rect 230768 1964 230796 1992
rect 231486 1980 231492 1992
rect 231544 2020 231550 2032
rect 231544 1992 235948 2020
rect 231544 1980 231550 1992
rect 230658 1912 230664 1964
rect 230716 1912 230722 1964
rect 230750 1912 230756 1964
rect 230808 1912 230814 1964
rect 230842 1912 230848 1964
rect 230900 1952 230906 1964
rect 231596 1961 231624 1992
rect 231397 1955 231455 1961
rect 231397 1952 231409 1955
rect 230900 1924 231409 1952
rect 230900 1912 230906 1924
rect 231397 1921 231409 1924
rect 231443 1921 231455 1955
rect 231397 1915 231455 1921
rect 231581 1955 231639 1961
rect 231581 1921 231593 1955
rect 231627 1921 231639 1955
rect 231581 1915 231639 1921
rect 232038 1912 232044 1964
rect 232096 1952 232102 1964
rect 232424 1961 232452 1992
rect 232225 1955 232283 1961
rect 232225 1952 232237 1955
rect 232096 1924 232237 1952
rect 232096 1912 232102 1924
rect 232225 1921 232237 1924
rect 232271 1921 232283 1955
rect 232225 1915 232283 1921
rect 232409 1955 232467 1961
rect 232409 1921 232421 1955
rect 232455 1921 232467 1955
rect 232409 1915 232467 1921
rect 232774 1912 232780 1964
rect 232832 1952 232838 1964
rect 233436 1961 233464 1992
rect 233237 1955 233295 1961
rect 233237 1952 233249 1955
rect 232832 1924 233249 1952
rect 232832 1912 232838 1924
rect 233237 1921 233249 1924
rect 233283 1921 233295 1955
rect 233237 1915 233295 1921
rect 233421 1955 233479 1961
rect 233421 1921 233433 1955
rect 233467 1921 233479 1955
rect 233421 1915 233479 1921
rect 233602 1912 233608 1964
rect 233660 1952 233666 1964
rect 234264 1961 234292 1992
rect 235092 1961 235120 1992
rect 234065 1955 234123 1961
rect 234065 1952 234077 1955
rect 233660 1924 234077 1952
rect 233660 1912 233666 1924
rect 234065 1921 234077 1924
rect 234111 1921 234123 1955
rect 234065 1915 234123 1921
rect 234249 1955 234307 1961
rect 234249 1921 234261 1955
rect 234295 1921 234307 1955
rect 234249 1915 234307 1921
rect 235077 1955 235135 1961
rect 235077 1921 235089 1955
rect 235123 1921 235135 1955
rect 235077 1915 235135 1921
rect 235626 1912 235632 1964
rect 235684 1952 235690 1964
rect 235920 1961 235948 1992
rect 236178 1980 236184 2032
rect 236236 2020 236242 2032
rect 236236 1992 237420 2020
rect 236236 1980 236242 1992
rect 235721 1955 235779 1961
rect 235721 1952 235733 1955
rect 235684 1924 235733 1952
rect 235684 1912 235690 1924
rect 235721 1921 235733 1924
rect 235767 1921 235779 1955
rect 235721 1915 235779 1921
rect 235905 1955 235963 1961
rect 235905 1921 235917 1955
rect 235951 1952 235963 1955
rect 235994 1952 236000 1964
rect 235951 1924 236000 1952
rect 235951 1921 235963 1924
rect 235905 1915 235963 1921
rect 235994 1912 236000 1924
rect 236052 1912 236058 1964
rect 236086 1912 236092 1964
rect 236144 1952 236150 1964
rect 237392 1961 237420 1992
rect 236549 1955 236607 1961
rect 236549 1952 236561 1955
rect 236144 1924 236561 1952
rect 236144 1912 236150 1924
rect 236549 1921 236561 1924
rect 236595 1921 236607 1955
rect 236549 1915 236607 1921
rect 236733 1955 236791 1961
rect 236733 1921 236745 1955
rect 236779 1921 236791 1955
rect 236733 1915 236791 1921
rect 237377 1955 237435 1961
rect 237377 1921 237389 1955
rect 237423 1921 237435 1955
rect 238726 1952 238754 2060
rect 239490 2048 239496 2100
rect 239548 2088 239554 2100
rect 241471 2091 241529 2097
rect 241471 2088 241483 2091
rect 239548 2060 241483 2088
rect 239548 2048 239554 2060
rect 241471 2057 241483 2060
rect 241517 2057 241529 2091
rect 241471 2051 241529 2057
rect 243630 2048 243636 2100
rect 243688 2088 243694 2100
rect 243688 2060 247540 2088
rect 243688 2048 243694 2060
rect 245013 2023 245071 2029
rect 245013 1989 245025 2023
rect 245059 2020 245071 2023
rect 245378 2020 245384 2032
rect 245059 1992 245384 2020
rect 245059 1989 245071 1992
rect 245013 1983 245071 1989
rect 245378 1980 245384 1992
rect 245436 1980 245442 2032
rect 243817 1955 243875 1961
rect 243817 1952 243829 1955
rect 238726 1924 243829 1952
rect 237377 1915 237435 1921
rect 243817 1921 243829 1924
rect 243863 1921 243875 1955
rect 243817 1915 243875 1921
rect 246224 1924 247264 1952
rect 231670 1884 231676 1896
rect 230032 1856 231676 1884
rect 227128 1844 227134 1856
rect 231670 1844 231676 1856
rect 231728 1844 231734 1896
rect 233510 1844 233516 1896
rect 233568 1884 233574 1896
rect 234893 1887 234951 1893
rect 234893 1884 234905 1887
rect 233568 1856 234905 1884
rect 233568 1844 233574 1856
rect 234893 1853 234905 1856
rect 234939 1853 234951 1887
rect 236012 1884 236040 1912
rect 236748 1884 236776 1915
rect 236012 1856 236776 1884
rect 234893 1847 234951 1853
rect 241238 1844 241244 1896
rect 241296 1844 241302 1896
rect 242802 1844 242808 1896
rect 242860 1884 242866 1896
rect 243541 1887 243599 1893
rect 243541 1884 243553 1887
rect 242860 1856 243553 1884
rect 242860 1844 242866 1856
rect 243541 1853 243553 1856
rect 243587 1853 243599 1887
rect 243541 1847 243599 1853
rect 244826 1844 244832 1896
rect 244884 1844 244890 1896
rect 245930 1844 245936 1896
rect 245988 1884 245994 1896
rect 246224 1884 246252 1924
rect 245988 1856 246252 1884
rect 245988 1844 245994 1856
rect 246666 1844 246672 1896
rect 246724 1844 246730 1896
rect 247129 1887 247187 1893
rect 247129 1853 247141 1887
rect 247175 1853 247187 1887
rect 247129 1847 247187 1853
rect 223040 1788 244274 1816
rect 219526 1748 219532 1760
rect 217980 1720 219532 1748
rect 214892 1708 214898 1720
rect 219526 1708 219532 1720
rect 219584 1708 219590 1760
rect 221366 1708 221372 1760
rect 221424 1748 221430 1760
rect 221918 1748 221924 1760
rect 221424 1720 221924 1748
rect 221424 1708 221430 1720
rect 221918 1708 221924 1720
rect 221976 1708 221982 1760
rect 223390 1708 223396 1760
rect 223448 1708 223454 1760
rect 225141 1751 225199 1757
rect 225141 1717 225153 1751
rect 225187 1748 225199 1751
rect 225506 1748 225512 1760
rect 225187 1720 225512 1748
rect 225187 1717 225199 1720
rect 225141 1711 225199 1717
rect 225506 1708 225512 1720
rect 225564 1708 225570 1760
rect 227438 1708 227444 1760
rect 227496 1708 227502 1760
rect 228542 1708 228548 1760
rect 228600 1748 228606 1760
rect 229281 1751 229339 1757
rect 229281 1748 229293 1751
rect 228600 1720 229293 1748
rect 228600 1708 228606 1720
rect 229281 1717 229293 1720
rect 229327 1717 229339 1751
rect 229281 1711 229339 1717
rect 230106 1708 230112 1760
rect 230164 1708 230170 1760
rect 233694 1708 233700 1760
rect 233752 1748 233758 1760
rect 234433 1751 234491 1757
rect 234433 1748 234445 1751
rect 233752 1720 234445 1748
rect 233752 1708 233758 1720
rect 234433 1717 234445 1720
rect 234479 1717 234491 1751
rect 234433 1711 234491 1717
rect 235258 1708 235264 1760
rect 235316 1708 235322 1760
rect 237374 1708 237380 1760
rect 237432 1748 237438 1760
rect 237561 1751 237619 1757
rect 237561 1748 237573 1751
rect 237432 1720 237573 1748
rect 237432 1708 237438 1720
rect 237561 1717 237573 1720
rect 237607 1717 237619 1751
rect 244246 1748 244274 1788
rect 245746 1776 245752 1828
rect 245804 1816 245810 1828
rect 247144 1816 247172 1847
rect 245804 1788 247172 1816
rect 247236 1816 247264 1924
rect 247402 1912 247408 1964
rect 247460 1912 247466 1964
rect 247512 1952 247540 2060
rect 248874 2048 248880 2100
rect 248932 2088 248938 2100
rect 248932 2060 255544 2088
rect 248932 2048 248938 2060
rect 252370 1980 252376 2032
rect 252428 2020 252434 2032
rect 255222 2020 255228 2032
rect 252428 1992 255228 2020
rect 252428 1980 252434 1992
rect 255222 1980 255228 1992
rect 255280 1980 255286 2032
rect 255516 1961 255544 2060
rect 260282 2048 260288 2100
rect 260340 2088 260346 2100
rect 260561 2091 260619 2097
rect 260561 2088 260573 2091
rect 260340 2060 260573 2088
rect 260340 2048 260346 2060
rect 260561 2057 260573 2060
rect 260607 2057 260619 2091
rect 260561 2051 260619 2057
rect 261110 2048 261116 2100
rect 261168 2088 261174 2100
rect 261665 2091 261723 2097
rect 261665 2088 261677 2091
rect 261168 2060 261677 2088
rect 261168 2048 261174 2060
rect 261665 2057 261677 2060
rect 261711 2057 261723 2091
rect 261665 2051 261723 2057
rect 263134 2048 263140 2100
rect 263192 2088 263198 2100
rect 263321 2091 263379 2097
rect 263321 2088 263333 2091
rect 263192 2060 263333 2088
rect 263192 2048 263198 2060
rect 263321 2057 263333 2060
rect 263367 2057 263379 2091
rect 268838 2088 268844 2100
rect 263321 2051 263379 2057
rect 263566 2060 268844 2088
rect 255682 1980 255688 2032
rect 255740 1980 255746 2032
rect 257341 2023 257399 2029
rect 257341 1989 257353 2023
rect 257387 2020 257399 2023
rect 263566 2020 263594 2060
rect 268838 2048 268844 2060
rect 268896 2048 268902 2100
rect 257387 1992 263594 2020
rect 257387 1989 257399 1992
rect 257341 1983 257399 1989
rect 263962 1980 263968 2032
rect 264020 2020 264026 2032
rect 268562 2020 268568 2032
rect 264020 1992 268568 2020
rect 264020 1980 264026 1992
rect 268562 1980 268568 1992
rect 268620 1980 268626 2032
rect 269942 2020 269948 2032
rect 269408 1992 269948 2020
rect 248693 1955 248751 1961
rect 248693 1952 248705 1955
rect 247512 1924 248705 1952
rect 248693 1921 248705 1924
rect 248739 1921 248751 1955
rect 254121 1955 254179 1961
rect 254121 1952 254133 1955
rect 248693 1915 248751 1921
rect 250088 1924 254133 1952
rect 247494 1844 247500 1896
rect 247552 1884 247558 1896
rect 248877 1887 248935 1893
rect 248877 1884 248889 1887
rect 247552 1856 248889 1884
rect 247552 1844 247558 1856
rect 248877 1853 248889 1856
rect 248923 1853 248935 1887
rect 250088 1884 250116 1924
rect 254121 1921 254133 1924
rect 254167 1921 254179 1955
rect 254121 1915 254179 1921
rect 255501 1955 255559 1961
rect 255501 1921 255513 1955
rect 255547 1921 255559 1955
rect 258077 1955 258135 1961
rect 258077 1952 258089 1955
rect 255501 1915 255559 1921
rect 257632 1924 258089 1952
rect 248877 1847 248935 1853
rect 248984 1856 250116 1884
rect 248984 1816 249012 1856
rect 250530 1844 250536 1896
rect 250588 1844 250594 1896
rect 250993 1887 251051 1893
rect 250993 1853 251005 1887
rect 251039 1853 251051 1887
rect 250993 1847 251051 1853
rect 247236 1788 249012 1816
rect 245804 1776 245810 1788
rect 249794 1776 249800 1828
rect 249852 1816 249858 1828
rect 251008 1816 251036 1847
rect 251266 1844 251272 1896
rect 251324 1844 251330 1896
rect 251358 1844 251364 1896
rect 251416 1884 251422 1896
rect 252281 1887 252339 1893
rect 252281 1884 252293 1887
rect 251416 1856 252293 1884
rect 251416 1844 251422 1856
rect 252281 1853 252293 1856
rect 252327 1853 252339 1887
rect 252281 1847 252339 1853
rect 252557 1887 252615 1893
rect 252557 1853 252569 1887
rect 252603 1853 252615 1887
rect 252557 1847 252615 1853
rect 253845 1887 253903 1893
rect 253845 1853 253857 1887
rect 253891 1853 253903 1887
rect 253845 1847 253903 1853
rect 252572 1816 252600 1847
rect 249852 1788 251036 1816
rect 251100 1788 252600 1816
rect 249852 1776 249858 1788
rect 251100 1748 251128 1788
rect 244246 1720 251128 1748
rect 237561 1711 237619 1717
rect 252554 1708 252560 1760
rect 252612 1748 252618 1760
rect 253860 1748 253888 1847
rect 252612 1720 253888 1748
rect 252612 1708 252618 1720
rect 255682 1708 255688 1760
rect 255740 1748 255746 1760
rect 257632 1757 257660 1924
rect 258077 1921 258089 1924
rect 258123 1952 258135 1955
rect 258442 1952 258448 1964
rect 258123 1924 258448 1952
rect 258123 1921 258135 1924
rect 258077 1915 258135 1921
rect 258442 1912 258448 1924
rect 258500 1912 258506 1964
rect 258534 1912 258540 1964
rect 258592 1952 258598 1964
rect 259273 1955 259331 1961
rect 259273 1952 259285 1955
rect 258592 1924 259285 1952
rect 258592 1912 258598 1924
rect 259273 1921 259285 1924
rect 259319 1921 259331 1955
rect 259273 1915 259331 1921
rect 260466 1912 260472 1964
rect 260524 1952 260530 1964
rect 261386 1952 261392 1964
rect 260524 1924 261392 1952
rect 260524 1912 260530 1924
rect 261386 1912 261392 1924
rect 261444 1912 261450 1964
rect 261478 1912 261484 1964
rect 261536 1912 261542 1964
rect 261754 1912 261760 1964
rect 261812 1952 261818 1964
rect 262125 1955 262183 1961
rect 262125 1952 262137 1955
rect 261812 1924 262137 1952
rect 261812 1912 261818 1924
rect 262125 1921 262137 1924
rect 262171 1921 262183 1955
rect 262125 1915 262183 1921
rect 262309 1955 262367 1961
rect 262309 1921 262321 1955
rect 262355 1921 262367 1955
rect 262309 1915 262367 1921
rect 258166 1844 258172 1896
rect 258224 1884 258230 1896
rect 258997 1887 259055 1893
rect 258997 1884 259009 1887
rect 258224 1856 259009 1884
rect 258224 1844 258230 1856
rect 258997 1853 259009 1856
rect 259043 1853 259055 1887
rect 258997 1847 259055 1853
rect 260190 1844 260196 1896
rect 260248 1884 260254 1896
rect 261297 1887 261355 1893
rect 261297 1884 261309 1887
rect 260248 1856 261309 1884
rect 260248 1844 260254 1856
rect 261297 1853 261309 1856
rect 261343 1853 261355 1887
rect 261496 1884 261524 1912
rect 262324 1884 262352 1915
rect 262858 1912 262864 1964
rect 262916 1952 262922 1964
rect 262953 1955 263011 1961
rect 262953 1952 262965 1955
rect 262916 1924 262965 1952
rect 262916 1912 262922 1924
rect 262953 1921 262965 1924
rect 262999 1921 263011 1955
rect 262953 1915 263011 1921
rect 263137 1955 263195 1961
rect 263137 1921 263149 1955
rect 263183 1921 263195 1955
rect 263137 1915 263195 1921
rect 263152 1884 263180 1915
rect 264054 1912 264060 1964
rect 264112 1952 264118 1964
rect 264149 1955 264207 1961
rect 264149 1952 264161 1955
rect 264112 1924 264161 1952
rect 264112 1912 264118 1924
rect 264149 1921 264161 1924
rect 264195 1921 264207 1955
rect 264149 1915 264207 1921
rect 264330 1912 264336 1964
rect 264388 1912 264394 1964
rect 264422 1912 264428 1964
rect 264480 1952 264486 1964
rect 264977 1955 265035 1961
rect 264977 1952 264989 1955
rect 264480 1924 264989 1952
rect 264480 1912 264486 1924
rect 264977 1921 264989 1924
rect 265023 1921 265035 1955
rect 264977 1915 265035 1921
rect 265158 1912 265164 1964
rect 265216 1912 265222 1964
rect 265802 1912 265808 1964
rect 265860 1912 265866 1964
rect 265989 1955 266047 1961
rect 265989 1921 266001 1955
rect 266035 1921 266047 1955
rect 265989 1915 266047 1921
rect 264348 1884 264376 1912
rect 261496 1856 264376 1884
rect 265176 1884 265204 1912
rect 266004 1884 266032 1915
rect 266538 1912 266544 1964
rect 266596 1952 266602 1964
rect 266633 1955 266691 1961
rect 266633 1952 266645 1955
rect 266596 1924 266645 1952
rect 266596 1912 266602 1924
rect 266633 1921 266645 1924
rect 266679 1921 266691 1955
rect 266633 1915 266691 1921
rect 266817 1955 266875 1961
rect 266817 1921 266829 1955
rect 266863 1921 266875 1955
rect 266817 1915 266875 1921
rect 266832 1884 266860 1915
rect 266998 1912 267004 1964
rect 267056 1912 267062 1964
rect 267366 1912 267372 1964
rect 267424 1952 267430 1964
rect 267461 1955 267519 1961
rect 267461 1952 267473 1955
rect 267424 1924 267473 1952
rect 267424 1912 267430 1924
rect 267461 1921 267473 1924
rect 267507 1921 267519 1955
rect 267461 1915 267519 1921
rect 267645 1955 267703 1961
rect 267645 1921 267657 1955
rect 267691 1921 267703 1955
rect 267645 1915 267703 1921
rect 267660 1884 267688 1915
rect 267734 1912 267740 1964
rect 267792 1952 267798 1964
rect 268289 1955 268347 1961
rect 268289 1952 268301 1955
rect 267792 1924 268301 1952
rect 267792 1912 267798 1924
rect 268289 1921 268301 1924
rect 268335 1921 268347 1955
rect 268289 1915 268347 1921
rect 268473 1955 268531 1961
rect 268473 1921 268485 1955
rect 268519 1952 268531 1955
rect 269114 1952 269120 1964
rect 268519 1924 269120 1952
rect 268519 1921 268531 1924
rect 268473 1915 268531 1921
rect 268488 1884 268516 1915
rect 269114 1912 269120 1924
rect 269172 1912 269178 1964
rect 269408 1961 269436 1992
rect 269942 1980 269948 1992
rect 270000 1980 270006 2032
rect 269393 1955 269451 1961
rect 269393 1921 269405 1955
rect 269439 1921 269451 1955
rect 269393 1915 269451 1921
rect 269485 1955 269543 1961
rect 269485 1921 269497 1955
rect 269531 1952 269543 1955
rect 269669 1955 269727 1961
rect 269531 1924 269620 1952
rect 269531 1921 269543 1924
rect 269485 1915 269543 1921
rect 265176 1856 268516 1884
rect 269132 1884 269160 1912
rect 269592 1884 269620 1924
rect 269669 1921 269681 1955
rect 269715 1952 269727 1955
rect 270129 1955 270187 1961
rect 270129 1952 270141 1955
rect 269715 1924 270141 1952
rect 269715 1921 269727 1924
rect 269669 1915 269727 1921
rect 270129 1921 270141 1924
rect 270175 1921 270187 1955
rect 270129 1915 270187 1921
rect 269132 1856 269620 1884
rect 261297 1847 261355 1853
rect 271138 1776 271144 1828
rect 271196 1816 271202 1828
rect 272150 1816 272156 1828
rect 271196 1788 272156 1816
rect 271196 1776 271202 1788
rect 272150 1776 272156 1788
rect 272208 1776 272214 1828
rect 257617 1751 257675 1757
rect 257617 1748 257629 1751
rect 255740 1720 257629 1748
rect 255740 1708 255746 1720
rect 257617 1717 257629 1720
rect 257663 1717 257675 1751
rect 257617 1711 257675 1717
rect 257706 1708 257712 1760
rect 257764 1748 257770 1760
rect 257982 1748 257988 1760
rect 257764 1720 257988 1748
rect 257764 1708 257770 1720
rect 257982 1708 257988 1720
rect 258040 1748 258046 1760
rect 258169 1751 258227 1757
rect 258169 1748 258181 1751
rect 258040 1720 258181 1748
rect 258040 1708 258046 1720
rect 258169 1717 258181 1720
rect 258215 1717 258227 1751
rect 258169 1711 258227 1717
rect 262493 1751 262551 1757
rect 262493 1717 262505 1751
rect 262539 1748 262551 1751
rect 263134 1748 263140 1760
rect 262539 1720 263140 1748
rect 262539 1717 262551 1720
rect 262493 1711 262551 1717
rect 263134 1708 263140 1720
rect 263192 1708 263198 1760
rect 264146 1708 264152 1760
rect 264204 1748 264210 1760
rect 264517 1751 264575 1757
rect 264517 1748 264529 1751
rect 264204 1720 264529 1748
rect 264204 1708 264210 1720
rect 264517 1717 264529 1720
rect 264563 1717 264575 1751
rect 264517 1711 264575 1717
rect 265345 1751 265403 1757
rect 265345 1717 265357 1751
rect 265391 1748 265403 1751
rect 265618 1748 265624 1760
rect 265391 1720 265624 1748
rect 265391 1717 265403 1720
rect 265345 1711 265403 1717
rect 265618 1708 265624 1720
rect 265676 1708 265682 1760
rect 266173 1751 266231 1757
rect 266173 1717 266185 1751
rect 266219 1748 266231 1751
rect 266722 1748 266728 1760
rect 266219 1720 266728 1748
rect 266219 1717 266231 1720
rect 266173 1711 266231 1717
rect 266722 1708 266728 1720
rect 266780 1708 266786 1760
rect 267826 1708 267832 1760
rect 267884 1708 267890 1760
rect 268194 1708 268200 1760
rect 268252 1748 268258 1760
rect 268657 1751 268715 1757
rect 268657 1748 268669 1751
rect 268252 1720 268669 1748
rect 268252 1708 268258 1720
rect 268657 1717 268669 1720
rect 268703 1717 268715 1751
rect 268657 1711 268715 1717
rect 269758 1708 269764 1760
rect 269816 1748 269822 1760
rect 270313 1751 270371 1757
rect 270313 1748 270325 1751
rect 269816 1720 270325 1748
rect 269816 1708 269822 1720
rect 270313 1717 270325 1720
rect 270359 1717 270371 1751
rect 270313 1711 270371 1717
rect 1104 1658 271492 1680
rect 1104 1606 34748 1658
rect 34800 1606 34812 1658
rect 34864 1606 34876 1658
rect 34928 1606 34940 1658
rect 34992 1606 35004 1658
rect 35056 1606 102345 1658
rect 102397 1606 102409 1658
rect 102461 1606 102473 1658
rect 102525 1606 102537 1658
rect 102589 1606 102601 1658
rect 102653 1606 169942 1658
rect 169994 1606 170006 1658
rect 170058 1606 170070 1658
rect 170122 1606 170134 1658
rect 170186 1606 170198 1658
rect 170250 1606 237539 1658
rect 237591 1606 237603 1658
rect 237655 1606 237667 1658
rect 237719 1606 237731 1658
rect 237783 1606 237795 1658
rect 237847 1606 271492 1658
rect 1104 1584 271492 1606
rect 20714 1504 20720 1556
rect 20772 1544 20778 1556
rect 25038 1544 25044 1556
rect 20772 1516 25044 1544
rect 20772 1504 20778 1516
rect 25038 1504 25044 1516
rect 25096 1504 25102 1556
rect 27430 1504 27436 1556
rect 27488 1544 27494 1556
rect 27525 1547 27583 1553
rect 27525 1544 27537 1547
rect 27488 1516 27537 1544
rect 27488 1504 27494 1516
rect 27525 1513 27537 1516
rect 27571 1513 27583 1547
rect 27525 1507 27583 1513
rect 27614 1504 27620 1556
rect 27672 1544 27678 1556
rect 54294 1544 54300 1556
rect 27672 1516 54300 1544
rect 27672 1504 27678 1516
rect 54294 1504 54300 1516
rect 54352 1504 54358 1556
rect 58066 1504 58072 1556
rect 58124 1544 58130 1556
rect 58713 1547 58771 1553
rect 58713 1544 58725 1547
rect 58124 1516 58725 1544
rect 58124 1504 58130 1516
rect 58713 1513 58725 1516
rect 58759 1513 58771 1547
rect 58713 1507 58771 1513
rect 62206 1504 62212 1556
rect 62264 1544 62270 1556
rect 62393 1547 62451 1553
rect 62393 1544 62405 1547
rect 62264 1516 62405 1544
rect 62264 1504 62270 1516
rect 62393 1513 62405 1516
rect 62439 1513 62451 1547
rect 62393 1507 62451 1513
rect 73430 1504 73436 1556
rect 73488 1544 73494 1556
rect 73488 1516 92796 1544
rect 73488 1504 73494 1516
rect 24762 1436 24768 1488
rect 24820 1476 24826 1488
rect 24820 1448 28994 1476
rect 24820 1436 24826 1448
rect 22646 1368 22652 1420
rect 22704 1408 22710 1420
rect 22833 1411 22891 1417
rect 22833 1408 22845 1411
rect 22704 1380 22845 1408
rect 22704 1368 22710 1380
rect 22833 1377 22845 1380
rect 22879 1377 22891 1411
rect 22833 1371 22891 1377
rect 23661 1411 23719 1417
rect 23661 1377 23673 1411
rect 23707 1408 23719 1411
rect 23750 1408 23756 1420
rect 23707 1380 23756 1408
rect 23707 1377 23719 1380
rect 23661 1371 23719 1377
rect 23750 1368 23756 1380
rect 23808 1368 23814 1420
rect 25041 1411 25099 1417
rect 25041 1377 25053 1411
rect 25087 1408 25099 1411
rect 25130 1408 25136 1420
rect 25087 1380 25136 1408
rect 25087 1377 25099 1380
rect 25041 1371 25099 1377
rect 25130 1368 25136 1380
rect 25188 1368 25194 1420
rect 25682 1368 25688 1420
rect 25740 1408 25746 1420
rect 25869 1411 25927 1417
rect 25869 1408 25881 1411
rect 25740 1380 25881 1408
rect 25740 1368 25746 1380
rect 25869 1377 25881 1380
rect 25915 1377 25927 1411
rect 25869 1371 25927 1377
rect 27062 1368 27068 1420
rect 27120 1408 27126 1420
rect 27157 1411 27215 1417
rect 27157 1408 27169 1411
rect 27120 1380 27169 1408
rect 27120 1368 27126 1380
rect 27157 1377 27169 1380
rect 27203 1377 27215 1411
rect 28966 1408 28994 1448
rect 31294 1436 31300 1488
rect 31352 1476 31358 1488
rect 65058 1476 65064 1488
rect 31352 1448 65064 1476
rect 31352 1436 31358 1448
rect 65058 1436 65064 1448
rect 65116 1436 65122 1488
rect 82630 1436 82636 1488
rect 82688 1476 82694 1488
rect 92382 1476 92388 1488
rect 82688 1448 92388 1476
rect 82688 1436 82694 1448
rect 92382 1436 92388 1448
rect 92440 1436 92446 1488
rect 92768 1476 92796 1516
rect 92842 1504 92848 1556
rect 92900 1544 92906 1556
rect 95329 1547 95387 1553
rect 95329 1544 95341 1547
rect 92900 1516 95341 1544
rect 92900 1504 92906 1516
rect 95329 1513 95341 1516
rect 95375 1513 95387 1547
rect 95329 1507 95387 1513
rect 95510 1504 95516 1556
rect 95568 1544 95574 1556
rect 96982 1544 96988 1556
rect 95568 1516 96988 1544
rect 95568 1504 95574 1516
rect 96982 1504 96988 1516
rect 97040 1504 97046 1556
rect 98549 1547 98607 1553
rect 97460 1516 98316 1544
rect 97460 1488 97488 1516
rect 96065 1479 96123 1485
rect 96065 1476 96077 1479
rect 92768 1448 96077 1476
rect 96065 1445 96077 1448
rect 96111 1445 96123 1479
rect 96065 1439 96123 1445
rect 97353 1479 97411 1485
rect 97353 1445 97365 1479
rect 97399 1476 97411 1479
rect 97442 1476 97448 1488
rect 97399 1448 97448 1476
rect 97399 1445 97411 1448
rect 97353 1439 97411 1445
rect 53834 1408 53840 1420
rect 28966 1380 53840 1408
rect 27157 1371 27215 1377
rect 53834 1368 53840 1380
rect 53892 1368 53898 1420
rect 54294 1368 54300 1420
rect 54352 1368 54358 1420
rect 58158 1368 58164 1420
rect 58216 1408 58222 1420
rect 58345 1411 58403 1417
rect 58345 1408 58357 1411
rect 58216 1380 58357 1408
rect 58216 1368 58222 1380
rect 58345 1377 58357 1380
rect 58391 1408 58403 1411
rect 59538 1408 59544 1420
rect 58391 1380 59544 1408
rect 58391 1377 58403 1380
rect 58345 1371 58403 1377
rect 59538 1368 59544 1380
rect 59596 1368 59602 1420
rect 62022 1368 62028 1420
rect 62080 1368 62086 1420
rect 65981 1411 66039 1417
rect 65981 1377 65993 1411
rect 66027 1408 66039 1411
rect 66070 1408 66076 1420
rect 66027 1380 66076 1408
rect 66027 1377 66039 1380
rect 65981 1371 66039 1377
rect 66070 1368 66076 1380
rect 66128 1368 66134 1420
rect 69106 1368 69112 1420
rect 69164 1368 69170 1420
rect 72896 1380 73108 1408
rect 2593 1343 2651 1349
rect 2593 1309 2605 1343
rect 2639 1309 2651 1343
rect 2593 1303 2651 1309
rect 1946 1232 1952 1284
rect 2004 1232 2010 1284
rect 2608 1272 2636 1303
rect 2866 1300 2872 1352
rect 2924 1300 2930 1352
rect 5169 1343 5227 1349
rect 5169 1309 5181 1343
rect 5215 1340 5227 1343
rect 5350 1340 5356 1352
rect 5215 1312 5356 1340
rect 5215 1309 5227 1312
rect 5169 1303 5227 1309
rect 5350 1300 5356 1312
rect 5408 1300 5414 1352
rect 5442 1300 5448 1352
rect 5500 1300 5506 1352
rect 7742 1300 7748 1352
rect 7800 1300 7806 1352
rect 8018 1300 8024 1352
rect 8076 1300 8082 1352
rect 10318 1300 10324 1352
rect 10376 1300 10382 1352
rect 10594 1300 10600 1352
rect 10652 1300 10658 1352
rect 11698 1300 11704 1352
rect 11756 1300 11762 1352
rect 11977 1343 12035 1349
rect 11977 1309 11989 1343
rect 12023 1340 12035 1343
rect 14274 1340 14280 1352
rect 12023 1312 14280 1340
rect 12023 1309 12035 1312
rect 11977 1303 12035 1309
rect 14274 1300 14280 1312
rect 14332 1300 14338 1352
rect 15473 1343 15531 1349
rect 15473 1309 15485 1343
rect 15519 1340 15531 1343
rect 15654 1340 15660 1352
rect 15519 1312 15660 1340
rect 15519 1309 15531 1312
rect 15473 1303 15531 1309
rect 15654 1300 15660 1312
rect 15712 1300 15718 1352
rect 15746 1300 15752 1352
rect 15804 1300 15810 1352
rect 17034 1300 17040 1352
rect 17092 1300 17098 1352
rect 17310 1300 17316 1352
rect 17368 1300 17374 1352
rect 22094 1300 22100 1352
rect 22152 1300 22158 1352
rect 23017 1343 23075 1349
rect 23017 1309 23029 1343
rect 23063 1309 23075 1343
rect 23017 1303 23075 1309
rect 2958 1272 2964 1284
rect 2608 1244 2964 1272
rect 2958 1232 2964 1244
rect 3016 1232 3022 1284
rect 13446 1232 13452 1284
rect 13504 1232 13510 1284
rect 18598 1232 18604 1284
rect 18656 1232 18662 1284
rect 23032 1272 23060 1303
rect 23198 1300 23204 1352
rect 23256 1300 23262 1352
rect 23845 1343 23903 1349
rect 23845 1309 23857 1343
rect 23891 1309 23903 1343
rect 23845 1303 23903 1309
rect 24029 1343 24087 1349
rect 24029 1309 24041 1343
rect 24075 1340 24087 1343
rect 24946 1340 24952 1352
rect 24075 1312 24952 1340
rect 24075 1309 24087 1312
rect 24029 1303 24087 1309
rect 23860 1272 23888 1303
rect 24946 1300 24952 1312
rect 25004 1300 25010 1352
rect 25225 1343 25283 1349
rect 25225 1309 25237 1343
rect 25271 1309 25283 1343
rect 25225 1303 25283 1309
rect 25240 1272 25268 1303
rect 25406 1300 25412 1352
rect 25464 1300 25470 1352
rect 26050 1300 26056 1352
rect 26108 1300 26114 1352
rect 26234 1300 26240 1352
rect 26292 1300 26298 1352
rect 27338 1300 27344 1352
rect 27396 1300 27402 1352
rect 27982 1300 27988 1352
rect 28040 1300 28046 1352
rect 28810 1300 28816 1352
rect 28868 1300 28874 1352
rect 30285 1343 30343 1349
rect 30285 1309 30297 1343
rect 30331 1340 30343 1343
rect 30374 1340 30380 1352
rect 30331 1312 30380 1340
rect 30331 1309 30343 1312
rect 30285 1303 30343 1309
rect 30374 1300 30380 1312
rect 30432 1300 30438 1352
rect 31018 1300 31024 1352
rect 31076 1300 31082 1352
rect 32306 1300 32312 1352
rect 32364 1300 32370 1352
rect 35618 1300 35624 1352
rect 35676 1300 35682 1352
rect 36262 1300 36268 1352
rect 36320 1300 36326 1352
rect 36906 1300 36912 1352
rect 36964 1300 36970 1352
rect 38197 1343 38255 1349
rect 38197 1309 38209 1343
rect 38243 1340 38255 1343
rect 38562 1340 38568 1352
rect 38243 1312 38568 1340
rect 38243 1309 38255 1312
rect 38197 1303 38255 1309
rect 38562 1300 38568 1312
rect 38620 1300 38626 1352
rect 38838 1300 38844 1352
rect 38896 1300 38902 1352
rect 39485 1343 39543 1349
rect 39485 1309 39497 1343
rect 39531 1340 39543 1343
rect 39942 1340 39948 1352
rect 39531 1312 39948 1340
rect 39531 1309 39543 1312
rect 39485 1303 39543 1309
rect 39942 1300 39948 1312
rect 40000 1300 40006 1352
rect 40770 1300 40776 1352
rect 40828 1300 40834 1352
rect 41414 1300 41420 1352
rect 41472 1300 41478 1352
rect 42058 1300 42064 1352
rect 42116 1300 42122 1352
rect 43254 1300 43260 1352
rect 43312 1300 43318 1352
rect 43990 1300 43996 1352
rect 44048 1300 44054 1352
rect 44634 1300 44640 1352
rect 44692 1300 44698 1352
rect 45922 1300 45928 1352
rect 45980 1300 45986 1352
rect 46566 1300 46572 1352
rect 46624 1300 46630 1352
rect 47210 1300 47216 1352
rect 47268 1300 47274 1352
rect 48222 1300 48228 1352
rect 48280 1340 48286 1352
rect 48409 1343 48467 1349
rect 48409 1340 48421 1343
rect 48280 1312 48421 1340
rect 48280 1300 48286 1312
rect 48409 1309 48421 1312
rect 48455 1309 48467 1343
rect 48409 1303 48467 1309
rect 49142 1300 49148 1352
rect 49200 1300 49206 1352
rect 49786 1300 49792 1352
rect 49844 1300 49850 1352
rect 50614 1300 50620 1352
rect 50672 1300 50678 1352
rect 51350 1300 51356 1352
rect 51408 1300 51414 1352
rect 52086 1300 52092 1352
rect 52144 1300 52150 1352
rect 53098 1300 53104 1352
rect 53156 1300 53162 1352
rect 54481 1343 54539 1349
rect 54481 1309 54493 1343
rect 54527 1340 54539 1343
rect 54570 1340 54576 1352
rect 54527 1312 54576 1340
rect 54527 1309 54539 1312
rect 54481 1303 54539 1309
rect 54570 1300 54576 1312
rect 54628 1300 54634 1352
rect 54662 1300 54668 1352
rect 54720 1300 54726 1352
rect 55030 1300 55036 1352
rect 55088 1340 55094 1352
rect 55493 1343 55551 1349
rect 55493 1340 55505 1343
rect 55088 1312 55505 1340
rect 55088 1300 55094 1312
rect 55493 1309 55505 1312
rect 55539 1309 55551 1343
rect 55493 1303 55551 1309
rect 56226 1300 56232 1352
rect 56284 1300 56290 1352
rect 56962 1300 56968 1352
rect 57020 1300 57026 1352
rect 58526 1300 58532 1352
rect 58584 1300 58590 1352
rect 59814 1300 59820 1352
rect 59872 1300 59878 1352
rect 60734 1300 60740 1352
rect 60792 1300 60798 1352
rect 62209 1343 62267 1349
rect 62209 1309 62221 1343
rect 62255 1340 62267 1343
rect 62482 1340 62488 1352
rect 62255 1312 62488 1340
rect 62255 1309 62267 1312
rect 62209 1303 62267 1309
rect 62482 1300 62488 1312
rect 62540 1300 62546 1352
rect 63678 1300 63684 1352
rect 63736 1300 63742 1352
rect 64414 1300 64420 1352
rect 64472 1300 64478 1352
rect 66162 1300 66168 1352
rect 66220 1300 66226 1352
rect 66349 1343 66407 1349
rect 66349 1309 66361 1343
rect 66395 1340 66407 1343
rect 66809 1343 66867 1349
rect 66809 1340 66821 1343
rect 66395 1312 66821 1340
rect 66395 1309 66407 1312
rect 66349 1303 66407 1309
rect 66809 1309 66821 1312
rect 66855 1309 66867 1343
rect 66809 1303 66867 1309
rect 69566 1300 69572 1352
rect 69624 1300 69630 1352
rect 69845 1343 69903 1349
rect 69845 1309 69857 1343
rect 69891 1340 69903 1343
rect 69891 1312 70394 1340
rect 69891 1309 69903 1312
rect 69845 1303 69903 1309
rect 26068 1272 26096 1300
rect 23032 1244 26096 1272
rect 43438 1232 43444 1284
rect 43496 1272 43502 1284
rect 43496 1244 44496 1272
rect 43496 1232 43502 1244
rect 2038 1164 2044 1216
rect 2096 1164 2102 1216
rect 13538 1164 13544 1216
rect 13596 1164 13602 1216
rect 18690 1164 18696 1216
rect 18748 1164 18754 1216
rect 21450 1164 21456 1216
rect 21508 1204 21514 1216
rect 22281 1207 22339 1213
rect 22281 1204 22293 1207
rect 21508 1176 22293 1204
rect 21508 1164 21514 1176
rect 22281 1173 22293 1176
rect 22327 1173 22339 1207
rect 22281 1167 22339 1173
rect 28166 1164 28172 1216
rect 28224 1164 28230 1216
rect 28994 1164 29000 1216
rect 29052 1164 29058 1216
rect 30282 1164 30288 1216
rect 30340 1204 30346 1216
rect 30469 1207 30527 1213
rect 30469 1204 30481 1207
rect 30340 1176 30481 1204
rect 30340 1164 30346 1176
rect 30469 1173 30481 1176
rect 30515 1173 30527 1207
rect 30469 1167 30527 1173
rect 31202 1164 31208 1216
rect 31260 1164 31266 1216
rect 32490 1164 32496 1216
rect 32548 1164 32554 1216
rect 35434 1164 35440 1216
rect 35492 1164 35498 1216
rect 36078 1164 36084 1216
rect 36136 1164 36142 1216
rect 36354 1164 36360 1216
rect 36412 1204 36418 1216
rect 36725 1207 36783 1213
rect 36725 1204 36737 1207
rect 36412 1176 36737 1204
rect 36412 1164 36418 1176
rect 36725 1173 36737 1176
rect 36771 1173 36783 1207
rect 36725 1167 36783 1173
rect 37826 1164 37832 1216
rect 37884 1204 37890 1216
rect 38013 1207 38071 1213
rect 38013 1204 38025 1207
rect 37884 1176 38025 1204
rect 37884 1164 37890 1176
rect 38013 1173 38025 1176
rect 38059 1173 38071 1207
rect 38013 1167 38071 1173
rect 38286 1164 38292 1216
rect 38344 1204 38350 1216
rect 38657 1207 38715 1213
rect 38657 1204 38669 1207
rect 38344 1176 38669 1204
rect 38344 1164 38350 1176
rect 38657 1173 38669 1176
rect 38703 1173 38715 1207
rect 38657 1167 38715 1173
rect 39298 1164 39304 1216
rect 39356 1164 39362 1216
rect 40218 1164 40224 1216
rect 40276 1204 40282 1216
rect 40589 1207 40647 1213
rect 40589 1204 40601 1207
rect 40276 1176 40601 1204
rect 40276 1164 40282 1176
rect 40589 1173 40601 1176
rect 40635 1173 40647 1207
rect 40589 1167 40647 1173
rect 41230 1164 41236 1216
rect 41288 1164 41294 1216
rect 41598 1164 41604 1216
rect 41656 1204 41662 1216
rect 41877 1207 41935 1213
rect 41877 1204 41889 1207
rect 41656 1176 41889 1204
rect 41656 1164 41662 1176
rect 41877 1173 41889 1176
rect 41923 1173 41935 1207
rect 41877 1167 41935 1173
rect 42242 1164 42248 1216
rect 42300 1204 42306 1216
rect 43073 1207 43131 1213
rect 43073 1204 43085 1207
rect 42300 1176 43085 1204
rect 42300 1164 42306 1176
rect 43073 1173 43085 1176
rect 43119 1173 43131 1207
rect 43073 1167 43131 1173
rect 43162 1164 43168 1216
rect 43220 1204 43226 1216
rect 44468 1213 44496 1244
rect 47578 1232 47584 1284
rect 47636 1272 47642 1284
rect 70366 1272 70394 1312
rect 70946 1300 70952 1352
rect 71004 1300 71010 1352
rect 71225 1343 71283 1349
rect 71225 1309 71237 1343
rect 71271 1340 71283 1343
rect 72896 1340 72924 1380
rect 71271 1312 72924 1340
rect 71271 1309 71283 1312
rect 71225 1303 71283 1309
rect 72970 1300 72976 1352
rect 73028 1300 73034 1352
rect 73080 1340 73108 1380
rect 74184 1380 74396 1408
rect 74184 1340 74212 1380
rect 73080 1312 74212 1340
rect 74258 1300 74264 1352
rect 74316 1300 74322 1352
rect 74368 1272 74396 1380
rect 89070 1368 89076 1420
rect 89128 1368 89134 1420
rect 89714 1408 89720 1420
rect 89180 1380 89720 1408
rect 74718 1300 74724 1352
rect 74776 1300 74782 1352
rect 74994 1300 75000 1352
rect 75052 1300 75058 1352
rect 77294 1300 77300 1352
rect 77352 1300 77358 1352
rect 77570 1300 77576 1352
rect 77628 1300 77634 1352
rect 79873 1343 79931 1349
rect 79873 1309 79885 1343
rect 79919 1340 79931 1343
rect 79962 1340 79968 1352
rect 79919 1312 79968 1340
rect 79919 1309 79931 1312
rect 79873 1303 79931 1309
rect 79962 1300 79968 1312
rect 80020 1300 80026 1352
rect 80146 1300 80152 1352
rect 80204 1300 80210 1352
rect 82449 1343 82507 1349
rect 82449 1309 82461 1343
rect 82495 1340 82507 1343
rect 82630 1340 82636 1352
rect 82495 1312 82636 1340
rect 82495 1309 82507 1312
rect 82449 1303 82507 1309
rect 82630 1300 82636 1312
rect 82688 1300 82694 1352
rect 82722 1300 82728 1352
rect 82780 1300 82786 1352
rect 85022 1300 85028 1352
rect 85080 1300 85086 1352
rect 85301 1343 85359 1349
rect 85301 1309 85313 1343
rect 85347 1340 85359 1343
rect 85482 1340 85488 1352
rect 85347 1312 85488 1340
rect 85347 1309 85359 1312
rect 85301 1303 85359 1309
rect 85482 1300 85488 1312
rect 85540 1300 85546 1352
rect 86770 1300 86776 1352
rect 86828 1300 86834 1352
rect 87049 1343 87107 1349
rect 87049 1309 87061 1343
rect 87095 1309 87107 1343
rect 87049 1303 87107 1309
rect 88153 1343 88211 1349
rect 88153 1309 88165 1343
rect 88199 1340 88211 1343
rect 88794 1340 88800 1352
rect 88199 1312 88800 1340
rect 88199 1309 88211 1312
rect 88153 1303 88211 1309
rect 84194 1272 84200 1284
rect 47636 1244 49004 1272
rect 70366 1244 74212 1272
rect 74368 1244 84200 1272
rect 47636 1232 47642 1244
rect 43809 1207 43867 1213
rect 43809 1204 43821 1207
rect 43220 1176 43821 1204
rect 43220 1164 43226 1176
rect 43809 1173 43821 1176
rect 43855 1173 43867 1207
rect 43809 1167 43867 1173
rect 44453 1207 44511 1213
rect 44453 1173 44465 1207
rect 44499 1173 44511 1207
rect 44453 1167 44511 1173
rect 45370 1164 45376 1216
rect 45428 1204 45434 1216
rect 45741 1207 45799 1213
rect 45741 1204 45753 1207
rect 45428 1176 45753 1204
rect 45428 1164 45434 1176
rect 45741 1173 45753 1176
rect 45787 1173 45799 1207
rect 45741 1167 45799 1173
rect 45830 1164 45836 1216
rect 45888 1204 45894 1216
rect 46385 1207 46443 1213
rect 46385 1204 46397 1207
rect 45888 1176 46397 1204
rect 45888 1164 45894 1176
rect 46385 1173 46397 1176
rect 46431 1173 46443 1207
rect 46385 1167 46443 1173
rect 47026 1164 47032 1216
rect 47084 1164 47090 1216
rect 47946 1164 47952 1216
rect 48004 1204 48010 1216
rect 48976 1213 49004 1244
rect 48225 1207 48283 1213
rect 48225 1204 48237 1207
rect 48004 1176 48237 1204
rect 48004 1164 48010 1176
rect 48225 1173 48237 1176
rect 48271 1173 48283 1207
rect 48225 1167 48283 1173
rect 48961 1207 49019 1213
rect 48961 1173 48973 1207
rect 49007 1173 49019 1207
rect 48961 1167 49019 1173
rect 49510 1164 49516 1216
rect 49568 1204 49574 1216
rect 49605 1207 49663 1213
rect 49605 1204 49617 1207
rect 49568 1176 49617 1204
rect 49568 1164 49574 1176
rect 49605 1173 49617 1176
rect 49651 1173 49663 1207
rect 49605 1167 49663 1173
rect 50430 1164 50436 1216
rect 50488 1164 50494 1216
rect 51074 1164 51080 1216
rect 51132 1204 51138 1216
rect 51169 1207 51227 1213
rect 51169 1204 51181 1207
rect 51132 1176 51181 1204
rect 51132 1164 51138 1176
rect 51169 1173 51181 1176
rect 51215 1173 51227 1207
rect 51169 1167 51227 1173
rect 51902 1164 51908 1216
rect 51960 1164 51966 1216
rect 51994 1164 52000 1216
rect 52052 1204 52058 1216
rect 52917 1207 52975 1213
rect 52917 1204 52929 1207
rect 52052 1176 52929 1204
rect 52052 1164 52058 1176
rect 52917 1173 52929 1176
rect 52963 1173 52975 1207
rect 52917 1167 52975 1173
rect 55674 1164 55680 1216
rect 55732 1164 55738 1216
rect 56410 1164 56416 1216
rect 56468 1164 56474 1216
rect 57146 1164 57152 1216
rect 57204 1164 57210 1216
rect 59998 1164 60004 1216
rect 60056 1164 60062 1216
rect 60918 1164 60924 1216
rect 60976 1164 60982 1216
rect 63862 1164 63868 1216
rect 63920 1164 63926 1216
rect 64598 1164 64604 1216
rect 64656 1164 64662 1216
rect 65886 1164 65892 1216
rect 65944 1204 65950 1216
rect 66993 1207 67051 1213
rect 66993 1204 67005 1207
rect 65944 1176 67005 1204
rect 65944 1164 65950 1176
rect 66993 1173 67005 1176
rect 67039 1173 67051 1207
rect 66993 1167 67051 1173
rect 72786 1164 72792 1216
rect 72844 1164 72850 1216
rect 74074 1164 74080 1216
rect 74132 1164 74138 1216
rect 74184 1204 74212 1244
rect 84194 1232 84200 1244
rect 84252 1232 84258 1284
rect 87064 1272 87092 1303
rect 88794 1300 88800 1312
rect 88852 1300 88858 1352
rect 89180 1272 89208 1380
rect 89714 1368 89720 1380
rect 89772 1368 89778 1420
rect 90542 1368 90548 1420
rect 90600 1368 90606 1420
rect 94133 1411 94191 1417
rect 94133 1377 94145 1411
rect 94179 1408 94191 1411
rect 94498 1408 94504 1420
rect 94179 1380 94504 1408
rect 94179 1377 94191 1380
rect 94133 1371 94191 1377
rect 94498 1368 94504 1380
rect 94556 1368 94562 1420
rect 94958 1368 94964 1420
rect 95016 1368 95022 1420
rect 95421 1411 95479 1417
rect 95421 1377 95433 1411
rect 95467 1408 95479 1411
rect 95786 1408 95792 1420
rect 95467 1380 95792 1408
rect 95467 1377 95479 1380
rect 95421 1371 95479 1377
rect 95786 1368 95792 1380
rect 95844 1368 95850 1420
rect 96080 1408 96108 1439
rect 97442 1436 97448 1448
rect 97500 1436 97506 1488
rect 98288 1476 98316 1516
rect 98549 1513 98561 1547
rect 98595 1544 98607 1547
rect 99282 1544 99288 1556
rect 98595 1516 99288 1544
rect 98595 1513 98607 1516
rect 98549 1507 98607 1513
rect 99282 1504 99288 1516
rect 99340 1504 99346 1556
rect 105170 1544 105176 1556
rect 100312 1516 105176 1544
rect 100312 1485 100340 1516
rect 105170 1504 105176 1516
rect 105228 1544 105234 1556
rect 107746 1544 107752 1556
rect 105228 1516 107752 1544
rect 105228 1504 105234 1516
rect 105280 1485 105308 1516
rect 107746 1504 107752 1516
rect 107804 1504 107810 1556
rect 111334 1544 111340 1556
rect 107856 1516 111340 1544
rect 107856 1488 107884 1516
rect 100297 1479 100355 1485
rect 100297 1476 100309 1479
rect 98288 1448 100309 1476
rect 100297 1445 100309 1448
rect 100343 1445 100355 1479
rect 100297 1439 100355 1445
rect 105265 1479 105323 1485
rect 105265 1445 105277 1479
rect 105311 1445 105323 1479
rect 105265 1439 105323 1445
rect 107838 1436 107844 1488
rect 107896 1436 107902 1488
rect 109034 1436 109040 1488
rect 109092 1436 109098 1488
rect 110432 1485 110460 1516
rect 111334 1504 111340 1516
rect 111392 1544 111398 1556
rect 111392 1516 112852 1544
rect 111392 1504 111398 1516
rect 112824 1485 112852 1516
rect 117406 1504 117412 1556
rect 117464 1504 117470 1556
rect 118510 1504 118516 1556
rect 118568 1504 118574 1556
rect 120074 1504 120080 1556
rect 120132 1544 120138 1556
rect 120169 1547 120227 1553
rect 120169 1544 120181 1547
rect 120132 1516 120181 1544
rect 120132 1504 120138 1516
rect 120169 1513 120181 1516
rect 120215 1513 120227 1547
rect 120169 1507 120227 1513
rect 126054 1504 126060 1556
rect 126112 1544 126118 1556
rect 126517 1547 126575 1553
rect 126517 1544 126529 1547
rect 126112 1516 126529 1544
rect 126112 1504 126118 1516
rect 126517 1513 126529 1516
rect 126563 1513 126575 1547
rect 126517 1507 126575 1513
rect 128998 1504 129004 1556
rect 129056 1544 129062 1556
rect 129277 1547 129335 1553
rect 129277 1544 129289 1547
rect 129056 1516 129289 1544
rect 129056 1504 129062 1516
rect 129277 1513 129289 1516
rect 129323 1513 129335 1547
rect 129277 1507 129335 1513
rect 132466 1516 138244 1544
rect 110417 1479 110475 1485
rect 110417 1445 110429 1479
rect 110463 1445 110475 1479
rect 110417 1439 110475 1445
rect 112809 1479 112867 1485
rect 112809 1445 112821 1479
rect 112855 1445 112867 1479
rect 112809 1439 112867 1445
rect 115569 1479 115627 1485
rect 115569 1445 115581 1479
rect 115615 1476 115627 1479
rect 115658 1476 115664 1488
rect 115615 1448 115664 1476
rect 115615 1445 115627 1448
rect 115569 1439 115627 1445
rect 115658 1436 115664 1448
rect 115716 1436 115722 1488
rect 117130 1436 117136 1488
rect 117188 1476 117194 1488
rect 120718 1476 120724 1488
rect 117188 1448 120724 1476
rect 117188 1436 117194 1448
rect 120718 1436 120724 1448
rect 120776 1436 120782 1488
rect 123110 1436 123116 1488
rect 123168 1476 123174 1488
rect 132466 1476 132494 1516
rect 123168 1448 132494 1476
rect 123168 1436 123174 1448
rect 133506 1436 133512 1488
rect 133564 1436 133570 1488
rect 138014 1436 138020 1488
rect 138072 1476 138078 1488
rect 138109 1479 138167 1485
rect 138109 1476 138121 1479
rect 138072 1448 138121 1476
rect 138072 1436 138078 1448
rect 138109 1445 138121 1448
rect 138155 1445 138167 1479
rect 138216 1476 138244 1516
rect 138290 1504 138296 1556
rect 138348 1544 138354 1556
rect 141234 1544 141240 1556
rect 138348 1516 141240 1544
rect 138348 1504 138354 1516
rect 141234 1504 141240 1516
rect 141292 1504 141298 1556
rect 142154 1504 142160 1556
rect 142212 1504 142218 1556
rect 143442 1504 143448 1556
rect 143500 1544 143506 1556
rect 144917 1547 144975 1553
rect 143500 1516 144868 1544
rect 143500 1504 143506 1516
rect 140866 1476 140872 1488
rect 138216 1448 140872 1476
rect 138109 1439 138167 1445
rect 140866 1436 140872 1448
rect 140924 1436 140930 1488
rect 140961 1479 141019 1485
rect 140961 1445 140973 1479
rect 141007 1476 141019 1479
rect 141050 1476 141056 1488
rect 141007 1448 141056 1476
rect 141007 1445 141019 1448
rect 140961 1439 141019 1445
rect 141050 1436 141056 1448
rect 141108 1436 141114 1488
rect 144840 1476 144868 1516
rect 144917 1513 144929 1547
rect 144963 1544 144975 1547
rect 145374 1544 145380 1556
rect 144963 1516 145380 1544
rect 144963 1513 144975 1516
rect 144917 1507 144975 1513
rect 145374 1504 145380 1516
rect 145432 1504 145438 1556
rect 146662 1504 146668 1556
rect 146720 1544 146726 1556
rect 146720 1516 149836 1544
rect 146720 1504 146726 1516
rect 146294 1476 146300 1488
rect 143368 1448 143856 1476
rect 144840 1448 146300 1476
rect 97629 1411 97687 1417
rect 96080 1380 96844 1408
rect 89257 1343 89315 1349
rect 89257 1309 89269 1343
rect 89303 1340 89315 1343
rect 90726 1340 90732 1352
rect 89303 1312 90732 1340
rect 89303 1309 89315 1312
rect 89257 1303 89315 1309
rect 90726 1300 90732 1312
rect 90784 1300 90790 1352
rect 90910 1300 90916 1352
rect 90968 1300 90974 1352
rect 91646 1300 91652 1352
rect 91704 1300 91710 1352
rect 92385 1343 92443 1349
rect 92385 1309 92397 1343
rect 92431 1340 92443 1343
rect 92431 1312 93072 1340
rect 92431 1309 92443 1312
rect 92385 1303 92443 1309
rect 87064 1244 89208 1272
rect 80238 1204 80244 1216
rect 74184 1176 80244 1204
rect 80238 1164 80244 1176
rect 80296 1164 80302 1216
rect 87506 1164 87512 1216
rect 87564 1204 87570 1216
rect 88337 1207 88395 1213
rect 88337 1204 88349 1207
rect 87564 1176 88349 1204
rect 87564 1164 87570 1176
rect 88337 1173 88349 1176
rect 88383 1173 88395 1207
rect 88337 1167 88395 1173
rect 88426 1164 88432 1216
rect 88484 1204 88490 1216
rect 89441 1207 89499 1213
rect 89441 1204 89453 1207
rect 88484 1176 89453 1204
rect 88484 1164 88490 1176
rect 89441 1173 89453 1176
rect 89487 1173 89499 1207
rect 89441 1167 89499 1173
rect 91833 1207 91891 1213
rect 91833 1173 91845 1207
rect 91879 1204 91891 1207
rect 92474 1204 92480 1216
rect 91879 1176 92480 1204
rect 91879 1173 91891 1176
rect 91833 1167 91891 1173
rect 92474 1164 92480 1176
rect 92532 1164 92538 1216
rect 92566 1164 92572 1216
rect 92624 1164 92630 1216
rect 93044 1204 93072 1312
rect 93210 1300 93216 1352
rect 93268 1300 93274 1352
rect 93302 1300 93308 1352
rect 93360 1300 93366 1352
rect 93394 1300 93400 1352
rect 93452 1340 93458 1352
rect 93489 1343 93547 1349
rect 93489 1340 93501 1343
rect 93452 1312 93501 1340
rect 93452 1300 93458 1312
rect 93489 1309 93501 1312
rect 93535 1309 93547 1343
rect 93489 1303 93547 1309
rect 93578 1300 93584 1352
rect 93636 1340 93642 1352
rect 94317 1343 94375 1349
rect 94317 1340 94329 1343
rect 93636 1312 94329 1340
rect 93636 1300 93642 1312
rect 94317 1309 94329 1312
rect 94363 1309 94375 1343
rect 94317 1303 94375 1309
rect 94406 1300 94412 1352
rect 94464 1340 94470 1352
rect 95145 1343 95203 1349
rect 94464 1312 94912 1340
rect 94464 1300 94470 1312
rect 94884 1272 94912 1312
rect 95145 1309 95157 1343
rect 95191 1340 95203 1343
rect 95602 1340 95608 1352
rect 95191 1312 95608 1340
rect 95191 1309 95203 1312
rect 95145 1303 95203 1309
rect 95602 1300 95608 1312
rect 95660 1300 95666 1352
rect 96522 1300 96528 1352
rect 96580 1340 96586 1352
rect 96709 1343 96767 1349
rect 96709 1340 96721 1343
rect 96580 1312 96721 1340
rect 96580 1300 96586 1312
rect 96709 1309 96721 1312
rect 96755 1309 96767 1343
rect 96816 1340 96844 1380
rect 97629 1377 97641 1411
rect 97675 1408 97687 1411
rect 98454 1408 98460 1420
rect 97675 1380 98460 1408
rect 97675 1377 97687 1380
rect 97629 1371 97687 1377
rect 98454 1368 98460 1380
rect 98512 1368 98518 1420
rect 98914 1368 98920 1420
rect 98972 1408 98978 1420
rect 99193 1411 99251 1417
rect 99193 1408 99205 1411
rect 98972 1380 99205 1408
rect 98972 1368 98978 1380
rect 99193 1377 99205 1380
rect 99239 1377 99251 1411
rect 99193 1371 99251 1377
rect 99300 1380 99512 1408
rect 97810 1349 97816 1352
rect 96893 1343 96951 1349
rect 96893 1340 96905 1343
rect 96816 1312 96905 1340
rect 96709 1303 96767 1309
rect 96893 1309 96905 1312
rect 96939 1309 96951 1343
rect 96893 1303 96951 1309
rect 97767 1343 97816 1349
rect 97767 1309 97779 1343
rect 97813 1309 97816 1343
rect 97767 1303 97816 1309
rect 97810 1300 97816 1303
rect 97868 1300 97874 1352
rect 97902 1300 97908 1352
rect 97960 1300 97966 1352
rect 98641 1343 98699 1349
rect 98641 1309 98653 1343
rect 98687 1309 98699 1343
rect 98641 1303 98699 1309
rect 95789 1275 95847 1281
rect 95789 1272 95801 1275
rect 94884 1244 95801 1272
rect 95789 1241 95801 1244
rect 95835 1241 95847 1275
rect 98656 1272 98684 1303
rect 98730 1300 98736 1352
rect 98788 1340 98794 1352
rect 99300 1340 99328 1380
rect 98788 1312 99328 1340
rect 98788 1300 98794 1312
rect 99374 1300 99380 1352
rect 99432 1300 99438 1352
rect 99484 1340 99512 1380
rect 100570 1368 100576 1420
rect 100628 1368 100634 1420
rect 100711 1411 100769 1417
rect 100711 1377 100723 1411
rect 100757 1408 100769 1411
rect 105817 1411 105875 1417
rect 100757 1380 101812 1408
rect 100757 1377 100769 1380
rect 100711 1371 100769 1377
rect 99653 1343 99711 1349
rect 99653 1340 99665 1343
rect 99484 1312 99665 1340
rect 99653 1309 99665 1312
rect 99699 1309 99711 1343
rect 99653 1303 99711 1309
rect 99834 1300 99840 1352
rect 99892 1300 99898 1352
rect 100846 1300 100852 1352
rect 100904 1300 100910 1352
rect 101490 1300 101496 1352
rect 101548 1300 101554 1352
rect 101674 1300 101680 1352
rect 101732 1300 101738 1352
rect 101784 1340 101812 1380
rect 105817 1377 105829 1411
rect 105863 1408 105875 1411
rect 105998 1408 106004 1420
rect 105863 1380 106004 1408
rect 105863 1377 105875 1380
rect 105817 1371 105875 1377
rect 105998 1368 106004 1380
rect 106056 1408 106062 1420
rect 108393 1411 108451 1417
rect 108393 1408 108405 1411
rect 106056 1380 108405 1408
rect 106056 1368 106062 1380
rect 108393 1377 108405 1380
rect 108439 1408 108451 1411
rect 109218 1408 109224 1420
rect 108439 1380 109224 1408
rect 108439 1377 108451 1380
rect 108393 1371 108451 1377
rect 109218 1368 109224 1380
rect 109276 1368 109282 1420
rect 110690 1368 110696 1420
rect 110748 1368 110754 1420
rect 111334 1408 111340 1420
rect 110984 1380 111340 1408
rect 103882 1340 103888 1352
rect 101784 1312 103888 1340
rect 103882 1300 103888 1312
rect 103940 1300 103946 1352
rect 104618 1300 104624 1352
rect 104676 1300 104682 1352
rect 104805 1343 104863 1349
rect 104805 1309 104817 1343
rect 104851 1309 104863 1343
rect 104805 1303 104863 1309
rect 99561 1275 99619 1281
rect 99561 1272 99573 1275
rect 98656 1244 99573 1272
rect 95789 1235 95847 1241
rect 99561 1241 99573 1244
rect 99607 1241 99619 1275
rect 104820 1272 104848 1303
rect 105538 1300 105544 1352
rect 105596 1300 105602 1352
rect 105722 1349 105728 1352
rect 105679 1343 105728 1349
rect 105679 1309 105691 1343
rect 105725 1309 105728 1343
rect 105679 1303 105728 1309
rect 105722 1300 105728 1303
rect 105780 1300 105786 1352
rect 106458 1300 106464 1352
rect 106516 1300 106522 1352
rect 107194 1300 107200 1352
rect 107252 1300 107258 1352
rect 107378 1300 107384 1352
rect 107436 1300 107442 1352
rect 108114 1300 108120 1352
rect 108172 1300 108178 1352
rect 108298 1349 108304 1352
rect 108255 1343 108304 1349
rect 108255 1309 108267 1343
rect 108301 1309 108304 1343
rect 108255 1303 108304 1309
rect 108298 1300 108304 1303
rect 108356 1300 108362 1352
rect 109773 1343 109831 1349
rect 109773 1340 109785 1343
rect 109006 1312 109785 1340
rect 109006 1284 109034 1312
rect 109773 1309 109785 1312
rect 109819 1309 109831 1343
rect 109773 1303 109831 1309
rect 109954 1300 109960 1352
rect 110012 1300 110018 1352
rect 110782 1300 110788 1352
rect 110840 1349 110846 1352
rect 110984 1349 111012 1380
rect 111334 1368 111340 1380
rect 111392 1408 111398 1420
rect 111794 1408 111800 1420
rect 111392 1380 111800 1408
rect 111392 1368 111398 1380
rect 111794 1368 111800 1380
rect 111852 1408 111858 1420
rect 113361 1411 113419 1417
rect 113361 1408 113373 1411
rect 111852 1380 113373 1408
rect 111852 1368 111858 1380
rect 113361 1377 113373 1380
rect 113407 1377 113419 1411
rect 113361 1371 113419 1377
rect 115983 1411 116041 1417
rect 115983 1377 115995 1411
rect 116029 1408 116041 1411
rect 116029 1380 116716 1408
rect 116029 1377 116041 1380
rect 115983 1371 116041 1377
rect 110840 1343 110868 1349
rect 110856 1309 110868 1343
rect 110840 1303 110868 1309
rect 110969 1343 111027 1349
rect 110969 1309 110981 1343
rect 111015 1309 111027 1343
rect 110969 1303 111027 1309
rect 110840 1300 110846 1303
rect 111610 1300 111616 1352
rect 111668 1300 111674 1352
rect 112165 1343 112223 1349
rect 112165 1309 112177 1343
rect 112211 1309 112223 1343
rect 112165 1303 112223 1309
rect 99561 1235 99619 1241
rect 101324 1244 101904 1272
rect 94501 1207 94559 1213
rect 94501 1204 94513 1207
rect 93044 1176 94513 1204
rect 94501 1173 94513 1176
rect 94547 1173 94559 1207
rect 94501 1167 94559 1173
rect 94590 1164 94596 1216
rect 94648 1204 94654 1216
rect 97350 1204 97356 1216
rect 94648 1176 97356 1204
rect 94648 1164 94654 1176
rect 97350 1164 97356 1176
rect 97408 1164 97414 1216
rect 98825 1207 98883 1213
rect 98825 1173 98837 1207
rect 98871 1204 98883 1207
rect 99282 1204 99288 1216
rect 98871 1176 99288 1204
rect 98871 1173 98883 1176
rect 98825 1167 98883 1173
rect 99282 1164 99288 1176
rect 99340 1164 99346 1216
rect 100754 1164 100760 1216
rect 100812 1204 100818 1216
rect 101324 1204 101352 1244
rect 101876 1213 101904 1244
rect 103808 1244 104848 1272
rect 103808 1216 103836 1244
rect 108942 1232 108948 1284
rect 109000 1244 109034 1284
rect 112180 1272 112208 1303
rect 112346 1300 112352 1352
rect 112404 1300 112410 1352
rect 113082 1300 113088 1352
rect 113140 1300 113146 1352
rect 113266 1349 113272 1352
rect 113223 1343 113272 1349
rect 113223 1309 113235 1343
rect 113269 1309 113272 1343
rect 113223 1303 113272 1309
rect 113266 1300 113272 1303
rect 113324 1300 113330 1352
rect 114922 1300 114928 1352
rect 114980 1300 114986 1352
rect 115106 1300 115112 1352
rect 115164 1300 115170 1352
rect 115842 1300 115848 1352
rect 115900 1300 115906 1352
rect 116118 1300 116124 1352
rect 116176 1300 116182 1352
rect 111444 1244 112208 1272
rect 116688 1272 116716 1380
rect 126146 1368 126152 1420
rect 126204 1368 126210 1420
rect 128906 1368 128912 1420
rect 128964 1368 128970 1420
rect 132770 1368 132776 1420
rect 132828 1408 132834 1420
rect 133141 1411 133199 1417
rect 133141 1408 133153 1411
rect 132828 1380 133153 1408
rect 132828 1368 132834 1380
rect 133141 1377 133153 1380
rect 133187 1377 133199 1411
rect 133141 1371 133199 1377
rect 140222 1368 140228 1420
rect 140280 1408 140286 1420
rect 141513 1411 141571 1417
rect 140280 1380 140544 1408
rect 140280 1368 140286 1380
rect 116765 1343 116823 1349
rect 116765 1309 116777 1343
rect 116811 1340 116823 1343
rect 117498 1340 117504 1352
rect 116811 1312 117504 1340
rect 116811 1309 116823 1312
rect 116765 1303 116823 1309
rect 117498 1300 117504 1312
rect 117556 1300 117562 1352
rect 118050 1300 118056 1352
rect 118108 1300 118114 1352
rect 118694 1300 118700 1352
rect 118752 1300 118758 1352
rect 119338 1300 119344 1352
rect 119396 1300 119402 1352
rect 120350 1300 120356 1352
rect 120408 1300 120414 1352
rect 121086 1300 121092 1352
rect 121144 1300 121150 1352
rect 121638 1300 121644 1352
rect 121696 1300 121702 1352
rect 122466 1300 122472 1352
rect 122524 1300 122530 1352
rect 123202 1300 123208 1352
rect 123260 1300 123266 1352
rect 124217 1343 124275 1349
rect 124217 1309 124229 1343
rect 124263 1340 124275 1343
rect 125134 1340 125140 1352
rect 124263 1312 125140 1340
rect 124263 1309 124275 1312
rect 124217 1303 124275 1309
rect 125134 1300 125140 1312
rect 125192 1300 125198 1352
rect 125413 1343 125471 1349
rect 125413 1309 125425 1343
rect 125459 1340 125471 1343
rect 125778 1340 125784 1352
rect 125459 1312 125784 1340
rect 125459 1309 125471 1312
rect 125413 1303 125471 1309
rect 125778 1300 125784 1312
rect 125836 1300 125842 1352
rect 126333 1343 126391 1349
rect 126333 1309 126345 1343
rect 126379 1340 126391 1343
rect 126422 1340 126428 1352
rect 126379 1312 126428 1340
rect 126379 1309 126391 1312
rect 126333 1303 126391 1309
rect 126422 1300 126428 1312
rect 126480 1300 126486 1352
rect 127618 1300 127624 1352
rect 127676 1300 127682 1352
rect 129090 1300 129096 1352
rect 129148 1300 129154 1352
rect 130654 1300 130660 1352
rect 130712 1300 130718 1352
rect 131945 1343 132003 1349
rect 131945 1309 131957 1343
rect 131991 1340 132003 1343
rect 132678 1340 132684 1352
rect 131991 1312 132684 1340
rect 131991 1309 132003 1312
rect 131945 1303 132003 1309
rect 132678 1300 132684 1312
rect 132736 1300 132742 1352
rect 133325 1343 133383 1349
rect 133325 1309 133337 1343
rect 133371 1340 133383 1343
rect 133414 1340 133420 1352
rect 133371 1312 133420 1340
rect 133371 1309 133383 1312
rect 133325 1303 133383 1309
rect 133414 1300 133420 1312
rect 133472 1300 133478 1352
rect 134334 1300 134340 1352
rect 134392 1300 134398 1352
rect 138750 1300 138756 1352
rect 138808 1300 138814 1352
rect 138842 1300 138848 1352
rect 138900 1340 138906 1352
rect 139397 1343 139455 1349
rect 139397 1340 139409 1343
rect 138900 1312 139409 1340
rect 138900 1300 138906 1312
rect 139397 1309 139409 1312
rect 139443 1309 139455 1343
rect 139397 1303 139455 1309
rect 140317 1343 140375 1349
rect 140317 1309 140329 1343
rect 140363 1340 140375 1343
rect 140406 1340 140412 1352
rect 140363 1312 140412 1340
rect 140363 1309 140375 1312
rect 140317 1303 140375 1309
rect 140406 1300 140412 1312
rect 140464 1300 140470 1352
rect 140516 1349 140544 1380
rect 141513 1377 141525 1411
rect 141559 1408 141571 1411
rect 141694 1408 141700 1420
rect 141559 1380 141700 1408
rect 141559 1377 141571 1380
rect 141513 1371 141571 1377
rect 141694 1368 141700 1380
rect 141752 1368 141758 1420
rect 143368 1408 143396 1448
rect 143000 1380 143396 1408
rect 140501 1343 140559 1349
rect 140501 1309 140513 1343
rect 140547 1309 140559 1343
rect 140501 1303 140559 1309
rect 141234 1300 141240 1352
rect 141292 1300 141298 1352
rect 141418 1349 141424 1352
rect 141375 1343 141424 1349
rect 141375 1309 141387 1343
rect 141421 1309 141424 1343
rect 141375 1303 141424 1309
rect 141418 1300 141424 1303
rect 141476 1300 141482 1352
rect 142525 1343 142583 1349
rect 142525 1309 142537 1343
rect 142571 1340 142583 1343
rect 143000 1340 143028 1380
rect 143442 1368 143448 1420
rect 143500 1408 143506 1420
rect 143721 1411 143779 1417
rect 143721 1408 143733 1411
rect 143500 1380 143733 1408
rect 143500 1368 143506 1380
rect 143721 1377 143733 1380
rect 143767 1377 143779 1411
rect 143828 1408 143856 1448
rect 146294 1436 146300 1448
rect 146352 1436 146358 1488
rect 146386 1436 146392 1488
rect 146444 1476 146450 1488
rect 146941 1479 146999 1485
rect 146941 1476 146953 1479
rect 146444 1448 146953 1476
rect 146444 1436 146450 1448
rect 146941 1445 146953 1448
rect 146987 1445 146999 1479
rect 146941 1439 146999 1445
rect 148318 1436 148324 1488
rect 148376 1476 148382 1488
rect 148873 1479 148931 1485
rect 148873 1476 148885 1479
rect 148376 1448 148885 1476
rect 148376 1436 148382 1448
rect 148873 1445 148885 1448
rect 148919 1445 148931 1479
rect 149808 1476 149836 1516
rect 151262 1504 151268 1556
rect 151320 1544 151326 1556
rect 151449 1547 151507 1553
rect 151449 1544 151461 1547
rect 151320 1516 151461 1544
rect 151320 1504 151326 1516
rect 151449 1513 151461 1516
rect 151495 1513 151507 1547
rect 151449 1507 151507 1513
rect 151722 1504 151728 1556
rect 151780 1544 151786 1556
rect 153286 1544 153292 1556
rect 151780 1516 153292 1544
rect 151780 1504 151786 1516
rect 153286 1504 153292 1516
rect 153344 1504 153350 1556
rect 156322 1504 156328 1556
rect 156380 1544 156386 1556
rect 156785 1547 156843 1553
rect 156785 1544 156797 1547
rect 156380 1516 156797 1544
rect 156380 1504 156386 1516
rect 156785 1513 156797 1516
rect 156831 1513 156843 1547
rect 176930 1544 176936 1556
rect 156785 1507 156843 1513
rect 156984 1516 176936 1544
rect 156874 1476 156880 1488
rect 149808 1448 156880 1476
rect 148873 1439 148931 1445
rect 156874 1436 156880 1448
rect 156932 1436 156938 1488
rect 143828 1380 144132 1408
rect 143721 1371 143779 1377
rect 144104 1352 144132 1380
rect 144270 1368 144276 1420
rect 144328 1368 144334 1420
rect 145760 1380 145972 1408
rect 142571 1312 143028 1340
rect 142571 1309 142583 1312
rect 142525 1303 142583 1309
rect 143074 1300 143080 1352
rect 143132 1300 143138 1352
rect 143261 1343 143319 1349
rect 143261 1309 143273 1343
rect 143307 1309 143319 1343
rect 143261 1303 143319 1309
rect 117590 1272 117596 1284
rect 116688 1244 117596 1272
rect 109000 1232 109006 1244
rect 100812 1176 101352 1204
rect 101861 1207 101919 1213
rect 100812 1164 100818 1176
rect 101861 1173 101873 1207
rect 101907 1173 101919 1207
rect 101861 1167 101919 1173
rect 103514 1164 103520 1216
rect 103572 1164 103578 1216
rect 103790 1164 103796 1216
rect 103848 1164 103854 1216
rect 107378 1164 107384 1216
rect 107436 1204 107442 1216
rect 109589 1207 109647 1213
rect 109589 1204 109601 1207
rect 107436 1176 109601 1204
rect 107436 1164 107442 1176
rect 109589 1173 109601 1176
rect 109635 1173 109647 1207
rect 109589 1167 109647 1173
rect 110322 1164 110328 1216
rect 110380 1204 110386 1216
rect 111444 1204 111472 1244
rect 117590 1232 117596 1244
rect 117648 1232 117654 1284
rect 118418 1232 118424 1284
rect 118476 1272 118482 1284
rect 118476 1244 120948 1272
rect 118476 1232 118482 1244
rect 110380 1176 111472 1204
rect 110380 1164 110386 1176
rect 112162 1164 112168 1216
rect 112220 1204 112226 1216
rect 114005 1207 114063 1213
rect 114005 1204 114017 1207
rect 112220 1176 114017 1204
rect 112220 1164 112226 1176
rect 114005 1173 114017 1176
rect 114051 1173 114063 1207
rect 114005 1167 114063 1173
rect 114922 1164 114928 1216
rect 114980 1204 114986 1216
rect 117685 1207 117743 1213
rect 117685 1204 117697 1207
rect 114980 1176 117697 1204
rect 114980 1164 114986 1176
rect 117685 1173 117697 1176
rect 117731 1173 117743 1207
rect 117685 1167 117743 1173
rect 117869 1207 117927 1213
rect 117869 1173 117881 1207
rect 117915 1204 117927 1207
rect 117958 1204 117964 1216
rect 117915 1176 117964 1204
rect 117915 1173 117927 1176
rect 117869 1167 117927 1173
rect 117958 1164 117964 1176
rect 118016 1164 118022 1216
rect 118878 1164 118884 1216
rect 118936 1204 118942 1216
rect 120920 1213 120948 1244
rect 119157 1207 119215 1213
rect 119157 1204 119169 1207
rect 118936 1176 119169 1204
rect 118936 1164 118942 1176
rect 119157 1173 119169 1176
rect 119203 1173 119215 1207
rect 119157 1167 119215 1173
rect 120905 1207 120963 1213
rect 120905 1173 120917 1207
rect 120951 1173 120963 1207
rect 120905 1167 120963 1173
rect 121822 1164 121828 1216
rect 121880 1164 121886 1216
rect 122650 1164 122656 1216
rect 122708 1164 122714 1216
rect 123386 1164 123392 1216
rect 123444 1164 123450 1216
rect 124398 1164 124404 1216
rect 124456 1164 124462 1216
rect 125318 1164 125324 1216
rect 125376 1204 125382 1216
rect 125597 1207 125655 1213
rect 125597 1204 125609 1207
rect 125376 1176 125609 1204
rect 125376 1164 125382 1176
rect 125597 1173 125609 1176
rect 125643 1173 125655 1207
rect 125597 1167 125655 1173
rect 127802 1164 127808 1216
rect 127860 1164 127866 1216
rect 130838 1164 130844 1216
rect 130896 1164 130902 1216
rect 132126 1164 132132 1216
rect 132184 1164 132190 1216
rect 134518 1164 134524 1216
rect 134576 1164 134582 1216
rect 138382 1164 138388 1216
rect 138440 1204 138446 1216
rect 138569 1207 138627 1213
rect 138569 1204 138581 1207
rect 138440 1176 138581 1204
rect 138440 1164 138446 1176
rect 138569 1173 138581 1176
rect 138615 1173 138627 1207
rect 138569 1167 138627 1173
rect 139210 1164 139216 1216
rect 139268 1164 139274 1216
rect 143276 1204 143304 1303
rect 143994 1300 144000 1352
rect 144052 1300 144058 1352
rect 144086 1300 144092 1352
rect 144144 1349 144150 1352
rect 144144 1343 144172 1349
rect 144160 1309 144172 1343
rect 144144 1303 144172 1309
rect 144144 1300 144150 1303
rect 144914 1300 144920 1352
rect 144972 1340 144978 1352
rect 145760 1340 145788 1380
rect 144972 1312 145788 1340
rect 144972 1300 144978 1312
rect 145834 1300 145840 1352
rect 145892 1300 145898 1352
rect 145944 1340 145972 1380
rect 146202 1368 146208 1420
rect 146260 1408 146266 1420
rect 150158 1408 150164 1420
rect 146260 1380 146616 1408
rect 146260 1368 146266 1380
rect 146481 1343 146539 1349
rect 146481 1340 146493 1343
rect 145944 1312 146493 1340
rect 146481 1309 146493 1312
rect 146527 1309 146539 1343
rect 146588 1340 146616 1380
rect 149465 1380 150164 1408
rect 147125 1343 147183 1349
rect 147125 1340 147137 1343
rect 146588 1312 147137 1340
rect 146481 1303 146539 1309
rect 147125 1309 147137 1312
rect 147171 1309 147183 1343
rect 147125 1303 147183 1309
rect 148042 1300 148048 1352
rect 148100 1340 148106 1352
rect 148229 1343 148287 1349
rect 148229 1340 148241 1343
rect 148100 1312 148241 1340
rect 148100 1300 148106 1312
rect 148229 1309 148241 1312
rect 148275 1309 148287 1343
rect 148229 1303 148287 1309
rect 148413 1343 148471 1349
rect 148413 1309 148425 1343
rect 148459 1309 148471 1343
rect 148413 1303 148471 1309
rect 144748 1244 146340 1272
rect 144748 1204 144776 1244
rect 143276 1176 144776 1204
rect 144822 1164 144828 1216
rect 144880 1204 144886 1216
rect 146312 1213 146340 1244
rect 145653 1207 145711 1213
rect 145653 1204 145665 1207
rect 144880 1176 145665 1204
rect 144880 1164 144886 1176
rect 145653 1173 145665 1176
rect 145699 1173 145711 1207
rect 145653 1167 145711 1173
rect 146297 1207 146355 1213
rect 146297 1173 146309 1207
rect 146343 1173 146355 1207
rect 148428 1204 148456 1303
rect 149146 1300 149152 1352
rect 149204 1300 149210 1352
rect 149330 1349 149336 1352
rect 149287 1343 149336 1349
rect 149287 1309 149299 1343
rect 149333 1309 149336 1343
rect 149287 1303 149336 1309
rect 149330 1300 149336 1303
rect 149388 1300 149394 1352
rect 149465 1349 149493 1380
rect 150158 1368 150164 1380
rect 150216 1368 150222 1420
rect 150342 1368 150348 1420
rect 150400 1408 150406 1420
rect 150400 1380 151124 1408
rect 150400 1368 150406 1380
rect 149425 1343 149493 1349
rect 149425 1309 149437 1343
rect 149471 1312 149493 1343
rect 150069 1343 150127 1349
rect 149471 1309 149483 1312
rect 149425 1303 149483 1309
rect 150069 1309 150081 1343
rect 150115 1340 150127 1343
rect 150894 1340 150900 1352
rect 150115 1312 150900 1340
rect 150115 1309 150127 1312
rect 150069 1303 150127 1309
rect 150894 1300 150900 1312
rect 150952 1300 150958 1352
rect 150986 1300 150992 1352
rect 151044 1300 151050 1352
rect 151096 1340 151124 1380
rect 151538 1368 151544 1420
rect 151596 1408 151602 1420
rect 151596 1380 151768 1408
rect 151596 1368 151602 1380
rect 151633 1343 151691 1349
rect 151633 1340 151645 1343
rect 151096 1312 151645 1340
rect 151633 1309 151645 1312
rect 151679 1309 151691 1343
rect 151740 1340 151768 1380
rect 154574 1368 154580 1420
rect 154632 1408 154638 1420
rect 156984 1408 157012 1516
rect 176930 1504 176936 1516
rect 176988 1504 176994 1556
rect 177022 1504 177028 1556
rect 177080 1544 177086 1556
rect 211890 1544 211896 1556
rect 177080 1516 211896 1544
rect 177080 1504 177086 1516
rect 211890 1504 211896 1516
rect 211948 1504 211954 1556
rect 216582 1504 216588 1556
rect 216640 1544 216646 1556
rect 219434 1544 219440 1556
rect 216640 1516 219440 1544
rect 216640 1504 216646 1516
rect 219434 1504 219440 1516
rect 219492 1504 219498 1556
rect 219526 1504 219532 1556
rect 219584 1544 219590 1556
rect 220357 1547 220415 1553
rect 220357 1544 220369 1547
rect 219584 1516 220369 1544
rect 219584 1504 219590 1516
rect 220357 1513 220369 1516
rect 220403 1513 220415 1547
rect 220357 1507 220415 1513
rect 220446 1504 220452 1556
rect 220504 1544 220510 1556
rect 223022 1544 223028 1556
rect 220504 1516 223028 1544
rect 220504 1504 220510 1516
rect 223022 1504 223028 1516
rect 223080 1544 223086 1556
rect 223390 1544 223396 1556
rect 223080 1516 223396 1544
rect 223080 1504 223086 1516
rect 223390 1504 223396 1516
rect 223448 1544 223454 1556
rect 243538 1544 243544 1556
rect 223448 1516 230244 1544
rect 223448 1504 223454 1516
rect 157058 1436 157064 1488
rect 157116 1476 157122 1488
rect 178126 1476 178132 1488
rect 157116 1448 178132 1476
rect 157116 1436 157122 1448
rect 178126 1436 178132 1448
rect 178184 1436 178190 1488
rect 196158 1436 196164 1488
rect 196216 1476 196222 1488
rect 196621 1479 196679 1485
rect 196621 1476 196633 1479
rect 196216 1448 196633 1476
rect 196216 1436 196222 1448
rect 196621 1445 196633 1448
rect 196667 1445 196679 1479
rect 196621 1439 196679 1445
rect 198274 1436 198280 1488
rect 198332 1436 198338 1488
rect 203058 1436 203064 1488
rect 203116 1436 203122 1488
rect 209590 1436 209596 1488
rect 209648 1476 209654 1488
rect 210694 1476 210700 1488
rect 209648 1448 210700 1476
rect 209648 1436 209654 1448
rect 210694 1436 210700 1448
rect 210752 1436 210758 1488
rect 213012 1448 213224 1476
rect 154632 1380 157012 1408
rect 157168 1380 157380 1408
rect 154632 1368 154638 1380
rect 151740 1312 152228 1340
rect 151633 1303 151691 1309
rect 152200 1272 152228 1312
rect 152274 1300 152280 1352
rect 152332 1300 152338 1352
rect 153562 1300 153568 1352
rect 153620 1300 153626 1352
rect 154206 1300 154212 1352
rect 154264 1300 154270 1352
rect 154850 1300 154856 1352
rect 154908 1300 154914 1352
rect 156414 1300 156420 1352
rect 156472 1300 156478 1352
rect 156601 1343 156659 1349
rect 156601 1309 156613 1343
rect 156647 1340 156659 1343
rect 157168 1340 157196 1380
rect 156647 1312 157196 1340
rect 156647 1309 156659 1312
rect 156601 1303 156659 1309
rect 157242 1300 157248 1352
rect 157300 1300 157306 1352
rect 157352 1340 157380 1380
rect 158530 1368 158536 1420
rect 158588 1368 158594 1420
rect 159361 1411 159419 1417
rect 159361 1377 159373 1411
rect 159407 1408 159419 1411
rect 159450 1408 159456 1420
rect 159407 1380 159456 1408
rect 159407 1377 159419 1380
rect 159361 1371 159419 1377
rect 159450 1368 159456 1380
rect 159508 1368 159514 1420
rect 162578 1368 162584 1420
rect 162636 1408 162642 1420
rect 162673 1411 162731 1417
rect 162673 1408 162685 1411
rect 162636 1380 162685 1408
rect 162636 1368 162642 1380
rect 162673 1377 162685 1380
rect 162719 1377 162731 1411
rect 163130 1408 163136 1420
rect 162673 1371 162731 1377
rect 162780 1380 163136 1408
rect 157429 1343 157487 1349
rect 157429 1340 157441 1343
rect 157352 1312 157441 1340
rect 157429 1309 157441 1312
rect 157475 1340 157487 1343
rect 158717 1343 158775 1349
rect 158717 1340 158729 1343
rect 157475 1312 158729 1340
rect 157475 1309 157487 1312
rect 157429 1303 157487 1309
rect 158717 1309 158729 1312
rect 158763 1340 158775 1343
rect 159266 1340 159272 1352
rect 158763 1312 159272 1340
rect 158763 1309 158775 1312
rect 158717 1303 158775 1309
rect 159266 1300 159272 1312
rect 159324 1340 159330 1352
rect 159545 1343 159603 1349
rect 159545 1340 159557 1343
rect 159324 1312 159557 1340
rect 159324 1300 159330 1312
rect 159545 1309 159557 1312
rect 159591 1309 159603 1343
rect 159545 1303 159603 1309
rect 159729 1343 159787 1349
rect 159729 1309 159741 1343
rect 159775 1340 159787 1343
rect 160189 1343 160247 1349
rect 160189 1340 160201 1343
rect 159775 1312 160201 1340
rect 159775 1309 159787 1312
rect 159729 1303 159787 1309
rect 160189 1309 160201 1312
rect 160235 1309 160247 1343
rect 160189 1303 160247 1309
rect 161109 1343 161167 1349
rect 161109 1309 161121 1343
rect 161155 1340 161167 1343
rect 161474 1340 161480 1352
rect 161155 1312 161480 1340
rect 161155 1309 161167 1312
rect 161109 1303 161167 1309
rect 161474 1300 161480 1312
rect 161532 1300 161538 1352
rect 161937 1343 161995 1349
rect 161937 1309 161949 1343
rect 161983 1340 161995 1343
rect 162780 1340 162808 1380
rect 163130 1368 163136 1380
rect 163188 1368 163194 1420
rect 166902 1368 166908 1420
rect 166960 1368 166966 1420
rect 166994 1368 167000 1420
rect 167052 1408 167058 1420
rect 169846 1408 169852 1420
rect 167052 1380 169852 1408
rect 167052 1368 167058 1380
rect 169846 1368 169852 1380
rect 169904 1368 169910 1420
rect 171686 1368 171692 1420
rect 171744 1368 171750 1420
rect 190641 1411 190699 1417
rect 190641 1377 190653 1411
rect 190687 1408 190699 1411
rect 190917 1411 190975 1417
rect 190917 1408 190929 1411
rect 190687 1380 190929 1408
rect 190687 1377 190699 1380
rect 190641 1371 190699 1377
rect 190917 1377 190929 1380
rect 190963 1408 190975 1411
rect 191374 1408 191380 1420
rect 190963 1380 191380 1408
rect 190963 1377 190975 1380
rect 190917 1371 190975 1377
rect 191374 1368 191380 1380
rect 191432 1368 191438 1420
rect 196250 1368 196256 1420
rect 196308 1368 196314 1420
rect 197906 1368 197912 1420
rect 197964 1368 197970 1420
rect 201310 1368 201316 1420
rect 201368 1368 201374 1420
rect 202877 1411 202935 1417
rect 202877 1377 202889 1411
rect 202923 1408 202935 1411
rect 203076 1408 203104 1436
rect 202923 1380 203104 1408
rect 202923 1377 202935 1380
rect 202877 1371 202935 1377
rect 205818 1368 205824 1420
rect 205876 1368 205882 1420
rect 210142 1368 210148 1420
rect 210200 1408 210206 1420
rect 211249 1411 211307 1417
rect 211249 1408 211261 1411
rect 210200 1380 211261 1408
rect 210200 1368 210206 1380
rect 211249 1377 211261 1380
rect 211295 1408 211307 1411
rect 213012 1408 213040 1448
rect 211295 1380 213040 1408
rect 211295 1377 211307 1380
rect 211249 1371 211307 1377
rect 213086 1368 213092 1420
rect 213144 1368 213150 1420
rect 213196 1408 213224 1448
rect 217962 1436 217968 1488
rect 218020 1476 218026 1488
rect 220630 1476 220636 1488
rect 218020 1448 220636 1476
rect 218020 1436 218026 1448
rect 220630 1436 220636 1448
rect 220688 1436 220694 1488
rect 220722 1436 220728 1488
rect 220780 1476 220786 1488
rect 229830 1476 229836 1488
rect 220780 1448 229836 1476
rect 220780 1436 220786 1448
rect 229830 1436 229836 1448
rect 229888 1436 229894 1488
rect 213641 1411 213699 1417
rect 213641 1408 213653 1411
rect 213196 1380 213653 1408
rect 213641 1377 213653 1380
rect 213687 1408 213699 1411
rect 213822 1408 213828 1420
rect 213687 1380 213828 1408
rect 213687 1377 213699 1380
rect 213641 1371 213699 1377
rect 213822 1368 213828 1380
rect 213880 1368 213886 1420
rect 215570 1368 215576 1420
rect 215628 1408 215634 1420
rect 215849 1411 215907 1417
rect 215849 1408 215861 1411
rect 215628 1380 215861 1408
rect 215628 1368 215634 1380
rect 215849 1377 215861 1380
rect 215895 1408 215907 1411
rect 218146 1408 218152 1420
rect 215895 1380 218152 1408
rect 215895 1377 215907 1380
rect 215849 1371 215907 1377
rect 218146 1368 218152 1380
rect 218204 1368 218210 1420
rect 218330 1368 218336 1420
rect 218388 1408 218394 1420
rect 222010 1408 222016 1420
rect 218388 1380 222016 1408
rect 218388 1368 218394 1380
rect 222010 1368 222016 1380
rect 222068 1368 222074 1420
rect 224402 1368 224408 1420
rect 224460 1368 224466 1420
rect 226889 1411 226947 1417
rect 226889 1377 226901 1411
rect 226935 1408 226947 1411
rect 227162 1408 227168 1420
rect 226935 1380 227168 1408
rect 226935 1377 226947 1380
rect 226889 1371 226947 1377
rect 227162 1368 227168 1380
rect 227220 1368 227226 1420
rect 227254 1368 227260 1420
rect 227312 1368 227318 1420
rect 161983 1312 162808 1340
rect 161983 1309 161995 1312
rect 161937 1303 161995 1309
rect 162854 1300 162860 1352
rect 162912 1300 162918 1352
rect 163041 1343 163099 1349
rect 163041 1309 163053 1343
rect 163087 1340 163099 1343
rect 163685 1343 163743 1349
rect 163685 1340 163697 1343
rect 163087 1312 163697 1340
rect 163087 1309 163099 1312
rect 163041 1303 163099 1309
rect 163685 1309 163697 1312
rect 163731 1309 163743 1343
rect 163685 1303 163743 1309
rect 164418 1300 164424 1352
rect 164476 1300 164482 1352
rect 167089 1343 167147 1349
rect 167089 1309 167101 1343
rect 167135 1340 167147 1343
rect 167178 1340 167184 1352
rect 167135 1312 167184 1340
rect 167135 1309 167147 1312
rect 167089 1303 167147 1309
rect 167178 1300 167184 1312
rect 167236 1300 167242 1352
rect 167273 1343 167331 1349
rect 167273 1309 167285 1343
rect 167319 1340 167331 1343
rect 167733 1343 167791 1349
rect 167733 1340 167745 1343
rect 167319 1312 167745 1340
rect 167319 1309 167331 1312
rect 167273 1303 167331 1309
rect 167733 1309 167745 1312
rect 167779 1309 167791 1343
rect 167733 1303 167791 1309
rect 168190 1300 168196 1352
rect 168248 1340 168254 1352
rect 168837 1343 168895 1349
rect 168837 1340 168849 1343
rect 168248 1312 168849 1340
rect 168248 1300 168254 1312
rect 168837 1309 168849 1312
rect 168883 1309 168895 1343
rect 168837 1303 168895 1309
rect 172238 1300 172244 1352
rect 172296 1300 172302 1352
rect 172514 1300 172520 1352
rect 172572 1300 172578 1352
rect 173894 1300 173900 1352
rect 173952 1340 173958 1352
rect 173989 1343 174047 1349
rect 173989 1340 174001 1343
rect 173952 1312 174001 1340
rect 173952 1300 173958 1312
rect 173989 1309 174001 1312
rect 174035 1309 174047 1343
rect 173989 1303 174047 1309
rect 174262 1300 174268 1352
rect 174320 1300 174326 1352
rect 175274 1300 175280 1352
rect 175332 1340 175338 1352
rect 176565 1343 176623 1349
rect 176565 1340 176577 1343
rect 175332 1312 176577 1340
rect 175332 1300 175338 1312
rect 176565 1309 176577 1312
rect 176611 1309 176623 1343
rect 176565 1303 176623 1309
rect 176838 1300 176844 1352
rect 176896 1300 176902 1352
rect 178494 1300 178500 1352
rect 178552 1340 178558 1352
rect 179141 1343 179199 1349
rect 179141 1340 179153 1343
rect 178552 1312 179153 1340
rect 178552 1300 178558 1312
rect 179141 1309 179153 1312
rect 179187 1309 179199 1343
rect 179141 1303 179199 1309
rect 179414 1300 179420 1352
rect 179472 1300 179478 1352
rect 180334 1300 180340 1352
rect 180392 1340 180398 1352
rect 181717 1343 181775 1349
rect 181717 1340 181729 1343
rect 180392 1312 181729 1340
rect 180392 1300 180398 1312
rect 181717 1309 181729 1312
rect 181763 1309 181775 1343
rect 181717 1303 181775 1309
rect 181990 1300 181996 1352
rect 182048 1300 182054 1352
rect 183278 1300 183284 1352
rect 183336 1340 183342 1352
rect 184293 1343 184351 1349
rect 184293 1340 184305 1343
rect 183336 1312 184305 1340
rect 183336 1300 183342 1312
rect 184293 1309 184305 1312
rect 184339 1309 184351 1343
rect 184293 1303 184351 1309
rect 184566 1300 184572 1352
rect 184624 1300 184630 1352
rect 185486 1300 185492 1352
rect 185544 1340 185550 1352
rect 186869 1343 186927 1349
rect 186869 1340 186881 1343
rect 185544 1312 186881 1340
rect 185544 1300 185550 1312
rect 186869 1309 186881 1312
rect 186915 1309 186927 1343
rect 186869 1303 186927 1309
rect 187142 1300 187148 1352
rect 187200 1300 187206 1352
rect 188614 1300 188620 1352
rect 188672 1300 188678 1352
rect 189442 1300 189448 1352
rect 189500 1300 189506 1352
rect 189718 1300 189724 1352
rect 189776 1300 189782 1352
rect 191006 1300 191012 1352
rect 191064 1340 191070 1352
rect 191101 1343 191159 1349
rect 191101 1340 191113 1343
rect 191064 1312 191113 1340
rect 191064 1300 191070 1312
rect 191101 1309 191113 1312
rect 191147 1309 191159 1343
rect 191101 1303 191159 1309
rect 191282 1300 191288 1352
rect 191340 1300 191346 1352
rect 192389 1343 192447 1349
rect 192389 1309 192401 1343
rect 192435 1309 192447 1343
rect 192389 1303 192447 1309
rect 193125 1343 193183 1349
rect 193125 1309 193137 1343
rect 193171 1340 193183 1343
rect 194042 1340 194048 1352
rect 193171 1312 194048 1340
rect 193171 1309 193183 1312
rect 193125 1303 193183 1309
rect 149900 1244 150940 1272
rect 152200 1244 152320 1272
rect 149900 1204 149928 1244
rect 148428 1176 149928 1204
rect 146297 1167 146355 1173
rect 150802 1164 150808 1216
rect 150860 1164 150866 1216
rect 150912 1204 150940 1244
rect 152093 1207 152151 1213
rect 152093 1204 152105 1207
rect 150912 1176 152105 1204
rect 152093 1173 152105 1176
rect 152139 1173 152151 1207
rect 152292 1204 152320 1244
rect 152366 1232 152372 1284
rect 152424 1272 152430 1284
rect 154942 1272 154948 1284
rect 152424 1244 154948 1272
rect 152424 1232 152430 1244
rect 154942 1232 154948 1244
rect 155000 1232 155006 1284
rect 155586 1232 155592 1284
rect 155644 1272 155650 1284
rect 157613 1275 157671 1281
rect 157613 1272 157625 1275
rect 155644 1244 157625 1272
rect 155644 1232 155650 1244
rect 157613 1241 157625 1244
rect 157659 1241 157671 1275
rect 157613 1235 157671 1241
rect 157702 1232 157708 1284
rect 157760 1272 157766 1284
rect 158901 1275 158959 1281
rect 158901 1272 158913 1275
rect 157760 1244 158913 1272
rect 157760 1232 157766 1244
rect 158901 1241 158913 1244
rect 158947 1241 158959 1275
rect 192404 1272 192432 1303
rect 194042 1300 194048 1312
rect 194100 1300 194106 1352
rect 194594 1300 194600 1352
rect 194652 1300 194658 1352
rect 195425 1343 195483 1349
rect 195425 1309 195437 1343
rect 195471 1340 195483 1343
rect 196066 1340 196072 1352
rect 195471 1312 196072 1340
rect 195471 1309 195483 1312
rect 195425 1303 195483 1309
rect 196066 1300 196072 1312
rect 196124 1300 196130 1352
rect 196434 1300 196440 1352
rect 196492 1300 196498 1352
rect 198093 1343 198151 1349
rect 198093 1309 198105 1343
rect 198139 1340 198151 1343
rect 198366 1340 198372 1352
rect 198139 1312 198372 1340
rect 198139 1309 198151 1312
rect 198093 1303 198151 1309
rect 198366 1300 198372 1312
rect 198424 1300 198430 1352
rect 199749 1343 199807 1349
rect 199749 1309 199761 1343
rect 199795 1340 199807 1343
rect 200574 1340 200580 1352
rect 199795 1312 200580 1340
rect 199795 1309 199807 1312
rect 199749 1303 199807 1309
rect 200574 1300 200580 1312
rect 200632 1300 200638 1352
rect 201494 1300 201500 1352
rect 201552 1340 201558 1352
rect 203061 1343 203119 1349
rect 203061 1340 203073 1343
rect 201552 1312 203073 1340
rect 201552 1300 201558 1312
rect 203061 1309 203073 1312
rect 203107 1309 203119 1343
rect 203061 1303 203119 1309
rect 203245 1343 203303 1349
rect 203245 1309 203257 1343
rect 203291 1340 203303 1343
rect 203705 1343 203763 1349
rect 203705 1340 203717 1343
rect 203291 1312 203717 1340
rect 203291 1309 203303 1312
rect 203245 1303 203303 1309
rect 203705 1309 203717 1312
rect 203751 1309 203763 1343
rect 203705 1303 203763 1309
rect 206554 1300 206560 1352
rect 206612 1300 206618 1352
rect 207658 1300 207664 1352
rect 207716 1300 207722 1352
rect 208302 1300 208308 1352
rect 208360 1300 208366 1352
rect 208946 1300 208952 1352
rect 209004 1300 209010 1352
rect 210050 1300 210056 1352
rect 210108 1300 210114 1352
rect 210234 1300 210240 1352
rect 210292 1300 210298 1352
rect 210970 1300 210976 1352
rect 211028 1300 211034 1352
rect 211062 1300 211068 1352
rect 211120 1349 211126 1352
rect 211120 1343 211148 1349
rect 211136 1309 211148 1343
rect 211120 1303 211148 1309
rect 211120 1300 211126 1303
rect 212442 1300 212448 1352
rect 212500 1300 212506 1352
rect 212626 1300 212632 1352
rect 212684 1300 212690 1352
rect 213362 1300 213368 1352
rect 213420 1300 213426 1352
rect 213546 1349 213552 1352
rect 213503 1343 213552 1349
rect 213503 1309 213515 1343
rect 213549 1309 213552 1343
rect 213503 1303 213552 1309
rect 213546 1300 213552 1303
rect 213604 1300 213610 1352
rect 215018 1300 215024 1352
rect 215076 1340 215082 1352
rect 215205 1343 215263 1349
rect 215205 1340 215217 1343
rect 215076 1312 215217 1340
rect 215076 1300 215082 1312
rect 215205 1309 215217 1312
rect 215251 1309 215263 1343
rect 215205 1303 215263 1309
rect 215389 1343 215447 1349
rect 215389 1309 215401 1343
rect 215435 1309 215447 1343
rect 215389 1303 215447 1309
rect 193214 1272 193220 1284
rect 192404 1244 193220 1272
rect 158901 1235 158959 1241
rect 193214 1232 193220 1244
rect 193272 1232 193278 1284
rect 201034 1232 201040 1284
rect 201092 1272 201098 1284
rect 201681 1275 201739 1281
rect 201681 1272 201693 1275
rect 201092 1244 201693 1272
rect 201092 1232 201098 1244
rect 201681 1241 201693 1244
rect 201727 1241 201739 1275
rect 208394 1272 208400 1284
rect 201681 1235 201739 1241
rect 207492 1244 208400 1272
rect 153381 1207 153439 1213
rect 153381 1204 153393 1207
rect 152292 1176 153393 1204
rect 152093 1167 152151 1173
rect 153381 1173 153393 1176
rect 153427 1173 153439 1207
rect 153381 1167 153439 1173
rect 153930 1164 153936 1216
rect 153988 1204 153994 1216
rect 154025 1207 154083 1213
rect 154025 1204 154037 1207
rect 153988 1176 154037 1204
rect 153988 1164 153994 1176
rect 154025 1173 154037 1176
rect 154071 1173 154083 1207
rect 154025 1167 154083 1173
rect 154666 1164 154672 1216
rect 154724 1164 154730 1216
rect 160094 1164 160100 1216
rect 160152 1204 160158 1216
rect 160373 1207 160431 1213
rect 160373 1204 160385 1207
rect 160152 1176 160385 1204
rect 160152 1164 160158 1176
rect 160373 1173 160385 1176
rect 160419 1173 160431 1207
rect 160373 1167 160431 1173
rect 161290 1164 161296 1216
rect 161348 1164 161354 1216
rect 162118 1164 162124 1216
rect 162176 1164 162182 1216
rect 163498 1164 163504 1216
rect 163556 1204 163562 1216
rect 163869 1207 163927 1213
rect 163869 1204 163881 1207
rect 163556 1176 163881 1204
rect 163556 1164 163562 1176
rect 163869 1173 163881 1176
rect 163915 1173 163927 1207
rect 163869 1167 163927 1173
rect 164602 1164 164608 1216
rect 164660 1164 164666 1216
rect 167914 1164 167920 1216
rect 167972 1164 167978 1216
rect 169018 1164 169024 1216
rect 169076 1164 169082 1216
rect 187602 1164 187608 1216
rect 187660 1204 187666 1216
rect 188433 1207 188491 1213
rect 188433 1204 188445 1207
rect 187660 1176 188445 1204
rect 187660 1164 187666 1176
rect 188433 1173 188445 1176
rect 188479 1173 188491 1207
rect 188433 1167 188491 1173
rect 192570 1164 192576 1216
rect 192628 1164 192634 1216
rect 192846 1164 192852 1216
rect 192904 1204 192910 1216
rect 193309 1207 193367 1213
rect 193309 1204 193321 1207
rect 192904 1176 193321 1204
rect 192904 1164 192910 1176
rect 193309 1173 193321 1176
rect 193355 1173 193367 1207
rect 193309 1167 193367 1173
rect 193582 1164 193588 1216
rect 193640 1204 193646 1216
rect 194781 1207 194839 1213
rect 194781 1204 194793 1207
rect 193640 1176 194793 1204
rect 193640 1164 193646 1176
rect 194781 1173 194793 1176
rect 194827 1173 194839 1207
rect 194781 1167 194839 1173
rect 195606 1164 195612 1216
rect 195664 1164 195670 1216
rect 199930 1164 199936 1216
rect 199988 1164 199994 1216
rect 202414 1164 202420 1216
rect 202472 1204 202478 1216
rect 203889 1207 203947 1213
rect 203889 1204 203901 1207
rect 202472 1176 203901 1204
rect 202472 1164 202478 1176
rect 203889 1173 203901 1176
rect 203935 1173 203947 1207
rect 203889 1167 203947 1173
rect 206373 1207 206431 1213
rect 206373 1173 206385 1207
rect 206419 1204 206431 1207
rect 207106 1204 207112 1216
rect 206419 1176 207112 1204
rect 206419 1173 206431 1176
rect 206373 1167 206431 1173
rect 207106 1164 207112 1176
rect 207164 1164 207170 1216
rect 207492 1213 207520 1244
rect 208394 1232 208400 1244
rect 208452 1232 208458 1284
rect 209038 1232 209044 1284
rect 209096 1272 209102 1284
rect 209096 1244 209774 1272
rect 209096 1232 209102 1244
rect 207477 1207 207535 1213
rect 207477 1173 207489 1207
rect 207523 1173 207535 1207
rect 207477 1167 207535 1173
rect 207566 1164 207572 1216
rect 207624 1204 207630 1216
rect 208121 1207 208179 1213
rect 208121 1204 208133 1207
rect 207624 1176 208133 1204
rect 207624 1164 207630 1176
rect 208121 1173 208133 1176
rect 208167 1173 208179 1207
rect 208121 1167 208179 1173
rect 208765 1207 208823 1213
rect 208765 1173 208777 1207
rect 208811 1204 208823 1207
rect 209130 1204 209136 1216
rect 208811 1176 209136 1204
rect 208811 1173 208823 1176
rect 208765 1167 208823 1173
rect 209130 1164 209136 1176
rect 209188 1164 209194 1216
rect 209498 1164 209504 1216
rect 209556 1164 209562 1216
rect 209746 1204 209774 1244
rect 211893 1207 211951 1213
rect 211893 1204 211905 1207
rect 209746 1176 211905 1204
rect 211893 1173 211905 1176
rect 211939 1173 211951 1207
rect 211893 1167 211951 1173
rect 212350 1164 212356 1216
rect 212408 1204 212414 1216
rect 214285 1207 214343 1213
rect 214285 1204 214297 1207
rect 212408 1176 214297 1204
rect 212408 1164 212414 1176
rect 214285 1173 214297 1176
rect 214331 1173 214343 1207
rect 214285 1167 214343 1173
rect 214650 1164 214656 1216
rect 214708 1164 214714 1216
rect 215404 1204 215432 1303
rect 216122 1300 216128 1352
rect 216180 1300 216186 1352
rect 216306 1349 216312 1352
rect 216263 1343 216312 1349
rect 216263 1309 216275 1343
rect 216309 1309 216312 1343
rect 216263 1303 216312 1309
rect 216306 1300 216312 1303
rect 216364 1300 216370 1352
rect 216398 1300 216404 1352
rect 216456 1300 216462 1352
rect 217870 1300 217876 1352
rect 217928 1300 217934 1352
rect 217962 1300 217968 1352
rect 218020 1300 218026 1352
rect 218054 1300 218060 1352
rect 218112 1300 218118 1352
rect 218238 1300 218244 1352
rect 218296 1340 218302 1352
rect 218885 1343 218943 1349
rect 218885 1340 218897 1343
rect 218296 1312 218897 1340
rect 218296 1300 218302 1312
rect 218885 1309 218897 1312
rect 218931 1309 218943 1343
rect 218885 1303 218943 1309
rect 219526 1300 219532 1352
rect 219584 1300 219590 1352
rect 220538 1300 220544 1352
rect 220596 1300 220602 1352
rect 221458 1300 221464 1352
rect 221516 1340 221522 1352
rect 221645 1343 221703 1349
rect 221645 1340 221657 1343
rect 221516 1312 221657 1340
rect 221516 1300 221522 1312
rect 221645 1309 221657 1312
rect 221691 1309 221703 1343
rect 221645 1303 221703 1309
rect 221734 1300 221740 1352
rect 221792 1300 221798 1352
rect 221921 1343 221979 1349
rect 221921 1309 221933 1343
rect 221967 1309 221979 1343
rect 221921 1303 221979 1309
rect 216876 1244 219388 1272
rect 216876 1204 216904 1244
rect 215404 1176 216904 1204
rect 217042 1164 217048 1216
rect 217100 1164 217106 1216
rect 218241 1207 218299 1213
rect 218241 1173 218253 1207
rect 218287 1204 218299 1207
rect 218422 1204 218428 1216
rect 218287 1176 218428 1204
rect 218287 1173 218299 1176
rect 218241 1167 218299 1173
rect 218422 1164 218428 1176
rect 218480 1164 218486 1216
rect 218698 1164 218704 1216
rect 218756 1164 218762 1216
rect 219360 1213 219388 1244
rect 220814 1232 220820 1284
rect 220872 1272 220878 1284
rect 221936 1272 221964 1303
rect 223114 1300 223120 1352
rect 223172 1300 223178 1352
rect 223942 1300 223948 1352
rect 224000 1340 224006 1352
rect 224221 1343 224279 1349
rect 224221 1340 224233 1343
rect 224000 1312 224233 1340
rect 224000 1300 224006 1312
rect 224221 1309 224233 1312
rect 224267 1309 224279 1343
rect 224221 1303 224279 1309
rect 225506 1300 225512 1352
rect 225564 1300 225570 1352
rect 226426 1300 226432 1352
rect 226484 1300 226490 1352
rect 227070 1300 227076 1352
rect 227128 1300 227134 1352
rect 228542 1300 228548 1352
rect 228600 1300 228606 1352
rect 229281 1343 229339 1349
rect 229281 1309 229293 1343
rect 229327 1340 229339 1343
rect 230106 1340 230112 1352
rect 229327 1312 230112 1340
rect 229327 1309 229339 1312
rect 229281 1303 229339 1309
rect 230106 1300 230112 1312
rect 230164 1300 230170 1352
rect 230216 1340 230244 1516
rect 230676 1516 243544 1544
rect 230290 1368 230296 1420
rect 230348 1408 230354 1420
rect 230676 1408 230704 1516
rect 243538 1504 243544 1516
rect 243596 1504 243602 1556
rect 246574 1504 246580 1556
rect 246632 1544 246638 1556
rect 247313 1547 247371 1553
rect 247313 1544 247325 1547
rect 246632 1516 247325 1544
rect 246632 1504 246638 1516
rect 247313 1513 247325 1516
rect 247359 1513 247371 1547
rect 247313 1507 247371 1513
rect 253106 1504 253112 1556
rect 253164 1544 253170 1556
rect 269850 1544 269856 1556
rect 253164 1516 269856 1544
rect 253164 1504 253170 1516
rect 269850 1504 269856 1516
rect 269908 1504 269914 1556
rect 230348 1380 230704 1408
rect 230860 1448 249104 1476
rect 230348 1368 230354 1380
rect 230860 1340 230888 1448
rect 231302 1368 231308 1420
rect 231360 1368 231366 1420
rect 235813 1411 235871 1417
rect 235813 1377 235825 1411
rect 235859 1408 235871 1411
rect 235902 1408 235908 1420
rect 235859 1380 235908 1408
rect 235859 1377 235871 1380
rect 235813 1371 235871 1377
rect 235902 1368 235908 1380
rect 235960 1368 235966 1420
rect 239950 1368 239956 1420
rect 240008 1368 240014 1420
rect 246117 1411 246175 1417
rect 246117 1377 246129 1411
rect 246163 1377 246175 1411
rect 246117 1371 246175 1377
rect 247497 1411 247555 1417
rect 247497 1377 247509 1411
rect 247543 1408 247555 1411
rect 247678 1408 247684 1420
rect 247543 1380 247684 1408
rect 247543 1377 247555 1380
rect 247497 1371 247555 1377
rect 230216 1312 230888 1340
rect 231486 1300 231492 1352
rect 231544 1300 231550 1352
rect 231673 1343 231731 1349
rect 231673 1309 231685 1343
rect 231719 1340 231731 1343
rect 232133 1343 232191 1349
rect 232133 1340 232145 1343
rect 231719 1312 232145 1340
rect 231719 1309 231731 1312
rect 231673 1303 231731 1309
rect 232133 1309 232145 1312
rect 232179 1309 232191 1343
rect 232133 1303 232191 1309
rect 233694 1300 233700 1352
rect 233752 1300 233758 1352
rect 234433 1343 234491 1349
rect 234433 1309 234445 1343
rect 234479 1340 234491 1343
rect 235258 1340 235264 1352
rect 234479 1312 235264 1340
rect 234479 1309 234491 1312
rect 234433 1303 234491 1309
rect 235258 1300 235264 1312
rect 235316 1300 235322 1352
rect 235994 1300 236000 1352
rect 236052 1300 236058 1352
rect 236181 1343 236239 1349
rect 236181 1309 236193 1343
rect 236227 1340 236239 1343
rect 236641 1343 236699 1349
rect 236641 1340 236653 1343
rect 236227 1312 236653 1340
rect 236227 1309 236239 1312
rect 236181 1303 236239 1309
rect 236641 1309 236653 1312
rect 236687 1309 236699 1343
rect 236641 1303 236699 1309
rect 240962 1300 240968 1352
rect 241020 1300 241026 1352
rect 241054 1300 241060 1352
rect 241112 1340 241118 1352
rect 241241 1343 241299 1349
rect 241241 1340 241253 1343
rect 241112 1312 241253 1340
rect 241112 1300 241118 1312
rect 241241 1309 241253 1312
rect 241287 1309 241299 1343
rect 241241 1303 241299 1309
rect 241974 1300 241980 1352
rect 242032 1340 242038 1352
rect 243541 1343 243599 1349
rect 243541 1340 243553 1343
rect 242032 1312 243553 1340
rect 242032 1300 242038 1312
rect 243541 1309 243553 1312
rect 243587 1309 243599 1343
rect 243541 1303 243599 1309
rect 243814 1300 243820 1352
rect 243872 1300 243878 1352
rect 245473 1343 245531 1349
rect 245473 1309 245485 1343
rect 245519 1340 245531 1343
rect 246022 1340 246028 1352
rect 245519 1312 246028 1340
rect 245519 1309 245531 1312
rect 245473 1303 245531 1309
rect 246022 1300 246028 1312
rect 246080 1300 246086 1352
rect 220872 1244 221964 1272
rect 222289 1275 222347 1281
rect 220872 1232 220878 1244
rect 222289 1241 222301 1275
rect 222335 1272 222347 1275
rect 225322 1272 225328 1284
rect 222335 1244 225328 1272
rect 222335 1241 222347 1244
rect 222289 1235 222347 1241
rect 225322 1232 225328 1244
rect 225380 1232 225386 1284
rect 244366 1272 244372 1284
rect 226536 1244 244372 1272
rect 219345 1207 219403 1213
rect 219345 1173 219357 1207
rect 219391 1173 219403 1207
rect 219345 1167 219403 1173
rect 222930 1164 222936 1216
rect 222988 1164 222994 1216
rect 224770 1164 224776 1216
rect 224828 1204 224834 1216
rect 225693 1207 225751 1213
rect 225693 1204 225705 1207
rect 224828 1176 225705 1204
rect 224828 1164 224834 1176
rect 225693 1173 225705 1176
rect 225739 1173 225751 1207
rect 225693 1167 225751 1173
rect 226242 1164 226248 1216
rect 226300 1164 226306 1216
rect 226334 1164 226340 1216
rect 226392 1204 226398 1216
rect 226536 1204 226564 1244
rect 244366 1232 244372 1244
rect 244424 1232 244430 1284
rect 244918 1232 244924 1284
rect 244976 1272 244982 1284
rect 246132 1272 246160 1371
rect 247678 1368 247684 1380
rect 247736 1368 247742 1420
rect 249076 1408 249104 1448
rect 250530 1436 250536 1488
rect 250588 1476 250594 1488
rect 268838 1476 268844 1488
rect 250588 1448 268844 1476
rect 250588 1436 250594 1448
rect 268838 1436 268844 1448
rect 268896 1436 268902 1488
rect 257706 1408 257712 1420
rect 249076 1380 257712 1408
rect 257706 1368 257712 1380
rect 257764 1368 257770 1420
rect 257908 1380 258304 1408
rect 246390 1300 246396 1352
rect 246448 1300 246454 1352
rect 247218 1300 247224 1352
rect 247276 1340 247282 1352
rect 247313 1343 247371 1349
rect 247313 1340 247325 1343
rect 247276 1312 247325 1340
rect 247276 1300 247282 1312
rect 247313 1309 247325 1312
rect 247359 1309 247371 1343
rect 247313 1303 247371 1309
rect 247586 1300 247592 1352
rect 247644 1300 247650 1352
rect 248785 1343 248843 1349
rect 248785 1340 248797 1343
rect 248064 1312 248797 1340
rect 244976 1244 246160 1272
rect 244976 1232 244982 1244
rect 246206 1232 246212 1284
rect 246264 1272 246270 1284
rect 246264 1244 246436 1272
rect 246264 1232 246270 1244
rect 226392 1176 226564 1204
rect 226392 1164 226398 1176
rect 228726 1164 228732 1216
rect 228784 1164 228790 1216
rect 229462 1164 229468 1216
rect 229520 1164 229526 1216
rect 231854 1164 231860 1216
rect 231912 1204 231918 1216
rect 232317 1207 232375 1213
rect 232317 1204 232329 1207
rect 231912 1176 232329 1204
rect 231912 1164 231918 1176
rect 232317 1173 232329 1176
rect 232363 1173 232375 1207
rect 232317 1167 232375 1173
rect 233878 1164 233884 1216
rect 233936 1164 233942 1216
rect 234614 1164 234620 1216
rect 234672 1164 234678 1216
rect 235810 1164 235816 1216
rect 235868 1204 235874 1216
rect 236825 1207 236883 1213
rect 236825 1204 236837 1207
rect 235868 1176 236837 1204
rect 235868 1164 235874 1176
rect 236825 1173 236837 1176
rect 236871 1173 236883 1207
rect 236825 1167 236883 1173
rect 245289 1207 245347 1213
rect 245289 1173 245301 1207
rect 245335 1204 245347 1207
rect 246298 1204 246304 1216
rect 245335 1176 246304 1204
rect 245335 1173 245347 1176
rect 245289 1167 245347 1173
rect 246298 1164 246304 1176
rect 246356 1164 246362 1216
rect 246408 1204 246436 1244
rect 248064 1216 248092 1312
rect 248785 1309 248797 1312
rect 248831 1309 248843 1343
rect 251269 1343 251327 1349
rect 251269 1340 251281 1343
rect 248785 1303 248843 1309
rect 250180 1312 251281 1340
rect 248966 1232 248972 1284
rect 249024 1232 249030 1284
rect 247773 1207 247831 1213
rect 247773 1204 247785 1207
rect 246408 1176 247785 1204
rect 247773 1173 247785 1176
rect 247819 1173 247831 1207
rect 247773 1167 247831 1173
rect 248046 1164 248052 1216
rect 248104 1164 248110 1216
rect 248414 1164 248420 1216
rect 248472 1204 248478 1216
rect 250180 1204 250208 1312
rect 251269 1309 251281 1312
rect 251315 1309 251327 1343
rect 251269 1303 251327 1309
rect 251542 1300 251548 1352
rect 251600 1300 251606 1352
rect 252738 1300 252744 1352
rect 252796 1300 252802 1352
rect 252830 1300 252836 1352
rect 252888 1340 252894 1352
rect 253845 1343 253903 1349
rect 253845 1340 253857 1343
rect 252888 1312 253857 1340
rect 252888 1300 252894 1312
rect 253845 1309 253857 1312
rect 253891 1309 253903 1343
rect 253845 1303 253903 1309
rect 254118 1300 254124 1352
rect 254176 1300 254182 1352
rect 255590 1300 255596 1352
rect 255648 1300 255654 1352
rect 255958 1300 255964 1352
rect 256016 1340 256022 1352
rect 256421 1343 256479 1349
rect 256421 1340 256433 1343
rect 256016 1312 256433 1340
rect 256016 1300 256022 1312
rect 256421 1309 256433 1312
rect 256467 1309 256479 1343
rect 256421 1303 256479 1309
rect 256694 1300 256700 1352
rect 256752 1300 256758 1352
rect 256786 1300 256792 1352
rect 256844 1340 256850 1352
rect 257908 1340 257936 1380
rect 256844 1312 257936 1340
rect 256844 1300 256850 1312
rect 257982 1300 257988 1352
rect 258040 1300 258046 1352
rect 258166 1300 258172 1352
rect 258224 1300 258230 1352
rect 258276 1340 258304 1380
rect 258350 1368 258356 1420
rect 258408 1408 258414 1420
rect 260285 1411 260343 1417
rect 260285 1408 260297 1411
rect 258408 1380 260297 1408
rect 258408 1368 258414 1380
rect 260285 1377 260297 1380
rect 260331 1377 260343 1411
rect 260285 1371 260343 1377
rect 261573 1411 261631 1417
rect 261573 1377 261585 1411
rect 261619 1408 261631 1411
rect 261846 1408 261852 1420
rect 261619 1380 261852 1408
rect 261619 1377 261631 1380
rect 261573 1371 261631 1377
rect 261846 1368 261852 1380
rect 261904 1368 261910 1420
rect 269301 1411 269359 1417
rect 269301 1377 269313 1411
rect 269347 1408 269359 1411
rect 271046 1408 271052 1420
rect 269347 1380 271052 1408
rect 269347 1377 269359 1380
rect 269301 1371 269359 1377
rect 271046 1368 271052 1380
rect 271104 1368 271110 1420
rect 258997 1343 259055 1349
rect 258997 1340 259009 1343
rect 258276 1312 259009 1340
rect 258997 1309 259009 1312
rect 259043 1309 259055 1343
rect 258997 1303 259055 1309
rect 259270 1300 259276 1352
rect 259328 1300 259334 1352
rect 260469 1343 260527 1349
rect 260469 1309 260481 1343
rect 260515 1309 260527 1343
rect 260469 1303 260527 1309
rect 250625 1275 250683 1281
rect 250625 1241 250637 1275
rect 250671 1272 250683 1275
rect 255314 1272 255320 1284
rect 250671 1244 255320 1272
rect 250671 1241 250683 1244
rect 250625 1235 250683 1241
rect 255314 1232 255320 1244
rect 255372 1232 255378 1284
rect 255866 1232 255872 1284
rect 255924 1272 255930 1284
rect 258353 1275 258411 1281
rect 258353 1272 258365 1275
rect 255924 1244 258365 1272
rect 255924 1232 255930 1244
rect 258353 1241 258365 1244
rect 258399 1241 258411 1275
rect 258353 1235 258411 1241
rect 260484 1272 260512 1303
rect 260650 1300 260656 1352
rect 260708 1300 260714 1352
rect 261757 1343 261815 1349
rect 261757 1309 261769 1343
rect 261803 1309 261815 1343
rect 261757 1303 261815 1309
rect 261941 1343 261999 1349
rect 261941 1309 261953 1343
rect 261987 1340 261999 1343
rect 262401 1343 262459 1349
rect 262401 1340 262413 1343
rect 261987 1312 262413 1340
rect 261987 1309 261999 1312
rect 261941 1303 261999 1309
rect 262401 1309 262413 1312
rect 262447 1309 262459 1343
rect 262401 1303 262459 1309
rect 261478 1272 261484 1284
rect 260484 1244 261484 1272
rect 248472 1176 250208 1204
rect 248472 1164 248478 1176
rect 251174 1164 251180 1216
rect 251232 1204 251238 1216
rect 252557 1207 252615 1213
rect 252557 1204 252569 1207
rect 251232 1176 252569 1204
rect 251232 1164 251238 1176
rect 252557 1173 252569 1176
rect 252603 1173 252615 1207
rect 252557 1167 252615 1173
rect 255777 1207 255835 1213
rect 255777 1173 255789 1207
rect 255823 1204 255835 1207
rect 258074 1204 258080 1216
rect 255823 1176 258080 1204
rect 255823 1173 255835 1176
rect 255777 1167 255835 1173
rect 258074 1164 258080 1176
rect 258132 1164 258138 1216
rect 258166 1164 258172 1216
rect 258224 1204 258230 1216
rect 260484 1204 260512 1244
rect 261478 1232 261484 1244
rect 261536 1272 261542 1284
rect 261772 1272 261800 1303
rect 263134 1300 263140 1352
rect 263192 1300 263198 1352
rect 264146 1300 264152 1352
rect 264204 1300 264210 1352
rect 264882 1300 264888 1352
rect 264940 1300 264946 1352
rect 265618 1300 265624 1352
rect 265676 1300 265682 1352
rect 266722 1300 266728 1352
rect 266780 1300 266786 1352
rect 267461 1343 267519 1349
rect 267461 1309 267473 1343
rect 267507 1340 267519 1343
rect 267826 1340 267832 1352
rect 267507 1312 267832 1340
rect 267507 1309 267519 1312
rect 267461 1303 267519 1309
rect 267826 1300 267832 1312
rect 267884 1300 267890 1352
rect 268194 1300 268200 1352
rect 268252 1300 268258 1352
rect 269114 1300 269120 1352
rect 269172 1340 269178 1352
rect 269485 1343 269543 1349
rect 269485 1340 269497 1343
rect 269172 1312 269497 1340
rect 269172 1300 269178 1312
rect 269485 1309 269497 1312
rect 269531 1309 269543 1343
rect 269485 1303 269543 1309
rect 269669 1343 269727 1349
rect 269669 1309 269681 1343
rect 269715 1340 269727 1343
rect 270034 1340 270040 1352
rect 269715 1312 270040 1340
rect 269715 1309 269727 1312
rect 269669 1303 269727 1309
rect 270034 1300 270040 1312
rect 270092 1300 270098 1352
rect 270126 1300 270132 1352
rect 270184 1300 270190 1352
rect 261536 1244 261800 1272
rect 261536 1232 261542 1244
rect 258224 1176 260512 1204
rect 258224 1164 258230 1176
rect 261110 1164 261116 1216
rect 261168 1204 261174 1216
rect 262585 1207 262643 1213
rect 262585 1204 262597 1207
rect 261168 1176 262597 1204
rect 261168 1164 261174 1176
rect 262585 1173 262597 1176
rect 262631 1173 262643 1207
rect 262585 1167 262643 1173
rect 262858 1164 262864 1216
rect 262916 1204 262922 1216
rect 263321 1207 263379 1213
rect 263321 1204 263333 1207
rect 262916 1176 263333 1204
rect 262916 1164 262922 1176
rect 263321 1173 263333 1176
rect 263367 1173 263379 1207
rect 263321 1167 263379 1173
rect 264330 1164 264336 1216
rect 264388 1164 264394 1216
rect 264974 1164 264980 1216
rect 265032 1204 265038 1216
rect 265069 1207 265127 1213
rect 265069 1204 265081 1207
rect 265032 1176 265081 1204
rect 265032 1164 265038 1176
rect 265069 1173 265081 1176
rect 265115 1173 265127 1207
rect 265069 1167 265127 1173
rect 265802 1164 265808 1216
rect 265860 1164 265866 1216
rect 266354 1164 266360 1216
rect 266412 1204 266418 1216
rect 266909 1207 266967 1213
rect 266909 1204 266921 1207
rect 266412 1176 266921 1204
rect 266412 1164 266418 1176
rect 266909 1173 266921 1176
rect 266955 1173 266967 1207
rect 266909 1167 266967 1173
rect 267642 1164 267648 1216
rect 267700 1164 267706 1216
rect 268378 1164 268384 1216
rect 268436 1164 268442 1216
rect 270310 1164 270316 1216
rect 270368 1164 270374 1216
rect 1104 1114 271651 1136
rect 1104 1062 68546 1114
rect 68598 1062 68610 1114
rect 68662 1062 68674 1114
rect 68726 1062 68738 1114
rect 68790 1062 68802 1114
rect 68854 1062 136143 1114
rect 136195 1062 136207 1114
rect 136259 1062 136271 1114
rect 136323 1062 136335 1114
rect 136387 1062 136399 1114
rect 136451 1062 203740 1114
rect 203792 1062 203804 1114
rect 203856 1062 203868 1114
rect 203920 1062 203932 1114
rect 203984 1062 203996 1114
rect 204048 1062 271337 1114
rect 271389 1062 271401 1114
rect 271453 1062 271465 1114
rect 271517 1062 271529 1114
rect 271581 1062 271593 1114
rect 271645 1062 271651 1114
rect 1104 1040 271651 1062
rect 2038 960 2044 1012
rect 2096 1000 2102 1012
rect 35986 1000 35992 1012
rect 2096 972 35992 1000
rect 2096 960 2102 972
rect 35986 960 35992 972
rect 36044 960 36050 1012
rect 77478 960 77484 1012
rect 77536 1000 77542 1012
rect 103790 1000 103796 1012
rect 77536 972 103796 1000
rect 77536 960 77542 972
rect 103790 960 103796 972
rect 103848 960 103854 1012
rect 103974 960 103980 1012
rect 104032 1000 104038 1012
rect 108942 1000 108948 1012
rect 104032 972 108948 1000
rect 104032 960 104038 972
rect 108942 960 108948 972
rect 109000 960 109006 1012
rect 110690 1000 110696 1012
rect 109052 972 110696 1000
rect 17310 892 17316 944
rect 17368 932 17374 944
rect 51718 932 51724 944
rect 17368 904 51724 932
rect 17368 892 17374 904
rect 51718 892 51724 904
rect 51776 892 51782 944
rect 74994 892 75000 944
rect 75052 932 75058 944
rect 99834 932 99840 944
rect 75052 904 99840 932
rect 75052 892 75058 904
rect 99834 892 99840 904
rect 99892 892 99898 944
rect 100846 892 100852 944
rect 100904 932 100910 944
rect 100904 904 103468 932
rect 100904 892 100910 904
rect 10594 824 10600 876
rect 10652 864 10658 876
rect 44358 864 44364 876
rect 10652 836 44364 864
rect 10652 824 10658 836
rect 44358 824 44364 836
rect 44416 824 44422 876
rect 77570 824 77576 876
rect 77628 864 77634 876
rect 77628 836 80054 864
rect 77628 824 77634 836
rect 14274 756 14280 808
rect 14332 796 14338 808
rect 45554 796 45560 808
rect 14332 768 45560 796
rect 14332 756 14338 768
rect 45554 756 45560 768
rect 45612 756 45618 808
rect 80026 796 80054 836
rect 92566 824 92572 876
rect 92624 864 92630 876
rect 94774 864 94780 876
rect 92624 836 94780 864
rect 92624 824 92630 836
rect 94774 824 94780 836
rect 94832 824 94838 876
rect 97810 824 97816 876
rect 97868 864 97874 876
rect 103330 864 103336 876
rect 97868 836 103336 864
rect 97868 824 97874 836
rect 103330 824 103336 836
rect 103388 824 103394 876
rect 103440 864 103468 904
rect 103514 892 103520 944
rect 103572 932 103578 944
rect 104618 932 104624 944
rect 103572 904 104624 932
rect 103572 892 103578 904
rect 104618 892 104624 904
rect 104676 892 104682 944
rect 105630 932 105636 944
rect 104728 904 105636 932
rect 104728 864 104756 904
rect 105630 892 105636 904
rect 105688 892 105694 944
rect 108298 892 108304 944
rect 108356 932 108362 944
rect 109052 932 109080 972
rect 110690 960 110696 972
rect 110748 960 110754 1012
rect 110782 960 110788 1012
rect 110840 1000 110846 1012
rect 118142 1000 118148 1012
rect 110840 972 118148 1000
rect 110840 960 110846 972
rect 118142 960 118148 972
rect 118200 960 118206 1012
rect 120534 1000 120540 1012
rect 118252 972 120540 1000
rect 108356 904 109080 932
rect 108356 892 108362 904
rect 109126 892 109132 944
rect 109184 932 109190 944
rect 109184 904 109816 932
rect 109184 892 109190 904
rect 103440 836 104756 864
rect 105538 824 105544 876
rect 105596 864 105602 876
rect 109678 864 109684 876
rect 105596 836 109684 864
rect 105596 824 105602 836
rect 109678 824 109684 836
rect 109736 824 109742 876
rect 109788 864 109816 904
rect 113266 892 113272 944
rect 113324 932 113330 944
rect 118252 932 118280 972
rect 120534 960 120540 972
rect 120592 960 120598 1012
rect 141694 1000 141700 1012
rect 125566 972 141700 1000
rect 125566 932 125594 972
rect 141694 960 141700 972
rect 141752 960 141758 1012
rect 141786 960 141792 1012
rect 141844 1000 141850 1012
rect 145834 1000 145840 1012
rect 141844 972 145840 1000
rect 141844 960 141850 972
rect 145834 960 145840 972
rect 145892 960 145898 1012
rect 147674 960 147680 1012
rect 147732 1000 147738 1012
rect 152274 1000 152280 1012
rect 147732 972 152280 1000
rect 147732 960 147738 972
rect 152274 960 152280 972
rect 152332 960 152338 1012
rect 154022 960 154028 1012
rect 154080 1000 154086 1012
rect 179414 1000 179420 1012
rect 154080 972 179420 1000
rect 154080 960 154086 972
rect 179414 960 179420 972
rect 179472 960 179478 1012
rect 214926 960 214932 1012
rect 214984 1000 214990 1012
rect 217042 1000 217048 1012
rect 214984 972 217048 1000
rect 214984 960 214990 972
rect 217042 960 217048 972
rect 217100 960 217106 1012
rect 218054 960 218060 1012
rect 218112 1000 218118 1012
rect 223114 1000 223120 1012
rect 218112 972 223120 1000
rect 218112 960 218118 972
rect 223114 960 223120 972
rect 223172 960 223178 1012
rect 223298 960 223304 1012
rect 223356 1000 223362 1012
rect 226242 1000 226248 1012
rect 223356 972 226248 1000
rect 223356 960 223362 972
rect 226242 960 226248 972
rect 226300 960 226306 1012
rect 240042 960 240048 1012
rect 240100 1000 240106 1012
rect 249058 1000 249064 1012
rect 240100 972 249064 1000
rect 240100 960 240106 972
rect 249058 960 249064 972
rect 249116 960 249122 1012
rect 250070 960 250076 1012
rect 250128 1000 250134 1012
rect 252830 1000 252836 1012
rect 250128 972 252836 1000
rect 250128 960 250134 972
rect 252830 960 252836 972
rect 252888 960 252894 1012
rect 252922 960 252928 1012
rect 252980 1000 252986 1012
rect 252980 972 253934 1000
rect 252980 960 252986 972
rect 113324 904 118280 932
rect 120736 904 125594 932
rect 113324 892 113330 904
rect 120736 864 120764 904
rect 138934 892 138940 944
rect 138992 932 138998 944
rect 150250 932 150256 944
rect 138992 904 150256 932
rect 138992 892 138998 904
rect 150250 892 150256 904
rect 150308 892 150314 944
rect 150434 892 150440 944
rect 150492 932 150498 944
rect 154850 932 154856 944
rect 150492 904 154856 932
rect 150492 892 150498 904
rect 154850 892 154856 904
rect 154908 892 154914 944
rect 154942 892 154948 944
rect 155000 932 155006 944
rect 155000 904 157334 932
rect 155000 892 155006 904
rect 109788 836 120764 864
rect 121454 824 121460 876
rect 121512 864 121518 876
rect 148318 864 148324 876
rect 121512 836 135254 864
rect 121512 824 121518 836
rect 95234 796 95240 808
rect 80026 768 95240 796
rect 95234 756 95240 768
rect 95292 756 95298 808
rect 96154 756 96160 808
rect 96212 796 96218 808
rect 98730 796 98736 808
rect 96212 768 98736 796
rect 96212 756 96218 768
rect 98730 756 98736 768
rect 98788 756 98794 808
rect 98822 756 98828 808
rect 98880 796 98886 808
rect 110874 796 110880 808
rect 98880 768 110880 796
rect 98880 756 98886 768
rect 110874 756 110880 768
rect 110932 756 110938 808
rect 18690 688 18696 740
rect 18748 728 18754 740
rect 51442 728 51448 740
rect 18748 700 51448 728
rect 18748 688 18754 700
rect 51442 688 51448 700
rect 51500 688 51506 740
rect 80146 688 80152 740
rect 80204 728 80210 740
rect 109954 728 109960 740
rect 80204 700 109960 728
rect 80204 688 80210 700
rect 109954 688 109960 700
rect 110012 688 110018 740
rect 110690 688 110696 740
rect 110748 728 110754 740
rect 112806 728 112812 740
rect 110748 700 112812 728
rect 110748 688 110754 700
rect 112806 688 112812 700
rect 112864 688 112870 740
rect 135226 728 135254 836
rect 143000 836 148324 864
rect 141694 756 141700 808
rect 141752 796 141758 808
rect 143000 796 143028 836
rect 148318 824 148324 836
rect 148376 824 148382 876
rect 148410 824 148416 876
rect 148468 864 148474 876
rect 154206 864 154212 876
rect 148468 836 154212 864
rect 148468 824 148474 836
rect 154206 824 154212 836
rect 154264 824 154270 876
rect 157306 864 157334 904
rect 214650 892 214656 944
rect 214708 932 214714 944
rect 216122 932 216128 944
rect 214708 904 216128 932
rect 214708 892 214714 904
rect 216122 892 216128 904
rect 216180 892 216186 944
rect 216674 892 216680 944
rect 216732 932 216738 944
rect 219526 932 219532 944
rect 216732 904 219532 932
rect 216732 892 216738 904
rect 219526 892 219532 904
rect 219584 892 219590 944
rect 246390 932 246396 944
rect 224926 904 246396 932
rect 213454 864 213460 876
rect 157306 836 213460 864
rect 213454 824 213460 836
rect 213512 824 213518 876
rect 213546 824 213552 876
rect 213604 864 213610 876
rect 224926 864 224954 904
rect 246390 892 246396 904
rect 246448 892 246454 944
rect 248966 892 248972 944
rect 249024 932 249030 944
rect 251726 932 251732 944
rect 249024 904 251732 932
rect 249024 892 249030 904
rect 251726 892 251732 904
rect 251784 892 251790 944
rect 253906 932 253934 972
rect 260742 960 260748 1012
rect 260800 1000 260806 1012
rect 267918 1000 267924 1012
rect 260800 972 267924 1000
rect 260800 960 260806 972
rect 267918 960 267924 972
rect 267976 960 267982 1012
rect 268010 932 268016 944
rect 253906 904 268016 932
rect 268010 892 268016 904
rect 268068 892 268074 944
rect 248782 864 248788 876
rect 213604 836 224954 864
rect 238726 836 248788 864
rect 213604 824 213610 836
rect 141752 768 143028 796
rect 141752 756 141758 768
rect 143994 756 144000 808
rect 144052 796 144058 808
rect 150986 796 150992 808
rect 144052 768 150992 796
rect 144052 756 144058 768
rect 150986 756 150992 768
rect 151044 756 151050 808
rect 151170 756 151176 808
rect 151228 796 151234 808
rect 154666 796 154672 808
rect 151228 768 154672 796
rect 151228 756 151234 768
rect 154666 756 154672 768
rect 154724 756 154730 808
rect 162946 756 162952 808
rect 163004 796 163010 808
rect 163004 768 209774 796
rect 163004 756 163010 768
rect 135226 700 147812 728
rect 7006 620 7012 672
rect 7064 660 7070 672
rect 41322 660 41328 672
rect 7064 632 41328 660
rect 7064 620 7070 632
rect 41322 620 41328 632
rect 41380 620 41386 672
rect 72786 620 72792 672
rect 72844 660 72850 672
rect 92934 660 92940 672
rect 72844 632 92940 660
rect 72844 620 72850 632
rect 92934 620 92940 632
rect 92992 620 92998 672
rect 94866 620 94872 672
rect 94924 660 94930 672
rect 107194 660 107200 672
rect 94924 632 107200 660
rect 94924 620 94930 632
rect 107194 620 107200 632
rect 107252 620 107258 672
rect 108114 620 108120 672
rect 108172 660 108178 672
rect 112622 660 112628 672
rect 108172 632 112628 660
rect 108172 620 108178 632
rect 112622 620 112628 632
rect 112680 620 112686 672
rect 113358 620 113364 672
rect 113416 660 113422 672
rect 113416 632 138014 660
rect 113416 620 113422 632
rect 15746 552 15752 604
rect 15804 592 15810 604
rect 51626 592 51632 604
rect 15804 564 51632 592
rect 15804 552 15810 564
rect 51626 552 51632 564
rect 51684 552 51690 604
rect 82722 552 82728 604
rect 82780 592 82786 604
rect 115198 592 115204 604
rect 82780 564 115204 592
rect 82780 552 82786 564
rect 115198 552 115204 564
rect 115256 552 115262 604
rect 13538 484 13544 536
rect 13596 524 13602 536
rect 47854 524 47860 536
rect 13596 496 47860 524
rect 13596 484 13602 496
rect 47854 484 47860 496
rect 47912 484 47918 536
rect 78950 484 78956 536
rect 79008 524 79014 536
rect 107378 524 107384 536
rect 79008 496 107384 524
rect 79008 484 79014 496
rect 107378 484 107384 496
rect 107436 484 107442 536
rect 137986 524 138014 632
rect 144914 620 144920 672
rect 144972 660 144978 672
rect 146202 660 146208 672
rect 144972 632 146208 660
rect 144972 620 144978 632
rect 146202 620 146208 632
rect 146260 620 146266 672
rect 147674 660 147680 672
rect 147646 620 147680 660
rect 147732 620 147738 672
rect 147784 660 147812 700
rect 147858 688 147864 740
rect 147916 728 147922 740
rect 151722 728 151728 740
rect 147916 700 151728 728
rect 147916 688 147922 700
rect 151722 688 151728 700
rect 151780 688 151786 740
rect 156414 728 156420 740
rect 152384 700 156420 728
rect 152384 660 152412 700
rect 156414 688 156420 700
rect 156472 688 156478 740
rect 160186 688 160192 740
rect 160244 728 160250 740
rect 208578 728 208584 740
rect 160244 700 208584 728
rect 160244 688 160250 700
rect 208578 688 208584 700
rect 208636 688 208642 740
rect 209746 728 209774 768
rect 213638 756 213644 808
rect 213696 796 213702 808
rect 218698 796 218704 808
rect 213696 768 218704 796
rect 213696 756 213702 768
rect 218698 756 218704 768
rect 218756 756 218762 808
rect 220814 756 220820 808
rect 220872 796 220878 808
rect 226426 796 226432 808
rect 220872 768 226432 796
rect 220872 756 220878 768
rect 226426 756 226432 768
rect 226484 756 226490 808
rect 228082 756 228088 808
rect 228140 796 228146 808
rect 238726 796 238754 836
rect 248782 824 248788 836
rect 248840 824 248846 876
rect 259270 864 259276 876
rect 248892 836 259276 864
rect 248892 796 248920 836
rect 259270 824 259276 836
rect 259328 824 259334 876
rect 228140 768 238754 796
rect 244246 768 248920 796
rect 249076 768 253934 796
rect 228140 756 228146 768
rect 215938 728 215944 740
rect 209746 700 215944 728
rect 215938 688 215944 700
rect 215996 688 216002 740
rect 216122 688 216128 740
rect 216180 728 216186 740
rect 226886 728 226892 740
rect 216180 700 226892 728
rect 216180 688 216186 700
rect 226886 688 226892 700
rect 226944 688 226950 740
rect 243354 688 243360 740
rect 243412 728 243418 740
rect 244246 728 244274 768
rect 249076 728 249104 768
rect 243412 700 244274 728
rect 248984 700 249104 728
rect 253906 728 253934 768
rect 255314 756 255320 808
rect 255372 796 255378 808
rect 272058 796 272064 808
rect 255372 768 272064 796
rect 255372 756 255378 768
rect 272058 756 272064 768
rect 272116 756 272122 808
rect 258258 728 258264 740
rect 253906 700 258264 728
rect 243412 688 243418 700
rect 147784 632 152412 660
rect 152458 620 152464 672
rect 152516 660 152522 672
rect 152516 632 157334 660
rect 152516 620 152522 632
rect 144086 552 144092 604
rect 144144 592 144150 604
rect 147646 592 147674 620
rect 153562 592 153568 604
rect 144144 564 147674 592
rect 147876 564 153568 592
rect 144144 552 144150 564
rect 147582 524 147588 536
rect 137986 496 147588 524
rect 147582 484 147588 496
rect 147640 484 147646 536
rect 2866 416 2872 468
rect 2924 456 2930 468
rect 37366 456 37372 468
rect 2924 428 37372 456
rect 2924 416 2930 428
rect 37366 416 37372 428
rect 37424 416 37430 468
rect 74074 416 74080 468
rect 74132 456 74138 468
rect 97074 456 97080 468
rect 74132 428 97080 456
rect 74132 416 74138 428
rect 97074 416 97080 428
rect 97132 416 97138 468
rect 105722 416 105728 468
rect 105780 456 105786 468
rect 110966 456 110972 468
rect 105780 428 110972 456
rect 105780 416 105786 428
rect 110966 416 110972 428
rect 111024 416 111030 468
rect 146938 416 146944 468
rect 146996 456 147002 468
rect 147876 456 147904 564
rect 153562 552 153568 564
rect 153620 552 153626 604
rect 157306 592 157334 632
rect 168374 620 168380 672
rect 168432 660 168438 672
rect 243538 660 243544 672
rect 168432 632 243544 660
rect 168432 620 168438 632
rect 243538 620 243544 632
rect 243596 620 243602 672
rect 243906 620 243912 672
rect 243964 660 243970 672
rect 248984 660 249012 700
rect 258258 688 258264 700
rect 258316 688 258322 740
rect 243964 632 249012 660
rect 243964 620 243970 632
rect 249058 620 249064 672
rect 249116 660 249122 672
rect 260190 660 260196 672
rect 249116 632 260196 660
rect 249116 620 249122 632
rect 260190 620 260196 632
rect 260248 620 260254 672
rect 177022 592 177028 604
rect 157306 564 177028 592
rect 177022 552 177028 564
rect 177080 552 177086 604
rect 208118 552 208124 604
rect 208176 592 208182 604
rect 212626 592 212632 604
rect 208176 564 212632 592
rect 208176 552 208182 564
rect 212626 552 212632 564
rect 212684 552 212690 604
rect 213454 552 213460 604
rect 213512 592 213518 604
rect 216766 592 216772 604
rect 213512 564 216772 592
rect 213512 552 213518 564
rect 216766 552 216772 564
rect 216824 552 216830 604
rect 217686 552 217692 604
rect 217744 592 217750 604
rect 222930 592 222936 604
rect 217744 564 222936 592
rect 217744 552 217750 564
rect 222930 552 222936 564
rect 222988 552 222994 604
rect 223022 552 223028 604
rect 223080 592 223086 604
rect 254118 592 254124 604
rect 223080 564 254124 592
rect 223080 552 223086 564
rect 254118 552 254124 564
rect 254176 552 254182 604
rect 151630 484 151636 536
rect 151688 524 151694 536
rect 153930 524 153936 536
rect 151688 496 153936 524
rect 151688 484 151694 496
rect 153930 484 153936 496
rect 153988 484 153994 536
rect 154298 484 154304 536
rect 154356 524 154362 536
rect 187142 524 187148 536
rect 154356 496 187148 524
rect 154356 484 154362 496
rect 187142 484 187148 496
rect 187200 484 187206 536
rect 209866 484 209872 536
rect 209924 524 209930 536
rect 243814 524 243820 536
rect 209924 496 243820 524
rect 209924 484 209930 496
rect 243814 484 243820 496
rect 243872 484 243878 536
rect 246850 484 246856 536
rect 246908 524 246914 536
rect 256694 524 256700 536
rect 246908 496 256700 524
rect 246908 484 246914 496
rect 256694 484 256700 496
rect 256752 484 256758 536
rect 146996 428 147904 456
rect 146996 416 147002 428
rect 148962 416 148968 468
rect 149020 456 149026 468
rect 172422 456 172428 468
rect 149020 428 172428 456
rect 149020 416 149026 428
rect 172422 416 172428 428
rect 172480 416 172486 468
rect 208670 416 208676 468
rect 208728 456 208734 468
rect 214558 456 214564 468
rect 208728 428 214564 456
rect 208728 416 208734 428
rect 214558 416 214564 428
rect 214616 416 214622 468
rect 216306 416 216312 468
rect 216364 456 216370 468
rect 251542 456 251548 468
rect 216364 428 251548 456
rect 216364 416 216370 428
rect 251542 416 251548 428
rect 251600 416 251606 468
rect 5442 348 5448 400
rect 5500 388 5506 400
rect 40034 388 40040 400
rect 5500 360 40040 388
rect 5500 348 5506 360
rect 40034 348 40040 360
rect 40092 348 40098 400
rect 92290 348 92296 400
rect 92348 388 92354 400
rect 98822 388 98828 400
rect 92348 360 98828 388
rect 92348 348 92354 360
rect 98822 348 98828 360
rect 98880 348 98886 400
rect 145006 348 145012 400
rect 145064 388 145070 400
rect 150802 388 150808 400
rect 145064 360 150808 388
rect 145064 348 145070 360
rect 150802 348 150808 360
rect 150860 348 150866 400
rect 158070 348 158076 400
rect 158128 388 158134 400
rect 172514 388 172520 400
rect 158128 360 172520 388
rect 158128 348 158134 360
rect 172514 348 172520 360
rect 172572 348 172578 400
rect 214466 348 214472 400
rect 214524 388 214530 400
rect 220538 388 220544 400
rect 214524 360 220544 388
rect 214524 348 214530 360
rect 220538 348 220544 360
rect 220596 348 220602 400
rect 222378 348 222384 400
rect 222436 388 222442 400
rect 241054 388 241060 400
rect 222436 360 241060 388
rect 222436 348 222442 360
rect 241054 348 241060 360
rect 241112 348 241118 400
rect 242986 348 242992 400
rect 243044 388 243050 400
rect 256418 388 256424 400
rect 243044 360 256424 388
rect 243044 348 243050 360
rect 256418 348 256424 360
rect 256476 348 256482 400
rect 147674 280 147680 332
rect 147732 320 147738 332
rect 154574 320 154580 332
rect 147732 292 154580 320
rect 147732 280 147738 292
rect 154574 280 154580 292
rect 154632 280 154638 332
rect 154758 280 154764 332
rect 154816 320 154822 332
rect 184566 320 184572 332
rect 154816 292 184572 320
rect 154816 280 154822 292
rect 184566 280 184572 292
rect 184624 280 184630 332
rect 212994 280 213000 332
rect 213052 320 213058 332
rect 218238 320 218244 332
rect 213052 292 218244 320
rect 213052 280 213058 292
rect 218238 280 218244 292
rect 218296 280 218302 332
rect 218790 280 218796 332
rect 218848 320 218854 332
rect 228174 320 228180 332
rect 218848 292 228180 320
rect 218848 280 218854 292
rect 228174 280 228180 292
rect 228232 280 228238 332
rect 230566 280 230572 332
rect 230624 320 230630 332
rect 248046 320 248052 332
rect 230624 292 248052 320
rect 230624 280 230630 292
rect 248046 280 248052 292
rect 248104 280 248110 332
rect 100478 212 100484 264
rect 100536 252 100542 264
rect 144730 252 144736 264
rect 100536 224 144736 252
rect 100536 212 100542 224
rect 144730 212 144736 224
rect 144788 212 144794 264
rect 155310 212 155316 264
rect 155368 252 155374 264
rect 213914 252 213920 264
rect 155368 224 213920 252
rect 155368 212 155374 224
rect 213914 212 213920 224
rect 213972 212 213978 264
rect 218606 212 218612 264
rect 218664 252 218670 264
rect 223022 252 223028 264
rect 218664 224 223028 252
rect 218664 212 218670 224
rect 223022 212 223028 224
rect 223080 212 223086 264
rect 224954 212 224960 264
rect 225012 252 225018 264
rect 244826 252 244832 264
rect 225012 224 244832 252
rect 225012 212 225018 224
rect 244826 212 244832 224
rect 244884 212 244890 264
rect 209498 144 209504 196
rect 209556 184 209562 196
rect 211062 184 211068 196
rect 209556 156 211068 184
rect 209556 144 209562 156
rect 211062 144 211068 156
rect 211120 184 211126 196
rect 243722 184 243728 196
rect 211120 156 243728 184
rect 211120 144 211126 156
rect 243722 144 243728 156
rect 243780 144 243786 196
rect 28810 76 28816 128
rect 28868 116 28874 128
rect 28994 116 29000 128
rect 28868 88 29000 116
rect 28868 76 28874 88
rect 28994 76 29000 88
rect 29052 76 29058 128
rect 149330 8 149336 60
rect 149388 48 149394 60
rect 181990 48 181996 60
rect 149388 20 181996 48
rect 149388 8 149394 20
rect 181990 8 181996 20
rect 182048 8 182054 60
<< via1 >>
rect 82084 10820 82136 10872
rect 94596 10820 94648 10872
rect 94780 10820 94832 10872
rect 100760 10820 100812 10872
rect 158536 10820 158588 10872
rect 166448 10820 166500 10872
rect 69848 10752 69900 10804
rect 81532 10752 81584 10804
rect 81716 10752 81768 10804
rect 93952 10752 94004 10804
rect 99196 10752 99248 10804
rect 132776 10752 132828 10804
rect 133788 10752 133840 10804
rect 146576 10752 146628 10804
rect 177580 10752 177632 10804
rect 92388 10684 92440 10736
rect 125876 10684 125928 10736
rect 151728 10684 151780 10736
rect 162768 10684 162820 10736
rect 165068 10684 165120 10736
rect 217876 10684 217928 10736
rect 60648 10616 60700 10668
rect 82084 10616 82136 10668
rect 94964 10616 95016 10668
rect 106188 10616 106240 10668
rect 21640 10412 21692 10464
rect 30656 10412 30708 10464
rect 27712 10344 27764 10396
rect 62028 10412 62080 10464
rect 96436 10548 96488 10600
rect 98644 10548 98696 10600
rect 100024 10548 100076 10600
rect 127624 10616 127676 10668
rect 131120 10616 131172 10668
rect 131856 10616 131908 10668
rect 158536 10616 158588 10668
rect 158628 10616 158680 10668
rect 164516 10616 164568 10668
rect 202328 10616 202380 10668
rect 220176 10820 220228 10872
rect 224960 10820 225012 10872
rect 219900 10752 219952 10804
rect 230664 10820 230716 10872
rect 225144 10752 225196 10804
rect 233608 10752 233660 10804
rect 257620 10820 257672 10872
rect 266912 10820 266964 10872
rect 264704 10752 264756 10804
rect 234712 10684 234764 10736
rect 236644 10684 236696 10736
rect 263784 10684 263836 10736
rect 218796 10616 218848 10668
rect 226708 10616 226760 10668
rect 226984 10616 227036 10668
rect 229100 10616 229152 10668
rect 258540 10616 258592 10668
rect 267556 10616 267608 10668
rect 148692 10548 148744 10600
rect 180708 10548 180760 10600
rect 200120 10548 200172 10600
rect 228640 10548 228692 10600
rect 91008 10480 91060 10532
rect 124220 10480 124272 10532
rect 124680 10480 124732 10532
rect 158812 10480 158864 10532
rect 160468 10480 160520 10532
rect 182088 10480 182140 10532
rect 193312 10480 193364 10532
rect 220084 10480 220136 10532
rect 223488 10480 223540 10532
rect 264428 10548 264480 10600
rect 228824 10480 228876 10532
rect 232780 10480 232832 10532
rect 233608 10480 233660 10532
rect 257620 10480 257672 10532
rect 258632 10480 258684 10532
rect 267004 10480 267056 10532
rect 74540 10412 74592 10464
rect 96620 10412 96672 10464
rect 98828 10412 98880 10464
rect 122840 10412 122892 10464
rect 145380 10412 145432 10464
rect 178040 10412 178092 10464
rect 223580 10412 223632 10464
rect 251272 10412 251324 10464
rect 259552 10412 259604 10464
rect 269028 10412 269080 10464
rect 24492 10276 24544 10328
rect 58532 10276 58584 10328
rect 29552 10208 29604 10260
rect 63224 10276 63276 10328
rect 80612 10344 80664 10396
rect 90732 10344 90784 10396
rect 91008 10344 91060 10396
rect 93308 10344 93360 10396
rect 105452 10344 105504 10396
rect 126704 10344 126756 10396
rect 161112 10344 161164 10396
rect 162124 10344 162176 10396
rect 216588 10344 216640 10396
rect 219072 10344 219124 10396
rect 244096 10344 244148 10396
rect 260196 10344 260248 10396
rect 268292 10344 268344 10396
rect 92848 10276 92900 10328
rect 92940 10276 92992 10328
rect 95516 10276 95568 10328
rect 95608 10276 95660 10328
rect 107016 10276 107068 10328
rect 140228 10276 140280 10328
rect 174268 10276 174320 10328
rect 196164 10276 196216 10328
rect 226984 10276 227036 10328
rect 227076 10276 227128 10328
rect 231860 10276 231912 10328
rect 231952 10276 232004 10328
rect 239312 10276 239364 10328
rect 96528 10208 96580 10260
rect 131120 10208 131172 10260
rect 133788 10208 133840 10260
rect 166724 10208 166776 10260
rect 203064 10208 203116 10260
rect 236000 10208 236052 10260
rect 268108 10276 268160 10328
rect 259644 10208 259696 10260
rect 267096 10208 267148 10260
rect 5908 10140 5960 10192
rect 39580 10140 39632 10192
rect 56324 10140 56376 10192
rect 80612 10140 80664 10192
rect 81072 10140 81124 10192
rect 92940 10140 92992 10192
rect 93032 10140 93084 10192
rect 126704 10140 126756 10192
rect 141424 10140 141476 10192
rect 175556 10140 175608 10192
rect 197084 10140 197136 10192
rect 204352 10140 204404 10192
rect 211252 10140 211304 10192
rect 227076 10140 227128 10192
rect 227168 10140 227220 10192
rect 22652 10072 22704 10124
rect 56876 10072 56928 10124
rect 22468 10004 22520 10056
rect 30564 10004 30616 10056
rect 30656 10004 30708 10056
rect 56416 10004 56468 10056
rect 91008 10072 91060 10124
rect 124680 10072 124732 10124
rect 125876 10072 125928 10124
rect 61476 10004 61528 10056
rect 95424 10004 95476 10056
rect 95516 10004 95568 10056
rect 95792 10004 95844 10056
rect 98552 10004 98604 10056
rect 98644 10004 98696 10056
rect 130108 10004 130160 10056
rect 25504 9936 25556 9988
rect 59728 9936 59780 9988
rect 81532 9936 81584 9988
rect 110512 9936 110564 9988
rect 142436 10072 142488 10124
rect 152556 10072 152608 10124
rect 159640 10072 159692 10124
rect 229008 10072 229060 10124
rect 159916 10004 159968 10056
rect 18052 9868 18104 9920
rect 27620 9868 27672 9920
rect 30104 9868 30156 9920
rect 64052 9868 64104 9920
rect 84016 9868 84068 9920
rect 117044 9868 117096 9920
rect 121644 9868 121696 9920
rect 130200 9868 130252 9920
rect 152464 9936 152516 9988
rect 161940 9936 161992 9988
rect 158628 9868 158680 9920
rect 158720 9868 158772 9920
rect 165344 10004 165396 10056
rect 166172 10004 166224 10056
rect 219992 10004 220044 10056
rect 220452 10004 220504 10056
rect 228732 10004 228784 10056
rect 231860 10140 231912 10192
rect 265624 10140 265676 10192
rect 229192 10072 229244 10124
rect 231952 10072 232004 10124
rect 233516 10072 233568 10124
rect 258540 10072 258592 10124
rect 258908 10072 258960 10124
rect 266544 10072 266596 10124
rect 261576 10004 261628 10056
rect 262680 10004 262732 10056
rect 268384 10004 268436 10056
rect 163872 9936 163924 9988
rect 216588 9936 216640 9988
rect 220084 9936 220136 9988
rect 227168 9936 227220 9988
rect 227812 9936 227864 9988
rect 262128 9936 262180 9988
rect 264796 9936 264848 9988
rect 268200 9936 268252 9988
rect 164240 9868 164292 9920
rect 176844 9868 176896 9920
rect 196348 9868 196400 9920
rect 204260 9868 204312 9920
rect 204352 9868 204404 9920
rect 220176 9868 220228 9920
rect 220268 9868 220320 9920
rect 229652 9868 229704 9920
rect 230940 9868 230992 9920
rect 231032 9868 231084 9920
rect 236644 9868 236696 9920
rect 236736 9868 236788 9920
rect 258724 9868 258776 9920
rect 258816 9868 258868 9920
rect 264244 9868 264296 9920
rect 265440 9868 265492 9920
rect 267740 9868 267792 9920
rect 68546 9766 68598 9818
rect 68610 9766 68662 9818
rect 68674 9766 68726 9818
rect 68738 9766 68790 9818
rect 68802 9766 68854 9818
rect 136143 9766 136195 9818
rect 136207 9766 136259 9818
rect 136271 9766 136323 9818
rect 136335 9766 136387 9818
rect 136399 9766 136451 9818
rect 203740 9766 203792 9818
rect 203804 9766 203856 9818
rect 203868 9766 203920 9818
rect 203932 9766 203984 9818
rect 203996 9766 204048 9818
rect 271337 9766 271389 9818
rect 271401 9766 271453 9818
rect 271465 9766 271517 9818
rect 271529 9766 271581 9818
rect 271593 9766 271645 9818
rect 5908 9707 5960 9716
rect 5908 9673 5917 9707
rect 5917 9673 5951 9707
rect 5951 9673 5960 9707
rect 5908 9664 5960 9673
rect 1676 9639 1728 9648
rect 1676 9605 1685 9639
rect 1685 9605 1719 9639
rect 1719 9605 1728 9639
rect 1676 9596 1728 9605
rect 2412 9639 2464 9648
rect 2412 9605 2421 9639
rect 2421 9605 2455 9639
rect 2455 9605 2464 9639
rect 2412 9596 2464 9605
rect 3240 9639 3292 9648
rect 3240 9605 3249 9639
rect 3249 9605 3283 9639
rect 3283 9605 3292 9639
rect 3240 9596 3292 9605
rect 4344 9639 4396 9648
rect 4344 9605 4353 9639
rect 4353 9605 4387 9639
rect 4387 9605 4396 9639
rect 4344 9596 4396 9605
rect 5080 9639 5132 9648
rect 5080 9605 5089 9639
rect 5089 9605 5123 9639
rect 5123 9605 5132 9639
rect 5080 9596 5132 9605
rect 5816 9639 5868 9648
rect 5816 9605 5825 9639
rect 5825 9605 5859 9639
rect 5859 9605 5868 9639
rect 5816 9596 5868 9605
rect 6828 9639 6880 9648
rect 6828 9605 6837 9639
rect 6837 9605 6871 9639
rect 6871 9605 6880 9639
rect 6828 9596 6880 9605
rect 7564 9639 7616 9648
rect 7564 9605 7573 9639
rect 7573 9605 7607 9639
rect 7607 9605 7616 9639
rect 7564 9596 7616 9605
rect 8392 9639 8444 9648
rect 8392 9605 8401 9639
rect 8401 9605 8435 9639
rect 8435 9605 8444 9639
rect 8392 9596 8444 9605
rect 9588 9596 9640 9648
rect 10232 9639 10284 9648
rect 10232 9605 10241 9639
rect 10241 9605 10275 9639
rect 10275 9605 10284 9639
rect 10232 9596 10284 9605
rect 10968 9639 11020 9648
rect 10968 9605 10977 9639
rect 10977 9605 11011 9639
rect 11011 9605 11020 9639
rect 10968 9596 11020 9605
rect 11980 9639 12032 9648
rect 11980 9605 11989 9639
rect 11989 9605 12023 9639
rect 12023 9605 12032 9639
rect 11980 9596 12032 9605
rect 12716 9639 12768 9648
rect 12716 9605 12725 9639
rect 12725 9605 12759 9639
rect 12759 9605 12768 9639
rect 12716 9596 12768 9605
rect 13728 9596 13780 9648
rect 14648 9639 14700 9648
rect 14648 9605 14657 9639
rect 14657 9605 14691 9639
rect 14691 9605 14700 9639
rect 14648 9596 14700 9605
rect 15384 9639 15436 9648
rect 15384 9605 15393 9639
rect 15393 9605 15427 9639
rect 15427 9605 15436 9639
rect 15384 9596 15436 9605
rect 16120 9639 16172 9648
rect 16120 9605 16129 9639
rect 16129 9605 16163 9639
rect 16163 9605 16172 9639
rect 16120 9596 16172 9605
rect 17132 9639 17184 9648
rect 17132 9605 17141 9639
rect 17141 9605 17175 9639
rect 17175 9605 17184 9639
rect 17132 9596 17184 9605
rect 17868 9639 17920 9648
rect 17868 9605 17877 9639
rect 17877 9605 17911 9639
rect 17911 9605 17920 9639
rect 17868 9596 17920 9605
rect 18052 9639 18104 9648
rect 18052 9605 18061 9639
rect 18061 9605 18095 9639
rect 18095 9605 18104 9639
rect 18052 9596 18104 9605
rect 18604 9639 18656 9648
rect 18604 9605 18613 9639
rect 18613 9605 18647 9639
rect 18647 9605 18656 9639
rect 18604 9596 18656 9605
rect 24400 9596 24452 9648
rect 22468 9571 22520 9580
rect 22468 9537 22477 9571
rect 22477 9537 22511 9571
rect 22511 9537 22520 9571
rect 22468 9528 22520 9537
rect 25688 9571 25740 9580
rect 25688 9537 25697 9571
rect 25697 9537 25731 9571
rect 25731 9537 25740 9571
rect 25688 9528 25740 9537
rect 16488 9460 16540 9512
rect 17224 9460 17276 9512
rect 7564 9392 7616 9444
rect 9680 9435 9732 9444
rect 9680 9401 9689 9435
rect 9689 9401 9723 9435
rect 9723 9401 9732 9435
rect 9680 9392 9732 9401
rect 12900 9435 12952 9444
rect 12900 9401 12909 9435
rect 12909 9401 12943 9435
rect 12943 9401 12952 9435
rect 12900 9392 12952 9401
rect 13728 9435 13780 9444
rect 13728 9401 13737 9435
rect 13737 9401 13771 9435
rect 13771 9401 13780 9435
rect 13728 9392 13780 9401
rect 15568 9435 15620 9444
rect 15568 9401 15577 9435
rect 15577 9401 15611 9435
rect 15611 9401 15620 9435
rect 15568 9392 15620 9401
rect 19156 9392 19208 9444
rect 23756 9460 23808 9512
rect 24308 9460 24360 9512
rect 25504 9503 25556 9512
rect 24584 9392 24636 9444
rect 25504 9469 25513 9503
rect 25513 9469 25547 9503
rect 25547 9469 25556 9503
rect 25504 9460 25556 9469
rect 25872 9664 25924 9716
rect 27344 9707 27396 9716
rect 27344 9673 27353 9707
rect 27353 9673 27387 9707
rect 27387 9673 27396 9707
rect 27344 9664 27396 9673
rect 29092 9707 29144 9716
rect 29092 9673 29101 9707
rect 29101 9673 29135 9707
rect 29135 9673 29144 9707
rect 29092 9664 29144 9673
rect 30288 9664 30340 9716
rect 32496 9707 32548 9716
rect 32496 9673 32505 9707
rect 32505 9673 32539 9707
rect 32539 9673 32548 9707
rect 32496 9664 32548 9673
rect 38200 9664 38252 9716
rect 39672 9664 39724 9716
rect 54760 9664 54812 9716
rect 54852 9664 54904 9716
rect 56508 9707 56560 9716
rect 56508 9673 56517 9707
rect 56517 9673 56551 9707
rect 56551 9673 56560 9707
rect 56508 9664 56560 9673
rect 57336 9707 57388 9716
rect 57336 9673 57345 9707
rect 57345 9673 57379 9707
rect 57379 9673 57388 9707
rect 57336 9664 57388 9673
rect 57796 9664 57848 9716
rect 61752 9707 61804 9716
rect 61752 9673 61761 9707
rect 61761 9673 61795 9707
rect 61795 9673 61804 9707
rect 61752 9664 61804 9673
rect 62488 9707 62540 9716
rect 62488 9673 62497 9707
rect 62497 9673 62531 9707
rect 62531 9673 62540 9707
rect 62488 9664 62540 9673
rect 63408 9707 63460 9716
rect 63408 9673 63417 9707
rect 63417 9673 63451 9707
rect 63451 9673 63460 9707
rect 63408 9664 63460 9673
rect 26148 9596 26200 9648
rect 54300 9596 54352 9648
rect 54576 9596 54628 9648
rect 60648 9596 60700 9648
rect 67364 9596 67416 9648
rect 76380 9596 76432 9648
rect 26516 9528 26568 9580
rect 29828 9528 29880 9580
rect 30380 9528 30432 9580
rect 32128 9528 32180 9580
rect 35624 9571 35676 9580
rect 35624 9537 35633 9571
rect 35633 9537 35667 9571
rect 35667 9537 35676 9571
rect 35624 9528 35676 9537
rect 36268 9571 36320 9580
rect 36268 9537 36277 9571
rect 36277 9537 36311 9571
rect 36311 9537 36320 9571
rect 36268 9528 36320 9537
rect 36912 9571 36964 9580
rect 36912 9537 36921 9571
rect 36921 9537 36955 9571
rect 36955 9537 36964 9571
rect 36912 9528 36964 9537
rect 38108 9571 38160 9580
rect 38108 9537 38117 9571
rect 38117 9537 38151 9571
rect 38151 9537 38160 9571
rect 38108 9528 38160 9537
rect 38844 9571 38896 9580
rect 38844 9537 38853 9571
rect 38853 9537 38887 9571
rect 38887 9537 38896 9571
rect 38844 9528 38896 9537
rect 39488 9571 39540 9580
rect 39488 9537 39497 9571
rect 39497 9537 39531 9571
rect 39531 9537 39540 9571
rect 39488 9528 39540 9537
rect 40776 9571 40828 9580
rect 40776 9537 40785 9571
rect 40785 9537 40819 9571
rect 40819 9537 40828 9571
rect 40776 9528 40828 9537
rect 41420 9571 41472 9580
rect 41420 9537 41429 9571
rect 41429 9537 41463 9571
rect 41463 9537 41472 9571
rect 41420 9528 41472 9537
rect 42064 9571 42116 9580
rect 42064 9537 42073 9571
rect 42073 9537 42107 9571
rect 42107 9537 42116 9571
rect 42064 9528 42116 9537
rect 43260 9571 43312 9580
rect 43260 9537 43269 9571
rect 43269 9537 43303 9571
rect 43303 9537 43312 9571
rect 43260 9528 43312 9537
rect 43996 9571 44048 9580
rect 43996 9537 44005 9571
rect 44005 9537 44039 9571
rect 44039 9537 44048 9571
rect 43996 9528 44048 9537
rect 44640 9571 44692 9580
rect 44640 9537 44649 9571
rect 44649 9537 44683 9571
rect 44683 9537 44692 9571
rect 44640 9528 44692 9537
rect 45928 9571 45980 9580
rect 45928 9537 45937 9571
rect 45937 9537 45971 9571
rect 45971 9537 45980 9571
rect 45928 9528 45980 9537
rect 46572 9571 46624 9580
rect 46572 9537 46581 9571
rect 46581 9537 46615 9571
rect 46615 9537 46624 9571
rect 46572 9528 46624 9537
rect 47216 9571 47268 9580
rect 47216 9537 47225 9571
rect 47225 9537 47259 9571
rect 47259 9537 47268 9571
rect 47216 9528 47268 9537
rect 48228 9528 48280 9580
rect 49148 9571 49200 9580
rect 49148 9537 49157 9571
rect 49157 9537 49191 9571
rect 49191 9537 49200 9571
rect 49148 9528 49200 9537
rect 49792 9571 49844 9580
rect 49792 9537 49801 9571
rect 49801 9537 49835 9571
rect 49835 9537 49844 9571
rect 49792 9528 49844 9537
rect 50620 9571 50672 9580
rect 50620 9537 50629 9571
rect 50629 9537 50663 9571
rect 50663 9537 50672 9571
rect 50620 9528 50672 9537
rect 51356 9571 51408 9580
rect 51356 9537 51365 9571
rect 51365 9537 51399 9571
rect 51399 9537 51408 9571
rect 51356 9528 51408 9537
rect 52092 9571 52144 9580
rect 52092 9537 52101 9571
rect 52101 9537 52135 9571
rect 52135 9537 52144 9571
rect 52092 9528 52144 9537
rect 53104 9571 53156 9580
rect 53104 9537 53113 9571
rect 53113 9537 53147 9571
rect 53147 9537 53156 9571
rect 53104 9528 53156 9537
rect 54668 9528 54720 9580
rect 54944 9528 54996 9580
rect 56600 9528 56652 9580
rect 57336 9528 57388 9580
rect 58072 9571 58124 9580
rect 58072 9537 58081 9571
rect 58081 9537 58115 9571
rect 58115 9537 58124 9571
rect 58072 9528 58124 9537
rect 62212 9528 62264 9580
rect 62580 9528 62632 9580
rect 62764 9528 62816 9580
rect 69112 9571 69164 9580
rect 69112 9537 69121 9571
rect 69121 9537 69155 9571
rect 69155 9537 69164 9571
rect 69112 9528 69164 9537
rect 70308 9528 70360 9580
rect 71504 9571 71556 9580
rect 71504 9537 71513 9571
rect 71513 9537 71547 9571
rect 71547 9537 71556 9571
rect 71504 9528 71556 9537
rect 72148 9571 72200 9580
rect 72148 9537 72157 9571
rect 72157 9537 72191 9571
rect 72191 9537 72200 9571
rect 72148 9528 72200 9537
rect 74724 9571 74776 9580
rect 74724 9537 74733 9571
rect 74733 9537 74767 9571
rect 74767 9537 74776 9571
rect 74724 9528 74776 9537
rect 77300 9571 77352 9580
rect 77300 9537 77309 9571
rect 77309 9537 77343 9571
rect 77343 9537 77352 9571
rect 77300 9528 77352 9537
rect 30472 9460 30524 9512
rect 30564 9460 30616 9512
rect 25228 9392 25280 9444
rect 46204 9392 46256 9444
rect 48596 9392 48648 9444
rect 51816 9392 51868 9444
rect 54300 9503 54352 9512
rect 54300 9469 54309 9503
rect 54309 9469 54343 9503
rect 54343 9469 54352 9503
rect 54300 9460 54352 9469
rect 54760 9460 54812 9512
rect 66076 9460 66128 9512
rect 69848 9503 69900 9512
rect 69848 9469 69857 9503
rect 69857 9469 69891 9503
rect 69891 9469 69900 9503
rect 69848 9460 69900 9469
rect 56324 9392 56376 9444
rect 59728 9392 59780 9444
rect 3240 9324 3292 9376
rect 4068 9324 4120 9376
rect 4436 9367 4488 9376
rect 4436 9333 4445 9367
rect 4445 9333 4479 9367
rect 4479 9333 4488 9367
rect 4436 9324 4488 9333
rect 5172 9367 5224 9376
rect 5172 9333 5181 9367
rect 5181 9333 5215 9367
rect 5215 9333 5224 9367
rect 5172 9324 5224 9333
rect 7656 9367 7708 9376
rect 7656 9333 7665 9367
rect 7665 9333 7699 9367
rect 7699 9333 7708 9367
rect 7656 9324 7708 9333
rect 10324 9367 10376 9376
rect 10324 9333 10333 9367
rect 10333 9333 10367 9367
rect 10367 9333 10376 9367
rect 10324 9324 10376 9333
rect 11060 9367 11112 9376
rect 11060 9333 11069 9367
rect 11069 9333 11103 9367
rect 11103 9333 11112 9367
rect 11060 9324 11112 9333
rect 14740 9367 14792 9376
rect 14740 9333 14749 9367
rect 14749 9333 14783 9367
rect 14783 9333 14792 9367
rect 14740 9324 14792 9333
rect 18604 9324 18656 9376
rect 18696 9367 18748 9376
rect 18696 9333 18705 9367
rect 18705 9333 18739 9367
rect 18739 9333 18748 9367
rect 18696 9324 18748 9333
rect 20260 9324 20312 9376
rect 22928 9324 22980 9376
rect 24676 9324 24728 9376
rect 25136 9367 25188 9376
rect 25136 9333 25145 9367
rect 25145 9333 25179 9367
rect 25179 9333 25188 9367
rect 25136 9324 25188 9333
rect 35624 9324 35676 9376
rect 35808 9324 35860 9376
rect 36636 9324 36688 9376
rect 37924 9367 37976 9376
rect 37924 9333 37933 9367
rect 37933 9333 37967 9367
rect 37967 9333 37976 9367
rect 37924 9324 37976 9333
rect 38660 9367 38712 9376
rect 38660 9333 38669 9367
rect 38669 9333 38703 9367
rect 38703 9333 38712 9367
rect 38660 9324 38712 9333
rect 40500 9324 40552 9376
rect 41052 9324 41104 9376
rect 41788 9324 41840 9376
rect 42892 9324 42944 9376
rect 43260 9324 43312 9376
rect 43904 9324 43956 9376
rect 45652 9324 45704 9376
rect 46020 9324 46072 9376
rect 47032 9367 47084 9376
rect 47032 9333 47041 9367
rect 47041 9333 47075 9367
rect 47075 9333 47084 9367
rect 47032 9324 47084 9333
rect 48228 9367 48280 9376
rect 48228 9333 48237 9367
rect 48237 9333 48271 9367
rect 48271 9333 48280 9367
rect 48228 9324 48280 9333
rect 48412 9324 48464 9376
rect 50436 9367 50488 9376
rect 50436 9333 50445 9367
rect 50445 9333 50479 9367
rect 50479 9333 50488 9367
rect 50436 9324 50488 9333
rect 51264 9324 51316 9376
rect 52276 9324 52328 9376
rect 53104 9324 53156 9376
rect 59912 9324 59964 9376
rect 73712 9392 73764 9444
rect 75828 9460 75880 9512
rect 77576 9503 77628 9512
rect 77576 9469 77585 9503
rect 77585 9469 77619 9503
rect 77619 9469 77628 9503
rect 77576 9460 77628 9469
rect 83188 9664 83240 9716
rect 84016 9707 84068 9716
rect 84016 9673 84025 9707
rect 84025 9673 84059 9707
rect 84059 9673 84068 9707
rect 84016 9664 84068 9673
rect 79232 9639 79284 9648
rect 79232 9605 79241 9639
rect 79241 9605 79275 9639
rect 79275 9605 79284 9639
rect 79232 9596 79284 9605
rect 79968 9528 80020 9580
rect 81624 9571 81676 9580
rect 81624 9537 81633 9571
rect 81633 9537 81667 9571
rect 81667 9537 81676 9571
rect 81624 9528 81676 9537
rect 83096 9639 83148 9648
rect 83096 9605 83105 9639
rect 83105 9605 83139 9639
rect 83139 9605 83148 9639
rect 83096 9596 83148 9605
rect 83924 9639 83976 9648
rect 83924 9605 83933 9639
rect 83933 9605 83967 9639
rect 83967 9605 83976 9639
rect 83924 9596 83976 9605
rect 84660 9639 84712 9648
rect 84660 9605 84669 9639
rect 84669 9605 84703 9639
rect 84703 9605 84712 9639
rect 84660 9596 84712 9605
rect 85396 9639 85448 9648
rect 85396 9605 85405 9639
rect 85405 9605 85439 9639
rect 85439 9605 85448 9639
rect 85396 9596 85448 9605
rect 92756 9707 92808 9716
rect 92756 9673 92765 9707
rect 92765 9673 92799 9707
rect 92799 9673 92808 9707
rect 92756 9664 92808 9673
rect 93492 9707 93544 9716
rect 93492 9673 93501 9707
rect 93501 9673 93535 9707
rect 93535 9673 93544 9707
rect 93492 9664 93544 9673
rect 94596 9664 94648 9716
rect 95976 9664 96028 9716
rect 96068 9707 96120 9716
rect 96068 9673 96077 9707
rect 96077 9673 96111 9707
rect 96111 9673 96120 9707
rect 96068 9664 96120 9673
rect 96344 9664 96396 9716
rect 99380 9664 99432 9716
rect 100484 9707 100536 9716
rect 100484 9673 100493 9707
rect 100493 9673 100527 9707
rect 100527 9673 100536 9707
rect 100484 9664 100536 9673
rect 100668 9664 100720 9716
rect 105452 9707 105504 9716
rect 105452 9673 105461 9707
rect 105461 9673 105495 9707
rect 105495 9673 105504 9707
rect 105452 9664 105504 9673
rect 106188 9707 106240 9716
rect 106188 9673 106197 9707
rect 106197 9673 106231 9707
rect 106231 9673 106240 9707
rect 106188 9664 106240 9673
rect 86776 9571 86828 9580
rect 86776 9537 86785 9571
rect 86785 9537 86819 9571
rect 86819 9537 86828 9571
rect 86776 9528 86828 9537
rect 80152 9503 80204 9512
rect 80152 9469 80161 9503
rect 80161 9469 80195 9503
rect 80195 9469 80204 9503
rect 80152 9460 80204 9469
rect 88984 9460 89036 9512
rect 89444 9528 89496 9580
rect 90088 9528 90140 9580
rect 91560 9571 91612 9580
rect 91560 9537 91569 9571
rect 91569 9537 91603 9571
rect 91603 9537 91612 9571
rect 91560 9528 91612 9537
rect 91652 9528 91704 9580
rect 83280 9435 83332 9444
rect 83280 9401 83289 9435
rect 83289 9401 83323 9435
rect 83323 9401 83332 9435
rect 83280 9392 83332 9401
rect 85488 9392 85540 9444
rect 89352 9392 89404 9444
rect 88340 9324 88392 9376
rect 88800 9324 88852 9376
rect 90364 9435 90416 9444
rect 90364 9401 90373 9435
rect 90373 9401 90407 9435
rect 90407 9401 90416 9435
rect 90364 9392 90416 9401
rect 92572 9571 92624 9580
rect 92572 9537 92581 9571
rect 92581 9537 92615 9571
rect 92615 9537 92624 9571
rect 92572 9528 92624 9537
rect 93676 9528 93728 9580
rect 94780 9571 94832 9580
rect 94780 9537 94789 9571
rect 94789 9537 94823 9571
rect 94823 9537 94832 9571
rect 94780 9528 94832 9537
rect 94872 9528 94924 9580
rect 96160 9528 96212 9580
rect 96896 9528 96948 9580
rect 98920 9528 98972 9580
rect 103060 9596 103112 9648
rect 108120 9664 108172 9716
rect 113824 9664 113876 9716
rect 121644 9664 121696 9716
rect 121736 9707 121788 9716
rect 121736 9673 121745 9707
rect 121745 9673 121779 9707
rect 121779 9673 121788 9707
rect 121736 9664 121788 9673
rect 125232 9707 125284 9716
rect 125232 9673 125241 9707
rect 125241 9673 125275 9707
rect 125275 9673 125284 9707
rect 125232 9664 125284 9673
rect 126336 9707 126388 9716
rect 126336 9673 126345 9707
rect 126345 9673 126379 9707
rect 126379 9673 126388 9707
rect 126336 9664 126388 9673
rect 129648 9664 129700 9716
rect 130752 9707 130804 9716
rect 130752 9673 130761 9707
rect 130761 9673 130795 9707
rect 130795 9673 130804 9707
rect 130752 9664 130804 9673
rect 131488 9707 131540 9716
rect 131488 9673 131497 9707
rect 131497 9673 131531 9707
rect 131531 9673 131540 9707
rect 131488 9664 131540 9673
rect 133420 9707 133472 9716
rect 133420 9673 133429 9707
rect 133429 9673 133463 9707
rect 133463 9673 133472 9707
rect 133420 9664 133472 9673
rect 134156 9707 134208 9716
rect 134156 9673 134165 9707
rect 134165 9673 134199 9707
rect 134199 9673 134208 9707
rect 134156 9664 134208 9673
rect 117320 9596 117372 9648
rect 123300 9596 123352 9648
rect 131120 9596 131172 9648
rect 158720 9664 158772 9716
rect 147864 9596 147916 9648
rect 155684 9596 155736 9648
rect 164332 9664 164384 9716
rect 100208 9528 100260 9580
rect 100576 9528 100628 9580
rect 100852 9528 100904 9580
rect 101496 9460 101548 9512
rect 103244 9571 103296 9580
rect 103244 9537 103253 9571
rect 103253 9537 103287 9571
rect 103287 9537 103296 9571
rect 103244 9528 103296 9537
rect 103888 9571 103940 9580
rect 103888 9537 103897 9571
rect 103897 9537 103931 9571
rect 103931 9537 103940 9571
rect 103888 9528 103940 9537
rect 104716 9528 104768 9580
rect 105636 9571 105688 9580
rect 105636 9537 105645 9571
rect 105645 9537 105679 9571
rect 105679 9537 105688 9571
rect 105636 9528 105688 9537
rect 106280 9528 106332 9580
rect 107752 9571 107804 9580
rect 107752 9537 107761 9571
rect 107761 9537 107795 9571
rect 107795 9537 107804 9571
rect 107752 9528 107804 9537
rect 108396 9571 108448 9580
rect 108396 9537 108405 9571
rect 108405 9537 108439 9571
rect 108439 9537 108448 9571
rect 108396 9528 108448 9537
rect 109040 9571 109092 9580
rect 109040 9537 109049 9571
rect 109049 9537 109083 9571
rect 109083 9537 109092 9571
rect 109040 9528 109092 9537
rect 110052 9571 110104 9580
rect 110052 9537 110061 9571
rect 110061 9537 110095 9571
rect 110095 9537 110104 9571
rect 110052 9528 110104 9537
rect 110788 9571 110840 9580
rect 110788 9537 110797 9571
rect 110797 9537 110831 9571
rect 110831 9537 110840 9571
rect 110788 9528 110840 9537
rect 111524 9571 111576 9580
rect 111524 9537 111533 9571
rect 111533 9537 111567 9571
rect 111567 9537 111576 9571
rect 111524 9528 111576 9537
rect 112904 9571 112956 9580
rect 112904 9537 112913 9571
rect 112913 9537 112947 9571
rect 112947 9537 112956 9571
rect 112904 9528 112956 9537
rect 113548 9571 113600 9580
rect 113548 9537 113557 9571
rect 113557 9537 113591 9571
rect 113591 9537 113600 9571
rect 113548 9528 113600 9537
rect 114192 9571 114244 9580
rect 114192 9537 114201 9571
rect 114201 9537 114235 9571
rect 114235 9537 114244 9571
rect 114192 9528 114244 9537
rect 115204 9571 115256 9580
rect 115204 9537 115213 9571
rect 115213 9537 115247 9571
rect 115247 9537 115256 9571
rect 115204 9528 115256 9537
rect 115756 9528 115808 9580
rect 116676 9571 116728 9580
rect 116676 9537 116685 9571
rect 116685 9537 116719 9571
rect 116719 9537 116728 9571
rect 116676 9528 116728 9537
rect 118056 9571 118108 9580
rect 118056 9537 118065 9571
rect 118065 9537 118099 9571
rect 118099 9537 118108 9571
rect 118056 9528 118108 9537
rect 118700 9571 118752 9580
rect 118700 9537 118709 9571
rect 118709 9537 118743 9571
rect 118743 9537 118752 9571
rect 118700 9528 118752 9537
rect 119344 9571 119396 9580
rect 119344 9537 119353 9571
rect 119353 9537 119387 9571
rect 119387 9537 119396 9571
rect 119344 9528 119396 9537
rect 120356 9571 120408 9580
rect 120356 9537 120365 9571
rect 120365 9537 120399 9571
rect 120399 9537 120408 9571
rect 120356 9528 120408 9537
rect 121092 9571 121144 9580
rect 121092 9537 121101 9571
rect 121101 9537 121135 9571
rect 121135 9537 121144 9571
rect 121092 9528 121144 9537
rect 121644 9528 121696 9580
rect 124404 9528 124456 9580
rect 126244 9528 126296 9580
rect 128820 9528 128872 9580
rect 129372 9571 129424 9580
rect 129372 9537 129381 9571
rect 129381 9537 129415 9571
rect 129415 9537 129424 9571
rect 129372 9528 129424 9537
rect 130568 9571 130620 9580
rect 130568 9537 130577 9571
rect 130577 9537 130611 9571
rect 130611 9537 130620 9571
rect 130568 9528 130620 9537
rect 131396 9528 131448 9580
rect 133052 9528 133104 9580
rect 134064 9528 134116 9580
rect 138020 9528 138072 9580
rect 138756 9571 138808 9580
rect 138756 9537 138765 9571
rect 138765 9537 138799 9571
rect 138799 9537 138808 9571
rect 138756 9528 138808 9537
rect 139400 9571 139452 9580
rect 139400 9537 139409 9571
rect 139409 9537 139443 9571
rect 139443 9537 139452 9571
rect 139400 9528 139452 9537
rect 140688 9571 140740 9580
rect 140688 9537 140697 9571
rect 140697 9537 140731 9571
rect 140731 9537 140740 9571
rect 140688 9528 140740 9537
rect 141332 9571 141384 9580
rect 141332 9537 141341 9571
rect 141341 9537 141375 9571
rect 141375 9537 141384 9571
rect 141332 9528 141384 9537
rect 141976 9571 142028 9580
rect 141976 9537 141985 9571
rect 141985 9537 142019 9571
rect 142019 9537 142028 9571
rect 141976 9528 142028 9537
rect 143264 9571 143316 9580
rect 143264 9537 143273 9571
rect 143273 9537 143307 9571
rect 143307 9537 143316 9571
rect 143264 9528 143316 9537
rect 143540 9528 143592 9580
rect 144552 9571 144604 9580
rect 144552 9537 144561 9571
rect 144561 9537 144595 9571
rect 144595 9537 144604 9571
rect 144552 9528 144604 9537
rect 145840 9571 145892 9580
rect 145840 9537 145849 9571
rect 145849 9537 145883 9571
rect 145883 9537 145892 9571
rect 145840 9528 145892 9537
rect 146300 9528 146352 9580
rect 147128 9571 147180 9580
rect 147128 9537 147137 9571
rect 147137 9537 147171 9571
rect 147171 9537 147180 9571
rect 147128 9528 147180 9537
rect 148416 9571 148468 9580
rect 148416 9537 148425 9571
rect 148425 9537 148459 9571
rect 148459 9537 148468 9571
rect 148416 9528 148468 9537
rect 149060 9571 149112 9580
rect 149060 9537 149069 9571
rect 149069 9537 149103 9571
rect 149103 9537 149112 9571
rect 149060 9528 149112 9537
rect 149704 9571 149756 9580
rect 149704 9537 149713 9571
rect 149713 9537 149747 9571
rect 149747 9537 149756 9571
rect 149704 9528 149756 9537
rect 150992 9571 151044 9580
rect 150992 9537 151001 9571
rect 151001 9537 151035 9571
rect 151035 9537 151044 9571
rect 150992 9528 151044 9537
rect 151636 9571 151688 9580
rect 151636 9537 151645 9571
rect 151645 9537 151679 9571
rect 151679 9537 151688 9571
rect 151636 9528 151688 9537
rect 152280 9571 152332 9580
rect 152280 9537 152289 9571
rect 152289 9537 152323 9571
rect 152323 9537 152332 9571
rect 152280 9528 152332 9537
rect 152832 9528 152884 9580
rect 154212 9571 154264 9580
rect 154212 9537 154221 9571
rect 154221 9537 154255 9571
rect 154255 9537 154264 9571
rect 154212 9528 154264 9537
rect 154304 9528 154356 9580
rect 92020 9392 92072 9444
rect 108120 9392 108172 9444
rect 127992 9460 128044 9512
rect 152464 9460 152516 9512
rect 157340 9528 157392 9580
rect 157524 9528 157576 9580
rect 161204 9528 161256 9580
rect 161296 9571 161348 9580
rect 161296 9537 161305 9571
rect 161305 9537 161339 9571
rect 161339 9537 161348 9571
rect 161296 9528 161348 9537
rect 162768 9571 162820 9580
rect 162768 9537 162777 9571
rect 162777 9537 162811 9571
rect 162811 9537 162820 9571
rect 162768 9528 162820 9537
rect 166540 9528 166592 9580
rect 166724 9528 166776 9580
rect 166908 9528 166960 9580
rect 168380 9664 168432 9716
rect 168748 9596 168800 9648
rect 215208 9664 215260 9716
rect 218520 9664 218572 9716
rect 220084 9664 220136 9716
rect 224776 9664 224828 9716
rect 225052 9664 225104 9716
rect 258816 9664 258868 9716
rect 259184 9707 259236 9716
rect 259184 9673 259193 9707
rect 259193 9673 259227 9707
rect 259227 9673 259236 9707
rect 259184 9664 259236 9673
rect 171232 9596 171284 9648
rect 169208 9528 169260 9580
rect 171692 9571 171744 9580
rect 171692 9537 171701 9571
rect 171701 9537 171735 9571
rect 171735 9537 171744 9571
rect 171692 9528 171744 9537
rect 172244 9571 172296 9580
rect 172244 9537 172253 9571
rect 172253 9537 172287 9571
rect 172287 9537 172296 9571
rect 172244 9528 172296 9537
rect 173992 9571 174044 9580
rect 173992 9537 174001 9571
rect 174001 9537 174035 9571
rect 174035 9537 174044 9571
rect 173992 9528 174044 9537
rect 174452 9596 174504 9648
rect 175556 9639 175608 9648
rect 175556 9605 175565 9639
rect 175565 9605 175599 9639
rect 175599 9605 175608 9639
rect 175556 9596 175608 9605
rect 220176 9596 220228 9648
rect 220360 9596 220412 9648
rect 175924 9528 175976 9580
rect 177948 9528 178000 9580
rect 178040 9571 178092 9580
rect 178040 9537 178049 9571
rect 178049 9537 178083 9571
rect 178083 9537 178092 9571
rect 178040 9528 178092 9537
rect 179144 9571 179196 9580
rect 179144 9537 179153 9571
rect 179153 9537 179187 9571
rect 179187 9537 179196 9571
rect 179144 9528 179196 9537
rect 109040 9392 109092 9444
rect 109684 9392 109736 9444
rect 112076 9392 112128 9444
rect 116032 9392 116084 9444
rect 121552 9392 121604 9444
rect 132684 9392 132736 9444
rect 103428 9324 103480 9376
rect 103704 9367 103756 9376
rect 103704 9333 103713 9367
rect 103713 9333 103747 9367
rect 103747 9333 103756 9367
rect 103704 9324 103756 9333
rect 104072 9324 104124 9376
rect 108948 9324 109000 9376
rect 110604 9367 110656 9376
rect 110604 9333 110613 9367
rect 110613 9333 110647 9367
rect 110647 9333 110656 9367
rect 110604 9324 110656 9333
rect 112628 9324 112680 9376
rect 113180 9324 113232 9376
rect 115020 9367 115072 9376
rect 115020 9333 115029 9367
rect 115029 9333 115063 9367
rect 115063 9333 115072 9367
rect 115020 9324 115072 9333
rect 115756 9367 115808 9376
rect 115756 9333 115765 9367
rect 115765 9333 115799 9367
rect 115799 9333 115808 9367
rect 115756 9324 115808 9333
rect 115848 9324 115900 9376
rect 117964 9324 118016 9376
rect 118332 9324 118384 9376
rect 119160 9367 119212 9376
rect 119160 9333 119169 9367
rect 119169 9333 119203 9367
rect 119203 9333 119212 9367
rect 119160 9324 119212 9333
rect 120908 9367 120960 9376
rect 120908 9333 120917 9367
rect 120917 9333 120951 9367
rect 120951 9333 120960 9367
rect 120908 9324 120960 9333
rect 128084 9324 128136 9376
rect 128728 9324 128780 9376
rect 142804 9392 142856 9444
rect 145196 9392 145248 9444
rect 148048 9392 148100 9444
rect 138572 9367 138624 9376
rect 138572 9333 138581 9367
rect 138581 9333 138615 9367
rect 138615 9333 138624 9367
rect 138572 9324 138624 9333
rect 140412 9324 140464 9376
rect 140504 9367 140556 9376
rect 140504 9333 140513 9367
rect 140513 9333 140547 9367
rect 140547 9333 140556 9367
rect 140504 9324 140556 9333
rect 140596 9324 140648 9376
rect 142712 9324 142764 9376
rect 143080 9367 143132 9376
rect 143080 9333 143089 9367
rect 143089 9333 143123 9367
rect 143123 9333 143132 9367
rect 143080 9324 143132 9333
rect 144368 9367 144420 9376
rect 144368 9333 144377 9367
rect 144377 9333 144411 9367
rect 144411 9333 144420 9367
rect 144368 9324 144420 9333
rect 145748 9324 145800 9376
rect 150716 9392 150768 9444
rect 153200 9392 153252 9444
rect 156972 9460 157024 9512
rect 158812 9503 158864 9512
rect 158812 9469 158821 9503
rect 158821 9469 158855 9503
rect 158855 9469 158864 9503
rect 158812 9460 158864 9469
rect 159548 9460 159600 9512
rect 159916 9460 159968 9512
rect 161664 9460 161716 9512
rect 161940 9503 161992 9512
rect 161940 9469 161949 9503
rect 161949 9469 161983 9503
rect 161983 9469 161992 9503
rect 161940 9460 161992 9469
rect 162676 9460 162728 9512
rect 163596 9460 163648 9512
rect 164516 9503 164568 9512
rect 164516 9469 164525 9503
rect 164525 9469 164559 9503
rect 164559 9469 164568 9503
rect 164516 9460 164568 9469
rect 165344 9503 165396 9512
rect 165344 9469 165353 9503
rect 165353 9469 165387 9503
rect 165387 9469 165396 9503
rect 165344 9460 165396 9469
rect 165804 9460 165856 9512
rect 167092 9460 167144 9512
rect 169484 9460 169536 9512
rect 148232 9367 148284 9376
rect 148232 9333 148241 9367
rect 148241 9333 148275 9367
rect 148275 9333 148284 9367
rect 148232 9324 148284 9333
rect 148876 9367 148928 9376
rect 148876 9333 148885 9367
rect 148885 9333 148919 9367
rect 148919 9333 148928 9367
rect 148876 9324 148928 9333
rect 150532 9324 150584 9376
rect 150808 9367 150860 9376
rect 150808 9333 150817 9367
rect 150817 9333 150851 9367
rect 150851 9333 150860 9367
rect 150808 9324 150860 9333
rect 153292 9324 153344 9376
rect 154028 9367 154080 9376
rect 154028 9333 154037 9367
rect 154037 9333 154071 9367
rect 154071 9333 154080 9367
rect 154028 9324 154080 9333
rect 156696 9435 156748 9444
rect 156696 9401 156705 9435
rect 156705 9401 156739 9435
rect 156739 9401 156748 9435
rect 156696 9392 156748 9401
rect 155592 9324 155644 9376
rect 155684 9324 155736 9376
rect 169576 9392 169628 9444
rect 171140 9460 171192 9512
rect 172612 9460 172664 9512
rect 180524 9571 180576 9580
rect 180524 9537 180533 9571
rect 180533 9537 180567 9571
rect 180567 9537 180576 9571
rect 180524 9528 180576 9537
rect 180708 9571 180760 9580
rect 180708 9537 180717 9571
rect 180717 9537 180751 9571
rect 180751 9537 180760 9571
rect 180708 9528 180760 9537
rect 181812 9571 181864 9580
rect 181812 9537 181821 9571
rect 181821 9537 181855 9571
rect 181855 9537 181864 9571
rect 181812 9528 181864 9537
rect 182548 9571 182600 9580
rect 182548 9537 182557 9571
rect 182557 9537 182591 9571
rect 182591 9537 182600 9571
rect 182548 9528 182600 9537
rect 183284 9528 183336 9580
rect 185492 9528 185544 9580
rect 188620 9571 188672 9580
rect 188620 9537 188629 9571
rect 188629 9537 188663 9571
rect 188663 9537 188672 9571
rect 188620 9528 188672 9537
rect 190184 9528 190236 9580
rect 190828 9571 190880 9580
rect 190828 9537 190837 9571
rect 190837 9537 190871 9571
rect 190871 9537 190880 9571
rect 190828 9528 190880 9537
rect 192024 9571 192076 9580
rect 192024 9537 192033 9571
rect 192033 9537 192067 9571
rect 192067 9537 192076 9571
rect 192024 9528 192076 9537
rect 192668 9528 192720 9580
rect 194600 9571 194652 9580
rect 194600 9537 194609 9571
rect 194609 9537 194643 9571
rect 194643 9537 194652 9571
rect 194600 9528 194652 9537
rect 195612 9528 195664 9580
rect 197544 9528 197596 9580
rect 197728 9528 197780 9580
rect 202696 9528 202748 9580
rect 203432 9528 203484 9580
rect 205824 9571 205876 9580
rect 205824 9537 205833 9571
rect 205833 9537 205867 9571
rect 205867 9537 205876 9571
rect 205824 9528 205876 9537
rect 206560 9571 206612 9580
rect 206560 9537 206569 9571
rect 206569 9537 206603 9571
rect 206603 9537 206612 9571
rect 206560 9528 206612 9537
rect 207664 9571 207716 9580
rect 207664 9537 207673 9571
rect 207673 9537 207707 9571
rect 207707 9537 207716 9571
rect 207664 9528 207716 9537
rect 208308 9571 208360 9580
rect 208308 9537 208317 9571
rect 208317 9537 208351 9571
rect 208351 9537 208360 9571
rect 208308 9528 208360 9537
rect 208952 9571 209004 9580
rect 208952 9537 208961 9571
rect 208961 9537 208995 9571
rect 208995 9537 209004 9571
rect 208952 9528 209004 9537
rect 209320 9528 209372 9580
rect 210884 9571 210936 9580
rect 210884 9537 210893 9571
rect 210893 9537 210927 9571
rect 210927 9537 210936 9571
rect 210884 9528 210936 9537
rect 211160 9528 211212 9580
rect 212540 9528 212592 9580
rect 213460 9571 213512 9580
rect 213460 9537 213469 9571
rect 213469 9537 213503 9571
rect 213503 9537 213512 9571
rect 213460 9528 213512 9537
rect 213920 9528 213972 9580
rect 214472 9528 214524 9580
rect 215484 9528 215536 9580
rect 216680 9571 216732 9580
rect 216680 9537 216689 9571
rect 216689 9537 216723 9571
rect 216723 9537 216732 9571
rect 216680 9528 216732 9537
rect 217968 9571 218020 9580
rect 217968 9537 217977 9571
rect 217977 9537 218011 9571
rect 218011 9537 218020 9571
rect 217968 9528 218020 9537
rect 218612 9571 218664 9580
rect 218612 9537 218621 9571
rect 218621 9537 218655 9571
rect 218655 9537 218664 9571
rect 218612 9528 218664 9537
rect 219256 9571 219308 9580
rect 219256 9537 219265 9571
rect 219265 9537 219299 9571
rect 219299 9537 219308 9571
rect 219256 9528 219308 9537
rect 220544 9571 220596 9580
rect 220544 9537 220553 9571
rect 220553 9537 220587 9571
rect 220587 9537 220596 9571
rect 220544 9528 220596 9537
rect 229008 9596 229060 9648
rect 221832 9571 221884 9580
rect 221832 9537 221841 9571
rect 221841 9537 221875 9571
rect 221875 9537 221884 9571
rect 221832 9528 221884 9537
rect 223120 9571 223172 9580
rect 223120 9537 223129 9571
rect 223129 9537 223163 9571
rect 223163 9537 223172 9571
rect 223120 9528 223172 9537
rect 223764 9528 223816 9580
rect 223948 9528 224000 9580
rect 224868 9528 224920 9580
rect 227812 9528 227864 9580
rect 228364 9528 228416 9580
rect 228456 9528 228508 9580
rect 230020 9528 230072 9580
rect 230664 9571 230716 9580
rect 230664 9537 230673 9571
rect 230673 9537 230707 9571
rect 230707 9537 230716 9571
rect 230664 9528 230716 9537
rect 230848 9571 230900 9580
rect 230848 9537 230857 9571
rect 230857 9537 230891 9571
rect 230891 9537 230900 9571
rect 230848 9528 230900 9537
rect 232320 9528 232372 9580
rect 233976 9528 234028 9580
rect 234804 9571 234856 9580
rect 234804 9537 234813 9571
rect 234813 9537 234847 9571
rect 234847 9537 234856 9571
rect 234804 9528 234856 9537
rect 239956 9571 240008 9580
rect 239956 9537 239965 9571
rect 239965 9537 239999 9571
rect 239999 9537 240008 9571
rect 239956 9528 240008 9537
rect 240968 9571 241020 9580
rect 240968 9537 240977 9571
rect 240977 9537 241011 9571
rect 241011 9537 241020 9571
rect 240968 9528 241020 9537
rect 242348 9571 242400 9580
rect 242348 9537 242357 9571
rect 242357 9537 242391 9571
rect 242391 9537 242400 9571
rect 242348 9528 242400 9537
rect 242900 9528 242952 9580
rect 169852 9392 169904 9444
rect 158536 9324 158588 9376
rect 160008 9324 160060 9376
rect 162216 9324 162268 9376
rect 162952 9324 163004 9376
rect 163688 9324 163740 9376
rect 164424 9324 164476 9376
rect 165160 9324 165212 9376
rect 165896 9324 165948 9376
rect 166724 9324 166776 9376
rect 169668 9324 169720 9376
rect 175556 9324 175608 9376
rect 178408 9324 178460 9376
rect 184572 9503 184624 9512
rect 184572 9469 184581 9503
rect 184581 9469 184615 9503
rect 184615 9469 184624 9503
rect 184572 9460 184624 9469
rect 186412 9460 186464 9512
rect 187700 9460 187752 9512
rect 184848 9392 184900 9444
rect 197912 9460 197964 9512
rect 219900 9460 219952 9512
rect 219992 9460 220044 9512
rect 191380 9392 191432 9444
rect 192944 9435 192996 9444
rect 192944 9401 192953 9435
rect 192953 9401 192987 9435
rect 192987 9401 192996 9435
rect 192944 9392 192996 9401
rect 194324 9392 194376 9444
rect 195520 9435 195572 9444
rect 195520 9401 195529 9435
rect 195529 9401 195563 9435
rect 195563 9401 195572 9435
rect 195520 9392 195572 9401
rect 196532 9435 196584 9444
rect 196532 9401 196541 9435
rect 196541 9401 196575 9435
rect 196575 9401 196584 9435
rect 196532 9392 196584 9401
rect 197268 9392 197320 9444
rect 202512 9435 202564 9444
rect 202512 9401 202521 9435
rect 202521 9401 202555 9435
rect 202555 9401 202564 9435
rect 202512 9392 202564 9401
rect 207020 9392 207072 9444
rect 215024 9392 215076 9444
rect 215116 9392 215168 9444
rect 186320 9324 186372 9376
rect 190920 9367 190972 9376
rect 190920 9333 190929 9367
rect 190929 9333 190963 9367
rect 190963 9333 190972 9367
rect 190920 9324 190972 9333
rect 194508 9324 194560 9376
rect 197176 9324 197228 9376
rect 202420 9324 202472 9376
rect 206836 9324 206888 9376
rect 207480 9367 207532 9376
rect 207480 9333 207489 9367
rect 207489 9333 207523 9367
rect 207523 9333 207532 9367
rect 207480 9324 207532 9333
rect 208768 9367 208820 9376
rect 208768 9333 208777 9367
rect 208777 9333 208811 9367
rect 208811 9333 208820 9367
rect 208768 9324 208820 9333
rect 210056 9367 210108 9376
rect 210056 9333 210065 9367
rect 210065 9333 210099 9367
rect 210099 9333 210108 9367
rect 210056 9324 210108 9333
rect 210700 9367 210752 9376
rect 210700 9333 210709 9367
rect 210709 9333 210743 9367
rect 210743 9333 210752 9367
rect 210700 9324 210752 9333
rect 212448 9324 212500 9376
rect 212632 9367 212684 9376
rect 212632 9333 212641 9367
rect 212641 9333 212675 9367
rect 212675 9333 212684 9367
rect 212632 9324 212684 9333
rect 213276 9367 213328 9376
rect 213276 9333 213285 9367
rect 213285 9333 213319 9367
rect 213319 9333 213328 9367
rect 213276 9324 213328 9333
rect 214840 9324 214892 9376
rect 217508 9324 217560 9376
rect 217784 9367 217836 9376
rect 217784 9333 217793 9367
rect 217793 9333 217827 9367
rect 217827 9333 217836 9367
rect 217784 9324 217836 9333
rect 218428 9367 218480 9376
rect 218428 9333 218437 9367
rect 218437 9333 218471 9367
rect 218471 9333 218480 9367
rect 218428 9324 218480 9333
rect 219348 9324 219400 9376
rect 220360 9367 220412 9376
rect 220360 9333 220369 9367
rect 220369 9333 220403 9367
rect 220403 9333 220412 9367
rect 220360 9324 220412 9333
rect 221004 9367 221056 9376
rect 221004 9333 221013 9367
rect 221013 9333 221047 9367
rect 221047 9333 221056 9367
rect 221004 9324 221056 9333
rect 221648 9367 221700 9376
rect 221648 9333 221657 9367
rect 221657 9333 221691 9367
rect 221691 9333 221700 9367
rect 221648 9324 221700 9333
rect 222936 9367 222988 9376
rect 222936 9333 222945 9367
rect 222945 9333 222979 9367
rect 222979 9333 222988 9367
rect 222936 9324 222988 9333
rect 224040 9367 224092 9376
rect 224040 9333 224049 9367
rect 224049 9333 224083 9367
rect 224083 9333 224092 9367
rect 224040 9324 224092 9333
rect 225236 9324 225288 9376
rect 228272 9435 228324 9444
rect 228272 9401 228281 9435
rect 228281 9401 228315 9435
rect 228315 9401 228324 9435
rect 228272 9392 228324 9401
rect 229008 9435 229060 9444
rect 229008 9401 229017 9435
rect 229017 9401 229051 9435
rect 229051 9401 229060 9435
rect 229008 9392 229060 9401
rect 229836 9435 229888 9444
rect 229836 9401 229845 9435
rect 229845 9401 229879 9435
rect 229879 9401 229888 9435
rect 229836 9392 229888 9401
rect 230296 9460 230348 9512
rect 235908 9460 235960 9512
rect 230296 9324 230348 9376
rect 231492 9324 231544 9376
rect 231952 9435 232004 9444
rect 231952 9401 231961 9435
rect 231961 9401 231995 9435
rect 231995 9401 232004 9435
rect 231952 9392 232004 9401
rect 233424 9435 233476 9444
rect 233424 9401 233433 9435
rect 233433 9401 233467 9435
rect 233467 9401 233476 9435
rect 233424 9392 233476 9401
rect 236000 9435 236052 9444
rect 236000 9401 236009 9435
rect 236009 9401 236043 9435
rect 236043 9401 236052 9435
rect 236000 9392 236052 9401
rect 237288 9460 237340 9512
rect 242532 9503 242584 9512
rect 242532 9469 242541 9503
rect 242541 9469 242575 9503
rect 242575 9469 242584 9503
rect 242532 9460 242584 9469
rect 243452 9460 243504 9512
rect 244188 9460 244240 9512
rect 246396 9571 246448 9580
rect 246396 9537 246405 9571
rect 246405 9537 246439 9571
rect 246439 9537 246448 9571
rect 246396 9528 246448 9537
rect 247960 9571 248012 9580
rect 247960 9537 247969 9571
rect 247969 9537 248003 9571
rect 248003 9537 248012 9571
rect 247960 9528 248012 9537
rect 249340 9571 249392 9580
rect 249340 9537 249349 9571
rect 249349 9537 249383 9571
rect 249383 9537 249392 9571
rect 249340 9528 249392 9537
rect 251548 9571 251600 9580
rect 251548 9537 251557 9571
rect 251557 9537 251591 9571
rect 251591 9537 251600 9571
rect 251548 9528 251600 9537
rect 253848 9571 253900 9580
rect 253848 9537 253857 9571
rect 253857 9537 253891 9571
rect 253891 9537 253900 9571
rect 253848 9528 253900 9537
rect 246672 9503 246724 9512
rect 246672 9469 246681 9503
rect 246681 9469 246715 9503
rect 246715 9469 246724 9503
rect 246672 9460 246724 9469
rect 249616 9503 249668 9512
rect 249616 9469 249625 9503
rect 249625 9469 249659 9503
rect 249659 9469 249668 9503
rect 249616 9460 249668 9469
rect 249708 9460 249760 9512
rect 254124 9503 254176 9512
rect 254124 9469 254133 9503
rect 254133 9469 254167 9503
rect 254167 9469 254176 9503
rect 254124 9460 254176 9469
rect 255228 9596 255280 9648
rect 266268 9707 266320 9716
rect 266268 9673 266277 9707
rect 266277 9673 266311 9707
rect 266311 9673 266320 9707
rect 266268 9664 266320 9673
rect 267004 9664 267056 9716
rect 270408 9664 270460 9716
rect 264980 9596 265032 9648
rect 255320 9528 255372 9580
rect 257896 9528 257948 9580
rect 257988 9571 258040 9580
rect 257988 9537 257997 9571
rect 257997 9537 258031 9571
rect 258031 9537 258040 9571
rect 257988 9528 258040 9537
rect 256884 9460 256936 9512
rect 259368 9528 259420 9580
rect 260196 9571 260248 9580
rect 260196 9537 260205 9571
rect 260205 9537 260239 9571
rect 260239 9537 260248 9571
rect 260196 9528 260248 9537
rect 259184 9460 259236 9512
rect 263600 9528 263652 9580
rect 264428 9528 264480 9580
rect 265256 9571 265308 9580
rect 265256 9537 265265 9571
rect 265265 9537 265299 9571
rect 265299 9537 265308 9571
rect 269948 9596 270000 9648
rect 265256 9528 265308 9537
rect 238852 9324 238904 9376
rect 240140 9392 240192 9444
rect 258632 9392 258684 9444
rect 258724 9392 258776 9444
rect 261392 9460 261444 9512
rect 261576 9503 261628 9512
rect 261576 9469 261585 9503
rect 261585 9469 261619 9503
rect 261619 9469 261628 9503
rect 261576 9460 261628 9469
rect 262128 9460 262180 9512
rect 263232 9503 263284 9512
rect 263232 9469 263241 9503
rect 263241 9469 263275 9503
rect 263275 9469 263284 9503
rect 263232 9460 263284 9469
rect 263968 9460 264020 9512
rect 264704 9460 264756 9512
rect 267648 9528 267700 9580
rect 268936 9528 268988 9580
rect 260840 9392 260892 9444
rect 263692 9392 263744 9444
rect 263784 9392 263836 9444
rect 266912 9503 266964 9512
rect 266912 9469 266921 9503
rect 266921 9469 266955 9503
rect 266955 9469 266964 9503
rect 266912 9460 266964 9469
rect 267464 9460 267516 9512
rect 267556 9460 267608 9512
rect 268476 9460 268528 9512
rect 268568 9503 268620 9512
rect 268568 9469 268577 9503
rect 268577 9469 268611 9503
rect 268611 9469 268620 9503
rect 268568 9460 268620 9469
rect 268844 9460 268896 9512
rect 270500 9528 270552 9580
rect 269856 9460 269908 9512
rect 244004 9324 244056 9376
rect 245200 9367 245252 9376
rect 245200 9333 245209 9367
rect 245209 9333 245243 9367
rect 245243 9333 245252 9367
rect 245200 9324 245252 9333
rect 245568 9324 245620 9376
rect 258080 9324 258132 9376
rect 261484 9324 261536 9376
rect 261576 9324 261628 9376
rect 262312 9324 262364 9376
rect 264152 9324 264204 9376
rect 265532 9324 265584 9376
rect 268752 9392 268804 9444
rect 270592 9392 270644 9444
rect 266360 9324 266412 9376
rect 269212 9367 269264 9376
rect 269212 9333 269221 9367
rect 269221 9333 269255 9367
rect 269255 9333 269264 9367
rect 269212 9324 269264 9333
rect 269672 9367 269724 9376
rect 269672 9333 269681 9367
rect 269681 9333 269715 9367
rect 269715 9333 269724 9367
rect 269672 9324 269724 9333
rect 34748 9222 34800 9274
rect 34812 9222 34864 9274
rect 34876 9222 34928 9274
rect 34940 9222 34992 9274
rect 35004 9222 35056 9274
rect 102345 9222 102397 9274
rect 102409 9222 102461 9274
rect 102473 9222 102525 9274
rect 102537 9222 102589 9274
rect 102601 9222 102653 9274
rect 169942 9222 169994 9274
rect 170006 9222 170058 9274
rect 170070 9222 170122 9274
rect 170134 9222 170186 9274
rect 170198 9222 170250 9274
rect 237539 9222 237591 9274
rect 237603 9222 237655 9274
rect 237667 9222 237719 9274
rect 237731 9222 237783 9274
rect 237795 9222 237847 9274
rect 1400 9120 1452 9172
rect 3240 9120 3292 9172
rect 7656 9052 7708 9104
rect 5172 8984 5224 9036
rect 17224 8984 17276 9036
rect 3148 8959 3200 8968
rect 3148 8925 3157 8959
rect 3157 8925 3191 8959
rect 3191 8925 3200 8959
rect 3148 8916 3200 8925
rect 8208 8916 8260 8968
rect 13452 8959 13504 8968
rect 13452 8925 13461 8959
rect 13461 8925 13495 8959
rect 13495 8925 13504 8959
rect 13452 8916 13504 8925
rect 14740 8916 14792 8968
rect 18420 8916 18472 8968
rect 20260 8959 20312 8968
rect 20260 8925 20269 8959
rect 20269 8925 20303 8959
rect 20303 8925 20312 8959
rect 20260 8916 20312 8925
rect 3332 8891 3384 8900
rect 3332 8857 3341 8891
rect 3341 8857 3375 8891
rect 3375 8857 3384 8891
rect 3332 8848 3384 8857
rect 8484 8891 8536 8900
rect 8484 8857 8493 8891
rect 8493 8857 8527 8891
rect 8527 8857 8536 8891
rect 8484 8848 8536 8857
rect 13636 8891 13688 8900
rect 13636 8857 13645 8891
rect 13645 8857 13679 8891
rect 13679 8857 13688 8891
rect 13636 8848 13688 8857
rect 7564 8780 7616 8832
rect 19340 8780 19392 8832
rect 21732 8984 21784 9036
rect 23204 9027 23256 9036
rect 23204 8993 23213 9027
rect 23213 8993 23247 9027
rect 23247 8993 23256 9027
rect 23204 8984 23256 8993
rect 21088 8959 21140 8968
rect 21088 8925 21097 8959
rect 21097 8925 21131 8959
rect 21131 8925 21140 8959
rect 21088 8916 21140 8925
rect 21456 8916 21508 8968
rect 21640 8959 21692 8968
rect 21640 8925 21649 8959
rect 21649 8925 21683 8959
rect 21683 8925 21692 8959
rect 21640 8916 21692 8925
rect 21640 8780 21692 8832
rect 22192 8959 22244 8968
rect 22192 8925 22201 8959
rect 22201 8925 22235 8959
rect 22235 8925 22244 8959
rect 22192 8916 22244 8925
rect 22928 8959 22980 8968
rect 22928 8925 22937 8959
rect 22937 8925 22971 8959
rect 22971 8925 22980 8959
rect 22928 8916 22980 8925
rect 23940 9163 23992 9172
rect 23940 9129 23949 9163
rect 23949 9129 23983 9163
rect 23983 9129 23992 9163
rect 23940 9120 23992 9129
rect 30380 9163 30432 9172
rect 30380 9129 30389 9163
rect 30389 9129 30423 9163
rect 30423 9129 30432 9163
rect 30380 9120 30432 9129
rect 32128 9163 32180 9172
rect 32128 9129 32137 9163
rect 32137 9129 32171 9163
rect 32171 9129 32180 9163
rect 32128 9120 32180 9129
rect 33048 9163 33100 9172
rect 33048 9129 33057 9163
rect 33057 9129 33091 9163
rect 33091 9129 33100 9163
rect 33048 9120 33100 9129
rect 35164 9163 35216 9172
rect 35164 9129 35173 9163
rect 35173 9129 35207 9163
rect 35207 9129 35216 9163
rect 35164 9120 35216 9129
rect 53288 9163 53340 9172
rect 53288 9129 53297 9163
rect 53297 9129 53331 9163
rect 53331 9129 53340 9163
rect 53288 9120 53340 9129
rect 53840 9163 53892 9172
rect 53840 9129 53849 9163
rect 53849 9129 53883 9163
rect 53883 9129 53892 9163
rect 53840 9120 53892 9129
rect 54944 9163 54996 9172
rect 54944 9129 54953 9163
rect 54953 9129 54987 9163
rect 54987 9129 54996 9163
rect 54944 9120 54996 9129
rect 55680 9163 55732 9172
rect 55680 9129 55689 9163
rect 55689 9129 55723 9163
rect 55723 9129 55732 9163
rect 55680 9120 55732 9129
rect 56600 9163 56652 9172
rect 56600 9129 56609 9163
rect 56609 9129 56643 9163
rect 56643 9129 56652 9163
rect 56600 9120 56652 9129
rect 58072 9120 58124 9172
rect 58532 9163 58584 9172
rect 58532 9129 58541 9163
rect 58541 9129 58575 9163
rect 58575 9129 58584 9163
rect 58532 9120 58584 9129
rect 62212 9163 62264 9172
rect 62212 9129 62221 9163
rect 62221 9129 62255 9163
rect 62255 9129 62264 9163
rect 62212 9120 62264 9129
rect 62764 9163 62816 9172
rect 62764 9129 62773 9163
rect 62773 9129 62807 9163
rect 62807 9129 62816 9163
rect 62764 9120 62816 9129
rect 64052 9120 64104 9172
rect 24032 9052 24084 9104
rect 41512 9052 41564 9104
rect 46204 9052 46256 9104
rect 57980 9052 58032 9104
rect 62304 9052 62356 9104
rect 73712 9120 73764 9172
rect 84844 9120 84896 9172
rect 88248 9120 88300 9172
rect 90088 9120 90140 9172
rect 90548 9120 90600 9172
rect 91652 9120 91704 9172
rect 91744 9163 91796 9172
rect 91744 9129 91753 9163
rect 91753 9129 91787 9163
rect 91787 9129 91796 9163
rect 91744 9120 91796 9129
rect 93676 9163 93728 9172
rect 93676 9129 93685 9163
rect 93685 9129 93719 9163
rect 93719 9129 93728 9163
rect 93676 9120 93728 9129
rect 24032 8916 24084 8968
rect 23940 8848 23992 8900
rect 24676 8959 24728 8968
rect 24676 8925 24685 8959
rect 24685 8925 24719 8959
rect 24719 8925 24728 8959
rect 24676 8916 24728 8925
rect 25688 8916 25740 8968
rect 27068 8959 27120 8968
rect 27068 8925 27077 8959
rect 27077 8925 27111 8959
rect 27111 8925 27120 8959
rect 27068 8916 27120 8925
rect 27160 8959 27212 8968
rect 27160 8925 27169 8959
rect 27169 8925 27203 8959
rect 27203 8925 27212 8959
rect 27160 8916 27212 8925
rect 27712 8916 27764 8968
rect 28540 8916 28592 8968
rect 30104 8959 30156 8968
rect 30104 8925 30113 8959
rect 30113 8925 30147 8959
rect 30147 8925 30156 8959
rect 30104 8916 30156 8925
rect 30748 8959 30800 8968
rect 30748 8925 30757 8959
rect 30757 8925 30791 8959
rect 30791 8925 30800 8959
rect 30748 8916 30800 8925
rect 31852 8984 31904 9036
rect 32772 8984 32824 9036
rect 32956 8984 33008 9036
rect 31944 8959 31996 8968
rect 31944 8925 31953 8959
rect 31953 8925 31987 8959
rect 31987 8925 31996 8959
rect 31944 8916 31996 8925
rect 33140 8916 33192 8968
rect 40316 8959 40368 8968
rect 40316 8925 40325 8959
rect 40325 8925 40359 8959
rect 40359 8925 40368 8959
rect 40316 8916 40368 8925
rect 36452 8848 36504 8900
rect 22100 8780 22152 8832
rect 22744 8780 22796 8832
rect 24768 8823 24820 8832
rect 24768 8789 24777 8823
rect 24777 8789 24811 8823
rect 24811 8789 24820 8823
rect 24768 8780 24820 8789
rect 27252 8780 27304 8832
rect 27988 8780 28040 8832
rect 28724 8780 28776 8832
rect 30840 8780 30892 8832
rect 32772 8780 32824 8832
rect 39672 8848 39724 8900
rect 45468 8959 45520 8968
rect 45468 8925 45477 8959
rect 45477 8925 45511 8959
rect 45511 8925 45520 8959
rect 45468 8916 45520 8925
rect 53104 8959 53156 8968
rect 53104 8925 53113 8959
rect 53113 8925 53147 8959
rect 53147 8925 53156 8959
rect 53104 8916 53156 8925
rect 53656 8959 53708 8968
rect 53656 8925 53665 8959
rect 53665 8925 53699 8959
rect 53699 8925 53708 8959
rect 53656 8916 53708 8925
rect 54116 8916 54168 8968
rect 54668 8916 54720 8968
rect 55680 8984 55732 9036
rect 55864 8916 55916 8968
rect 56324 8959 56376 8968
rect 56324 8925 56333 8959
rect 56333 8925 56367 8959
rect 56367 8925 56376 8959
rect 56324 8916 56376 8925
rect 56876 8959 56928 8968
rect 56876 8925 56885 8959
rect 56885 8925 56919 8959
rect 56919 8925 56928 8959
rect 56876 8916 56928 8925
rect 57152 8984 57204 9036
rect 57980 8916 58032 8968
rect 58532 8916 58584 8968
rect 60648 9027 60700 9036
rect 60648 8993 60657 9027
rect 60657 8993 60691 9027
rect 60691 8993 60700 9027
rect 60648 8984 60700 8993
rect 59728 8959 59780 8968
rect 59728 8925 59737 8959
rect 59737 8925 59771 8959
rect 59771 8925 59780 8959
rect 59728 8916 59780 8925
rect 59912 8959 59964 8968
rect 59912 8925 59921 8959
rect 59921 8925 59955 8959
rect 59955 8925 59964 8959
rect 59912 8916 59964 8925
rect 61476 8916 61528 8968
rect 62304 8848 62356 8900
rect 62488 8916 62540 8968
rect 63224 8959 63276 8968
rect 63224 8925 63233 8959
rect 63233 8925 63267 8959
rect 63267 8925 63276 8959
rect 63224 8916 63276 8925
rect 64052 8959 64104 8968
rect 64052 8925 64061 8959
rect 64061 8925 64095 8959
rect 64095 8925 64104 8959
rect 64052 8916 64104 8925
rect 64972 8959 65024 8968
rect 64972 8925 64981 8959
rect 64981 8925 65015 8959
rect 65015 8925 65024 8959
rect 64972 8916 65024 8925
rect 65984 8984 66036 9036
rect 66076 8959 66128 8968
rect 66076 8925 66085 8959
rect 66085 8925 66119 8959
rect 66119 8925 66128 8959
rect 66076 8916 66128 8925
rect 66352 8916 66404 8968
rect 70400 8984 70452 9036
rect 72056 9027 72108 9036
rect 72056 8993 72065 9027
rect 72065 8993 72099 9027
rect 72099 8993 72108 9027
rect 72056 8984 72108 8993
rect 73436 9027 73488 9036
rect 73436 8993 73445 9027
rect 73445 8993 73479 9027
rect 73479 8993 73488 9027
rect 73436 8984 73488 8993
rect 81072 9052 81124 9104
rect 94228 9120 94280 9172
rect 96068 9120 96120 9172
rect 96252 9120 96304 9172
rect 96528 9120 96580 9172
rect 97724 9120 97776 9172
rect 98920 9163 98972 9172
rect 98920 9129 98929 9163
rect 98929 9129 98963 9163
rect 98963 9129 98972 9163
rect 98920 9120 98972 9129
rect 100576 9163 100628 9172
rect 100576 9129 100585 9163
rect 100585 9129 100619 9163
rect 100619 9129 100628 9163
rect 100576 9120 100628 9129
rect 101220 9163 101272 9172
rect 101220 9129 101229 9163
rect 101229 9129 101263 9163
rect 101263 9129 101272 9163
rect 101220 9120 101272 9129
rect 107016 9163 107068 9172
rect 107016 9129 107025 9163
rect 107025 9129 107059 9163
rect 107059 9129 107068 9163
rect 107016 9120 107068 9129
rect 111892 9120 111944 9172
rect 115020 9120 115072 9172
rect 121000 9120 121052 9172
rect 94044 9052 94096 9104
rect 103704 9052 103756 9104
rect 104992 9052 105044 9104
rect 108948 9052 109000 9104
rect 111156 9052 111208 9104
rect 115756 9052 115808 9104
rect 121828 9052 121880 9104
rect 124404 9163 124456 9172
rect 124404 9129 124413 9163
rect 124413 9129 124447 9163
rect 124447 9129 124456 9163
rect 124404 9120 124456 9129
rect 124680 9163 124732 9172
rect 124680 9129 124689 9163
rect 124689 9129 124723 9163
rect 124723 9129 124732 9163
rect 124680 9120 124732 9129
rect 126244 9163 126296 9172
rect 126244 9129 126253 9163
rect 126253 9129 126287 9163
rect 126287 9129 126296 9163
rect 126244 9120 126296 9129
rect 127624 9120 127676 9172
rect 128728 9120 128780 9172
rect 130568 9163 130620 9172
rect 130568 9129 130577 9163
rect 130577 9129 130611 9163
rect 130611 9129 130620 9163
rect 130568 9120 130620 9129
rect 131396 9163 131448 9172
rect 131396 9129 131405 9163
rect 131405 9129 131439 9163
rect 131439 9129 131448 9163
rect 131396 9120 131448 9129
rect 133052 9163 133104 9172
rect 133052 9129 133061 9163
rect 133061 9129 133095 9163
rect 133095 9129 133104 9163
rect 133052 9120 133104 9129
rect 134064 9163 134116 9172
rect 134064 9129 134073 9163
rect 134073 9129 134107 9163
rect 134107 9129 134116 9163
rect 134064 9120 134116 9129
rect 134708 9163 134760 9172
rect 134708 9129 134717 9163
rect 134717 9129 134751 9163
rect 134751 9129 134760 9163
rect 134708 9120 134760 9129
rect 142804 9120 142856 9172
rect 148600 9120 148652 9172
rect 152464 9120 152516 9172
rect 175556 9120 175608 9172
rect 176844 9163 176896 9172
rect 176844 9129 176853 9163
rect 176853 9129 176887 9163
rect 176887 9129 176896 9163
rect 176844 9120 176896 9129
rect 177580 9163 177632 9172
rect 177580 9129 177589 9163
rect 177589 9129 177623 9163
rect 177623 9129 177632 9163
rect 177580 9120 177632 9129
rect 81256 9027 81308 9036
rect 81256 8993 81265 9027
rect 81265 8993 81299 9027
rect 81299 8993 81308 9027
rect 81256 8984 81308 8993
rect 81532 9027 81584 9036
rect 81532 8993 81541 9027
rect 81541 8993 81575 9027
rect 81575 8993 81584 9027
rect 81532 8984 81584 8993
rect 66996 8959 67048 8968
rect 66996 8925 67005 8959
rect 67005 8925 67039 8959
rect 67039 8925 67048 8959
rect 66996 8916 67048 8925
rect 70032 8959 70084 8968
rect 70032 8925 70041 8959
rect 70041 8925 70075 8959
rect 70075 8925 70084 8959
rect 70032 8916 70084 8925
rect 72332 8959 72384 8968
rect 72332 8925 72341 8959
rect 72341 8925 72375 8959
rect 72375 8925 72384 8959
rect 72332 8916 72384 8925
rect 73712 8959 73764 8968
rect 73712 8925 73721 8959
rect 73721 8925 73755 8959
rect 73755 8925 73764 8959
rect 73712 8916 73764 8925
rect 74724 8959 74776 8968
rect 74724 8925 74733 8959
rect 74733 8925 74767 8959
rect 74767 8925 74776 8959
rect 74724 8916 74776 8925
rect 75000 8959 75052 8968
rect 75000 8925 75009 8959
rect 75009 8925 75043 8959
rect 75043 8925 75052 8959
rect 75000 8916 75052 8925
rect 77208 8959 77260 8968
rect 77208 8925 77217 8959
rect 77217 8925 77251 8959
rect 77251 8925 77260 8959
rect 77208 8916 77260 8925
rect 77484 8959 77536 8968
rect 77484 8925 77493 8959
rect 77493 8925 77527 8959
rect 77527 8925 77536 8959
rect 77484 8916 77536 8925
rect 78680 8959 78732 8968
rect 78680 8925 78689 8959
rect 78689 8925 78723 8959
rect 78723 8925 78732 8959
rect 78680 8916 78732 8925
rect 78956 8959 79008 8968
rect 78956 8925 78965 8959
rect 78965 8925 78999 8959
rect 78999 8925 79008 8959
rect 78956 8916 79008 8925
rect 62672 8848 62724 8900
rect 82636 8959 82688 8968
rect 82636 8925 82645 8959
rect 82645 8925 82679 8959
rect 82679 8925 82688 8959
rect 82636 8916 82688 8925
rect 82820 9027 82872 9036
rect 82820 8993 82829 9027
rect 82829 8993 82863 9027
rect 82863 8993 82872 9027
rect 82820 8984 82872 8993
rect 86408 9027 86460 9036
rect 86408 8993 86417 9027
rect 86417 8993 86451 9027
rect 86451 8993 86460 9027
rect 86408 8984 86460 8993
rect 89536 8984 89588 9036
rect 86684 8959 86736 8968
rect 86684 8925 86693 8959
rect 86693 8925 86727 8959
rect 86727 8925 86736 8959
rect 86684 8916 86736 8925
rect 89076 8959 89128 8968
rect 89076 8925 89085 8959
rect 89085 8925 89119 8959
rect 89119 8925 89128 8959
rect 89076 8916 89128 8925
rect 89444 8916 89496 8968
rect 89904 8959 89956 8968
rect 89904 8925 89913 8959
rect 89913 8925 89947 8959
rect 89947 8925 89956 8959
rect 89904 8916 89956 8925
rect 89996 8959 90048 8968
rect 89996 8925 90005 8959
rect 90005 8925 90039 8959
rect 90039 8925 90048 8959
rect 89996 8916 90048 8925
rect 90732 8959 90784 8968
rect 90732 8925 90741 8959
rect 90741 8925 90775 8959
rect 90775 8925 90784 8959
rect 90732 8916 90784 8925
rect 39396 8780 39448 8832
rect 44732 8780 44784 8832
rect 54116 8780 54168 8832
rect 56876 8780 56928 8832
rect 57428 8780 57480 8832
rect 58256 8823 58308 8832
rect 58256 8789 58265 8823
rect 58265 8789 58299 8823
rect 58299 8789 58308 8823
rect 58256 8780 58308 8789
rect 59360 8780 59412 8832
rect 60096 8823 60148 8832
rect 60096 8789 60105 8823
rect 60105 8789 60139 8823
rect 60139 8789 60148 8823
rect 60096 8780 60148 8789
rect 60832 8780 60884 8832
rect 61476 8823 61528 8832
rect 61476 8789 61485 8823
rect 61485 8789 61519 8823
rect 61519 8789 61528 8823
rect 61476 8780 61528 8789
rect 63776 8780 63828 8832
rect 64512 8780 64564 8832
rect 65340 8780 65392 8832
rect 66076 8780 66128 8832
rect 67180 8823 67232 8832
rect 67180 8789 67189 8823
rect 67189 8789 67223 8823
rect 67223 8789 67232 8823
rect 67180 8780 67232 8789
rect 91100 8848 91152 8900
rect 91652 8916 91704 8968
rect 92388 8959 92440 8968
rect 92388 8925 92397 8959
rect 92397 8925 92431 8959
rect 92431 8925 92440 8959
rect 92388 8916 92440 8925
rect 92848 8916 92900 8968
rect 93400 8959 93452 8968
rect 93400 8925 93409 8959
rect 93409 8925 93443 8959
rect 93443 8925 93452 8959
rect 93400 8916 93452 8925
rect 93492 8959 93544 8968
rect 93492 8925 93501 8959
rect 93501 8925 93535 8959
rect 93535 8925 93544 8959
rect 93492 8916 93544 8925
rect 94596 8984 94648 9036
rect 92940 8848 92992 8900
rect 93124 8848 93176 8900
rect 94872 8916 94924 8968
rect 95240 8984 95292 9036
rect 95976 9027 96028 9036
rect 95976 8993 95985 9027
rect 95985 8993 96019 9027
rect 96019 8993 96028 9027
rect 95976 8984 96028 8993
rect 96528 8984 96580 9036
rect 99196 9027 99248 9036
rect 99196 8993 99205 9027
rect 99205 8993 99239 9027
rect 99239 8993 99248 9027
rect 99196 8984 99248 8993
rect 99288 8984 99340 9036
rect 123300 8984 123352 9036
rect 123484 8984 123536 9036
rect 96620 8916 96672 8968
rect 96988 8959 97040 8968
rect 96988 8925 96997 8959
rect 96997 8925 97031 8959
rect 97031 8925 97040 8959
rect 96988 8916 97040 8925
rect 89536 8780 89588 8832
rect 90548 8780 90600 8832
rect 90640 8780 90692 8832
rect 94412 8780 94464 8832
rect 94872 8780 94924 8832
rect 96068 8780 96120 8832
rect 97724 8959 97776 8968
rect 97724 8925 97733 8959
rect 97733 8925 97767 8959
rect 97767 8925 97776 8959
rect 97724 8916 97776 8925
rect 97356 8848 97408 8900
rect 97540 8848 97592 8900
rect 98092 8959 98144 8968
rect 98092 8925 98101 8959
rect 98101 8925 98135 8959
rect 98135 8925 98144 8959
rect 98092 8916 98144 8925
rect 98552 8959 98604 8968
rect 98552 8925 98561 8959
rect 98561 8925 98595 8959
rect 98595 8925 98604 8959
rect 98552 8916 98604 8925
rect 100300 8959 100352 8968
rect 100300 8925 100309 8959
rect 100309 8925 100343 8959
rect 100343 8925 100352 8959
rect 100300 8916 100352 8925
rect 100944 8916 100996 8968
rect 101036 8959 101088 8968
rect 101036 8925 101045 8959
rect 101045 8925 101079 8959
rect 101079 8925 101088 8959
rect 101036 8916 101088 8925
rect 101496 8916 101548 8968
rect 106372 8916 106424 8968
rect 107200 8959 107252 8968
rect 107200 8925 107209 8959
rect 107209 8925 107243 8959
rect 107243 8925 107252 8959
rect 107200 8916 107252 8925
rect 112352 8959 112404 8968
rect 112352 8925 112361 8959
rect 112361 8925 112395 8959
rect 112395 8925 112404 8959
rect 112352 8916 112404 8925
rect 117228 8916 117280 8968
rect 121000 8916 121052 8968
rect 105084 8848 105136 8900
rect 110604 8848 110656 8900
rect 97264 8823 97316 8832
rect 97264 8789 97273 8823
rect 97273 8789 97307 8823
rect 97307 8789 97316 8823
rect 97264 8780 97316 8789
rect 99656 8780 99708 8832
rect 100208 8780 100260 8832
rect 111340 8780 111392 8832
rect 112168 8823 112220 8832
rect 112168 8789 112177 8823
rect 112177 8789 112211 8823
rect 112211 8789 112220 8823
rect 112168 8780 112220 8789
rect 116492 8780 116544 8832
rect 122656 8959 122708 8968
rect 122656 8925 122665 8959
rect 122665 8925 122699 8959
rect 122699 8925 122708 8959
rect 122656 8916 122708 8925
rect 121828 8848 121880 8900
rect 124128 8959 124180 8968
rect 124128 8925 124137 8959
rect 124137 8925 124171 8959
rect 124171 8925 124180 8959
rect 124128 8916 124180 8925
rect 124680 8916 124732 8968
rect 125048 8959 125100 8968
rect 125048 8925 125057 8959
rect 125057 8925 125091 8959
rect 125091 8925 125100 8959
rect 125048 8916 125100 8925
rect 125876 8959 125928 8968
rect 125876 8925 125885 8959
rect 125885 8925 125919 8959
rect 125919 8925 125928 8959
rect 125876 8916 125928 8925
rect 126336 8916 126388 8968
rect 126704 8959 126756 8968
rect 126704 8925 126713 8959
rect 126713 8925 126747 8959
rect 126747 8925 126756 8959
rect 126704 8916 126756 8925
rect 127624 8959 127676 8968
rect 127624 8925 127633 8959
rect 127633 8925 127667 8959
rect 127667 8925 127676 8959
rect 127624 8916 127676 8925
rect 127808 8959 127860 8968
rect 127808 8925 127817 8959
rect 127817 8925 127851 8959
rect 127851 8925 127860 8959
rect 127808 8916 127860 8925
rect 122840 8848 122892 8900
rect 123392 8848 123444 8900
rect 133880 9052 133932 9104
rect 141424 9052 141476 9104
rect 169668 9052 169720 9104
rect 169760 9052 169812 9104
rect 174268 9095 174320 9104
rect 174268 9061 174277 9095
rect 174277 9061 174311 9095
rect 174311 9061 174320 9095
rect 174268 9052 174320 9061
rect 175280 9052 175332 9104
rect 184572 9120 184624 9172
rect 192024 9120 192076 9172
rect 194600 9120 194652 9172
rect 198004 9120 198056 9172
rect 199752 9120 199804 9172
rect 200120 9120 200172 9172
rect 200672 9120 200724 9172
rect 203340 9120 203392 9172
rect 203432 9163 203484 9172
rect 203432 9129 203441 9163
rect 203441 9129 203475 9163
rect 203475 9129 203484 9163
rect 203432 9120 203484 9129
rect 204076 9163 204128 9172
rect 204076 9129 204085 9163
rect 204085 9129 204119 9163
rect 204119 9129 204128 9163
rect 204076 9120 204128 9129
rect 182088 9095 182140 9104
rect 182088 9061 182097 9095
rect 182097 9061 182131 9095
rect 182131 9061 182140 9095
rect 182088 9052 182140 9061
rect 128820 9027 128872 9036
rect 128820 8993 128829 9027
rect 128829 8993 128863 9027
rect 128863 8993 128872 9027
rect 128820 8984 128872 8993
rect 130108 8916 130160 8968
rect 131120 8916 131172 8968
rect 131856 8959 131908 8968
rect 131856 8925 131865 8959
rect 131865 8925 131899 8959
rect 131899 8925 131908 8959
rect 131856 8916 131908 8925
rect 132592 8916 132644 8968
rect 132776 8959 132828 8968
rect 132776 8925 132785 8959
rect 132785 8925 132819 8959
rect 132819 8925 132828 8959
rect 132776 8916 132828 8925
rect 132868 8959 132920 8968
rect 132868 8925 132877 8959
rect 132877 8925 132911 8959
rect 132911 8925 132920 8959
rect 132868 8916 132920 8925
rect 133788 8959 133840 8968
rect 133788 8925 133797 8959
rect 133797 8925 133831 8959
rect 133831 8925 133840 8959
rect 133788 8916 133840 8925
rect 134524 8959 134576 8968
rect 134524 8925 134533 8959
rect 134533 8925 134567 8959
rect 134567 8925 134576 8959
rect 134524 8916 134576 8925
rect 130844 8848 130896 8900
rect 145012 8984 145064 9036
rect 149612 8984 149664 9036
rect 139768 8959 139820 8968
rect 139768 8925 139777 8959
rect 139777 8925 139811 8959
rect 139811 8925 139820 8959
rect 139768 8916 139820 8925
rect 144920 8959 144972 8968
rect 144920 8925 144929 8959
rect 144929 8925 144963 8959
rect 144963 8925 144972 8959
rect 144920 8916 144972 8925
rect 150072 8959 150124 8968
rect 150072 8925 150081 8959
rect 150081 8925 150115 8959
rect 150115 8925 150124 8959
rect 150072 8916 150124 8925
rect 150808 8984 150860 9036
rect 153476 8984 153528 9036
rect 156052 8984 156104 9036
rect 156696 8984 156748 9036
rect 157340 9027 157392 9036
rect 157340 8993 157349 9027
rect 157349 8993 157383 9027
rect 157383 8993 157392 9027
rect 157340 8984 157392 8993
rect 157432 8984 157484 9036
rect 155224 8959 155276 8968
rect 155224 8925 155233 8959
rect 155233 8925 155267 8959
rect 155267 8925 155276 8959
rect 155224 8916 155276 8925
rect 142804 8848 142856 8900
rect 156236 8848 156288 8900
rect 157064 8959 157116 8968
rect 157064 8925 157073 8959
rect 157073 8925 157107 8959
rect 157107 8925 157116 8959
rect 157064 8916 157116 8925
rect 157524 8916 157576 8968
rect 159640 8959 159692 8968
rect 159640 8925 159649 8959
rect 159649 8925 159683 8959
rect 159683 8925 159692 8959
rect 159640 8916 159692 8925
rect 157800 8848 157852 8900
rect 159180 8891 159232 8900
rect 159180 8857 159189 8891
rect 159189 8857 159223 8891
rect 159223 8857 159232 8891
rect 159180 8848 159232 8857
rect 161112 8848 161164 8900
rect 161940 8959 161992 8968
rect 161940 8925 161949 8959
rect 161949 8925 161983 8959
rect 161983 8925 161992 8959
rect 161940 8916 161992 8925
rect 162860 8916 162912 8968
rect 163780 8959 163832 8968
rect 163780 8925 163789 8959
rect 163789 8925 163823 8959
rect 163823 8925 163832 8959
rect 163780 8916 163832 8925
rect 162308 8891 162360 8900
rect 162308 8857 162317 8891
rect 162317 8857 162351 8891
rect 162351 8857 162360 8891
rect 162308 8848 162360 8857
rect 162584 8848 162636 8900
rect 162768 8848 162820 8900
rect 164516 8848 164568 8900
rect 121736 8780 121788 8832
rect 122196 8780 122248 8832
rect 123024 8780 123076 8832
rect 123852 8780 123904 8832
rect 125416 8823 125468 8832
rect 125416 8789 125425 8823
rect 125425 8789 125459 8823
rect 125459 8789 125468 8823
rect 125416 8780 125468 8789
rect 126796 8780 126848 8832
rect 127532 8780 127584 8832
rect 131948 8780 132000 8832
rect 133880 8780 133932 8832
rect 134156 8780 134208 8832
rect 139308 8780 139360 8832
rect 144736 8823 144788 8832
rect 144736 8789 144745 8823
rect 144745 8789 144779 8823
rect 144779 8789 144788 8823
rect 144736 8780 144788 8789
rect 150348 8780 150400 8832
rect 155040 8823 155092 8832
rect 155040 8789 155049 8823
rect 155049 8789 155083 8823
rect 155083 8789 155092 8823
rect 155040 8780 155092 8789
rect 155960 8780 156012 8832
rect 161848 8780 161900 8832
rect 165804 8780 165856 8832
rect 166172 8959 166224 8968
rect 166172 8925 166181 8959
rect 166181 8925 166215 8959
rect 166215 8925 166224 8959
rect 166172 8916 166224 8925
rect 166448 8916 166500 8968
rect 168748 8916 168800 8968
rect 168932 8959 168984 8968
rect 168932 8925 168941 8959
rect 168941 8925 168975 8959
rect 168975 8925 168984 8959
rect 168932 8916 168984 8925
rect 169024 8916 169076 8968
rect 167092 8848 167144 8900
rect 167828 8848 167880 8900
rect 171876 8984 171928 9036
rect 194508 9052 194560 9104
rect 194692 9052 194744 9104
rect 195336 9052 195388 9104
rect 195520 9052 195572 9104
rect 184296 9027 184348 9036
rect 184296 8993 184305 9027
rect 184305 8993 184339 9027
rect 184339 8993 184348 9027
rect 184296 8984 184348 8993
rect 184756 8984 184808 9036
rect 186228 8984 186280 9036
rect 189448 9027 189500 9036
rect 189448 8993 189457 9027
rect 189457 8993 189491 9027
rect 189491 8993 189500 9027
rect 189448 8984 189500 8993
rect 190828 8984 190880 9036
rect 197728 8984 197780 9036
rect 201316 9052 201368 9104
rect 204260 9052 204312 9104
rect 220268 9052 220320 9104
rect 173900 8916 173952 8968
rect 175188 8916 175240 8968
rect 176752 8959 176804 8968
rect 176752 8925 176761 8959
rect 176761 8925 176795 8959
rect 176795 8925 176804 8959
rect 176752 8916 176804 8925
rect 177488 8959 177540 8968
rect 177488 8925 177497 8959
rect 177497 8925 177531 8959
rect 177531 8925 177540 8959
rect 177488 8916 177540 8925
rect 180432 8959 180484 8968
rect 180432 8925 180441 8959
rect 180441 8925 180475 8959
rect 180475 8925 180484 8959
rect 180432 8916 180484 8925
rect 181904 8959 181956 8968
rect 181904 8925 181913 8959
rect 181913 8925 181947 8959
rect 181947 8925 181956 8959
rect 181904 8916 181956 8925
rect 185860 8959 185912 8968
rect 185860 8925 185869 8959
rect 185869 8925 185903 8959
rect 185903 8925 185912 8959
rect 185860 8916 185912 8925
rect 168840 8780 168892 8832
rect 168932 8780 168984 8832
rect 171048 8780 171100 8832
rect 172704 8780 172756 8832
rect 177672 8780 177724 8832
rect 182088 8780 182140 8832
rect 189724 8959 189776 8968
rect 189724 8925 189733 8959
rect 189733 8925 189767 8959
rect 189767 8925 189776 8959
rect 189724 8916 189776 8925
rect 190644 8916 190696 8968
rect 190920 8959 190972 8968
rect 190920 8925 190929 8959
rect 190929 8925 190963 8959
rect 190963 8925 190972 8959
rect 190920 8916 190972 8925
rect 191012 8916 191064 8968
rect 192116 8916 192168 8968
rect 192484 8848 192536 8900
rect 193312 8959 193364 8968
rect 193312 8925 193321 8959
rect 193321 8925 193355 8959
rect 193355 8925 193364 8959
rect 193312 8916 193364 8925
rect 194692 8959 194744 8968
rect 194692 8925 194701 8959
rect 194701 8925 194735 8959
rect 194735 8925 194744 8959
rect 194692 8916 194744 8925
rect 195520 8959 195572 8968
rect 195520 8925 195529 8959
rect 195529 8925 195563 8959
rect 195563 8925 195572 8959
rect 195520 8916 195572 8925
rect 196348 8959 196400 8968
rect 196348 8925 196357 8959
rect 196357 8925 196391 8959
rect 196391 8925 196400 8959
rect 196348 8916 196400 8925
rect 195980 8848 196032 8900
rect 198556 8916 198608 8968
rect 199752 8959 199804 8968
rect 199752 8925 199761 8959
rect 199761 8925 199795 8959
rect 199795 8925 199804 8959
rect 199752 8916 199804 8925
rect 220084 8984 220136 9036
rect 220176 8984 220228 9036
rect 223672 9052 223724 9104
rect 223764 9095 223816 9104
rect 223764 9061 223773 9095
rect 223773 9061 223807 9095
rect 223807 9061 223816 9095
rect 223764 9052 223816 9061
rect 221648 8984 221700 9036
rect 225420 9052 225472 9104
rect 228364 9163 228416 9172
rect 228364 9129 228373 9163
rect 228373 9129 228407 9163
rect 228407 9129 228416 9163
rect 228364 9120 228416 9129
rect 228548 9120 228600 9172
rect 230572 9052 230624 9104
rect 230940 9120 230992 9172
rect 233976 9163 234028 9172
rect 233976 9129 233985 9163
rect 233985 9129 234019 9163
rect 234019 9129 234028 9163
rect 233976 9120 234028 9129
rect 234712 9120 234764 9172
rect 235632 9120 235684 9172
rect 236460 9120 236512 9172
rect 236828 9163 236880 9172
rect 236828 9129 236837 9163
rect 236837 9129 236871 9163
rect 236871 9129 236880 9163
rect 236828 9120 236880 9129
rect 244924 9120 244976 9172
rect 249708 9120 249760 9172
rect 249800 9120 249852 9172
rect 254676 9120 254728 9172
rect 258724 9120 258776 9172
rect 259368 9163 259420 9172
rect 259368 9129 259377 9163
rect 259377 9129 259411 9163
rect 259411 9129 259420 9163
rect 259368 9120 259420 9129
rect 261668 9120 261720 9172
rect 262128 9120 262180 9172
rect 265072 9120 265124 9172
rect 268660 9120 268712 9172
rect 270408 9120 270460 9172
rect 200672 8959 200724 8968
rect 200672 8925 200681 8959
rect 200681 8925 200715 8959
rect 200715 8925 200724 8959
rect 200672 8916 200724 8925
rect 201316 8916 201368 8968
rect 202328 8959 202380 8968
rect 202328 8925 202337 8959
rect 202337 8925 202371 8959
rect 202371 8925 202380 8959
rect 202328 8916 202380 8925
rect 203064 8959 203116 8968
rect 203064 8925 203073 8959
rect 203073 8925 203107 8959
rect 203107 8925 203116 8959
rect 203064 8916 203116 8925
rect 202512 8848 202564 8900
rect 203524 8916 203576 8968
rect 211712 8959 211764 8968
rect 211712 8925 211721 8959
rect 211721 8925 211755 8959
rect 211755 8925 211764 8959
rect 211712 8916 211764 8925
rect 211804 8916 211856 8968
rect 215116 8916 215168 8968
rect 216864 8959 216916 8968
rect 216864 8925 216873 8959
rect 216873 8925 216907 8959
rect 216907 8925 216916 8959
rect 216864 8916 216916 8925
rect 222016 8959 222068 8968
rect 222016 8925 222025 8959
rect 222025 8925 222059 8959
rect 222059 8925 222068 8959
rect 222016 8916 222068 8925
rect 223028 8916 223080 8968
rect 224592 8984 224644 9036
rect 232780 9027 232832 9036
rect 232780 8993 232789 9027
rect 232789 8993 232823 9027
rect 232823 8993 232832 9027
rect 232780 8984 232832 8993
rect 254768 9052 254820 9104
rect 254952 9052 255004 9104
rect 263232 9052 263284 9104
rect 263692 9052 263744 9104
rect 267924 9052 267976 9104
rect 268476 9052 268528 9104
rect 254676 8984 254728 9036
rect 255044 9027 255096 9036
rect 255044 8993 255053 9027
rect 255053 8993 255087 9027
rect 255087 8993 255096 9027
rect 255044 8984 255096 8993
rect 256424 9027 256476 9036
rect 256424 8993 256433 9027
rect 256433 8993 256467 9027
rect 256467 8993 256476 9027
rect 256424 8984 256476 8993
rect 257712 9027 257764 9036
rect 257712 8993 257721 9027
rect 257721 8993 257755 9027
rect 257755 8993 257764 9027
rect 257712 8984 257764 8993
rect 257896 8984 257948 9036
rect 260748 8984 260800 9036
rect 224316 8959 224368 8968
rect 224316 8925 224325 8959
rect 224325 8925 224359 8959
rect 224359 8925 224368 8959
rect 224316 8916 224368 8925
rect 224408 8959 224460 8968
rect 224408 8925 224417 8959
rect 224417 8925 224451 8959
rect 224451 8925 224460 8959
rect 224408 8916 224460 8925
rect 203340 8848 203392 8900
rect 225144 8848 225196 8900
rect 225604 8959 225656 8968
rect 225604 8925 225613 8959
rect 225613 8925 225647 8959
rect 225647 8925 225656 8959
rect 225604 8916 225656 8925
rect 226432 8959 226484 8968
rect 226432 8925 226441 8959
rect 226441 8925 226475 8959
rect 226475 8925 226484 8959
rect 226432 8916 226484 8925
rect 227168 8959 227220 8968
rect 227168 8925 227177 8959
rect 227177 8925 227211 8959
rect 227211 8925 227220 8959
rect 227168 8916 227220 8925
rect 228088 8959 228140 8968
rect 228088 8925 228097 8959
rect 228097 8925 228131 8959
rect 228131 8925 228140 8959
rect 228088 8916 228140 8925
rect 228824 8959 228876 8968
rect 228824 8925 228833 8959
rect 228833 8925 228867 8959
rect 228867 8925 228876 8959
rect 228824 8916 228876 8925
rect 228272 8848 228324 8900
rect 229652 8959 229704 8968
rect 229652 8925 229661 8959
rect 229661 8925 229695 8959
rect 229695 8925 229704 8959
rect 229652 8916 229704 8925
rect 230020 8959 230072 8968
rect 230020 8925 230029 8959
rect 230029 8925 230063 8959
rect 230063 8925 230072 8959
rect 230020 8916 230072 8925
rect 230112 8916 230164 8968
rect 230848 8916 230900 8968
rect 230204 8848 230256 8900
rect 230664 8848 230716 8900
rect 231860 8916 231912 8968
rect 232044 8916 232096 8968
rect 232320 8959 232372 8968
rect 232320 8925 232329 8959
rect 232329 8925 232363 8959
rect 232363 8925 232372 8959
rect 232320 8916 232372 8925
rect 233608 8959 233660 8968
rect 233608 8925 233617 8959
rect 233617 8925 233651 8959
rect 233651 8925 233660 8959
rect 233608 8916 233660 8925
rect 233700 8848 233752 8900
rect 234528 8959 234580 8968
rect 234528 8925 234537 8959
rect 234537 8925 234571 8959
rect 234571 8925 234580 8959
rect 234528 8916 234580 8925
rect 234804 8916 234856 8968
rect 235816 8959 235868 8968
rect 235816 8925 235825 8959
rect 235825 8925 235859 8959
rect 235859 8925 235868 8959
rect 235816 8916 235868 8925
rect 241244 8959 241296 8968
rect 241244 8925 241253 8959
rect 241253 8925 241287 8959
rect 241287 8925 241296 8959
rect 241244 8916 241296 8925
rect 241612 8916 241664 8968
rect 245016 8959 245068 8968
rect 245016 8925 245025 8959
rect 245025 8925 245059 8959
rect 245059 8925 245068 8959
rect 245016 8916 245068 8925
rect 246212 8959 246264 8968
rect 246212 8925 246221 8959
rect 246221 8925 246255 8959
rect 246255 8925 246264 8959
rect 246212 8916 246264 8925
rect 247132 8959 247184 8968
rect 247132 8925 247141 8959
rect 247141 8925 247175 8959
rect 247175 8925 247184 8959
rect 247132 8916 247184 8925
rect 247408 8959 247460 8968
rect 247408 8925 247417 8959
rect 247417 8925 247451 8959
rect 247451 8925 247460 8959
rect 247408 8916 247460 8925
rect 248696 8959 248748 8968
rect 248696 8925 248705 8959
rect 248705 8925 248739 8959
rect 248739 8925 248748 8959
rect 248696 8916 248748 8925
rect 250168 8959 250220 8968
rect 250168 8925 250177 8959
rect 250177 8925 250211 8959
rect 250211 8925 250220 8959
rect 250168 8916 250220 8925
rect 251180 8916 251232 8968
rect 252284 8959 252336 8968
rect 252284 8925 252293 8959
rect 252293 8925 252327 8959
rect 252327 8925 252336 8959
rect 252284 8916 252336 8925
rect 253756 8959 253808 8968
rect 253756 8925 253765 8959
rect 253765 8925 253799 8959
rect 253799 8925 253808 8959
rect 253756 8916 253808 8925
rect 238852 8848 238904 8900
rect 246948 8848 247000 8900
rect 249064 8848 249116 8900
rect 255320 8959 255372 8968
rect 255320 8925 255329 8959
rect 255329 8925 255363 8959
rect 255363 8925 255372 8959
rect 255320 8916 255372 8925
rect 256792 8916 256844 8968
rect 190368 8780 190420 8832
rect 191932 8823 191984 8832
rect 191932 8789 191941 8823
rect 191941 8789 191975 8823
rect 191975 8789 191984 8823
rect 191932 8780 191984 8789
rect 193128 8780 193180 8832
rect 193864 8780 193916 8832
rect 195336 8823 195388 8832
rect 195336 8789 195345 8823
rect 195345 8789 195379 8823
rect 195379 8789 195388 8823
rect 195336 8780 195388 8789
rect 196072 8780 196124 8832
rect 199200 8780 199252 8832
rect 200212 8780 200264 8832
rect 201040 8780 201092 8832
rect 201868 8780 201920 8832
rect 214564 8780 214616 8832
rect 217692 8780 217744 8832
rect 217968 8780 218020 8832
rect 221280 8780 221332 8832
rect 223396 8780 223448 8832
rect 224500 8780 224552 8832
rect 225328 8780 225380 8832
rect 226064 8780 226116 8832
rect 226800 8780 226852 8832
rect 228088 8780 228140 8832
rect 228548 8780 228600 8832
rect 229008 8780 229060 8832
rect 231308 8780 231360 8832
rect 232412 8780 232464 8832
rect 234712 8780 234764 8832
rect 245108 8823 245160 8832
rect 245108 8789 245117 8823
rect 245117 8789 245151 8823
rect 245151 8789 245160 8823
rect 245108 8780 245160 8789
rect 246304 8823 246356 8832
rect 246304 8789 246313 8823
rect 246313 8789 246347 8823
rect 246347 8789 246356 8823
rect 246304 8780 246356 8789
rect 247040 8780 247092 8832
rect 250260 8823 250312 8832
rect 250260 8789 250269 8823
rect 250269 8789 250303 8823
rect 250303 8789 250312 8823
rect 250260 8780 250312 8789
rect 250352 8780 250404 8832
rect 251548 8780 251600 8832
rect 259092 8959 259144 8968
rect 259092 8925 259101 8959
rect 259101 8925 259135 8959
rect 259135 8925 259144 8959
rect 259092 8916 259144 8925
rect 259184 8959 259236 8968
rect 259184 8925 259193 8959
rect 259193 8925 259227 8959
rect 259227 8925 259236 8959
rect 259184 8916 259236 8925
rect 259828 8959 259880 8968
rect 259828 8925 259837 8959
rect 259837 8925 259871 8959
rect 259871 8925 259880 8959
rect 259828 8916 259880 8925
rect 260564 8916 260616 8968
rect 264060 8984 264112 9036
rect 267188 8984 267240 9036
rect 267280 8984 267332 9036
rect 269672 8984 269724 9036
rect 262956 8916 263008 8968
rect 263600 8959 263652 8968
rect 263600 8925 263609 8959
rect 263609 8925 263643 8959
rect 263643 8925 263652 8959
rect 263600 8916 263652 8925
rect 263876 8916 263928 8968
rect 265256 8916 265308 8968
rect 266452 8916 266504 8968
rect 267924 8916 267976 8968
rect 262036 8848 262088 8900
rect 266728 8848 266780 8900
rect 267188 8848 267240 8900
rect 267372 8848 267424 8900
rect 268016 8848 268068 8900
rect 270868 8848 270920 8900
rect 259736 8780 259788 8832
rect 260288 8780 260340 8832
rect 263140 8780 263192 8832
rect 266452 8780 266504 8832
rect 266544 8780 266596 8832
rect 267464 8780 267516 8832
rect 269028 8780 269080 8832
rect 269212 8780 269264 8832
rect 270408 8780 270460 8832
rect 68546 8678 68598 8730
rect 68610 8678 68662 8730
rect 68674 8678 68726 8730
rect 68738 8678 68790 8730
rect 68802 8678 68854 8730
rect 136143 8678 136195 8730
rect 136207 8678 136259 8730
rect 136271 8678 136323 8730
rect 136335 8678 136387 8730
rect 136399 8678 136451 8730
rect 203740 8678 203792 8730
rect 203804 8678 203856 8730
rect 203868 8678 203920 8730
rect 203932 8678 203984 8730
rect 203996 8678 204048 8730
rect 271337 8678 271389 8730
rect 271401 8678 271453 8730
rect 271465 8678 271517 8730
rect 271529 8678 271581 8730
rect 271593 8678 271645 8730
rect 10324 8576 10376 8628
rect 20812 8576 20864 8628
rect 21364 8619 21416 8628
rect 21364 8585 21373 8619
rect 21373 8585 21407 8619
rect 21407 8585 21416 8619
rect 21364 8576 21416 8585
rect 21456 8576 21508 8628
rect 22192 8576 22244 8628
rect 24032 8619 24084 8628
rect 24032 8585 24041 8619
rect 24041 8585 24075 8619
rect 24075 8585 24084 8619
rect 24032 8576 24084 8585
rect 26516 8619 26568 8628
rect 26516 8585 26525 8619
rect 26525 8585 26559 8619
rect 26559 8585 26568 8619
rect 26516 8576 26568 8585
rect 27436 8619 27488 8628
rect 27436 8585 27445 8619
rect 27445 8585 27479 8619
rect 27479 8585 27488 8619
rect 27436 8576 27488 8585
rect 28172 8619 28224 8628
rect 28172 8585 28181 8619
rect 28181 8585 28215 8619
rect 28215 8585 28224 8619
rect 28172 8576 28224 8585
rect 28908 8619 28960 8628
rect 28908 8585 28917 8619
rect 28917 8585 28951 8619
rect 28951 8585 28960 8619
rect 28908 8576 28960 8585
rect 29828 8619 29880 8628
rect 29828 8585 29837 8619
rect 29837 8585 29871 8619
rect 29871 8585 29880 8619
rect 29828 8576 29880 8585
rect 31024 8619 31076 8628
rect 31024 8585 31033 8619
rect 31033 8585 31067 8619
rect 31067 8585 31076 8619
rect 31024 8576 31076 8585
rect 33140 8619 33192 8628
rect 33140 8585 33149 8619
rect 33149 8585 33183 8619
rect 33183 8585 33192 8619
rect 33140 8576 33192 8585
rect 53656 8576 53708 8628
rect 55864 8619 55916 8628
rect 55864 8585 55873 8619
rect 55873 8585 55907 8619
rect 55907 8585 55916 8619
rect 55864 8576 55916 8585
rect 56416 8576 56468 8628
rect 57336 8619 57388 8628
rect 57336 8585 57345 8619
rect 57345 8585 57379 8619
rect 57379 8585 57388 8619
rect 57336 8576 57388 8585
rect 58808 8619 58860 8628
rect 58808 8585 58817 8619
rect 58817 8585 58851 8619
rect 58851 8585 58860 8619
rect 58808 8576 58860 8585
rect 59268 8576 59320 8628
rect 60280 8619 60332 8628
rect 60280 8585 60289 8619
rect 60289 8585 60323 8619
rect 60323 8585 60332 8619
rect 60280 8576 60332 8585
rect 60648 8576 60700 8628
rect 62580 8619 62632 8628
rect 62580 8585 62589 8619
rect 62589 8585 62623 8619
rect 62623 8585 62632 8619
rect 62580 8576 62632 8585
rect 63960 8619 64012 8628
rect 63960 8585 63969 8619
rect 63969 8585 64003 8619
rect 64003 8585 64012 8619
rect 63960 8576 64012 8585
rect 64696 8619 64748 8628
rect 64696 8585 64705 8619
rect 64705 8585 64739 8619
rect 64739 8585 64748 8619
rect 64696 8576 64748 8585
rect 11060 8508 11112 8560
rect 20720 8508 20772 8560
rect 23388 8551 23440 8560
rect 23388 8517 23397 8551
rect 23397 8517 23431 8551
rect 23431 8517 23440 8551
rect 23388 8508 23440 8517
rect 22192 8483 22244 8492
rect 22192 8449 22201 8483
rect 22201 8449 22235 8483
rect 22235 8449 22244 8483
rect 25228 8508 25280 8560
rect 25688 8508 25740 8560
rect 27068 8508 27120 8560
rect 22192 8440 22244 8449
rect 22284 8372 22336 8424
rect 22652 8415 22704 8424
rect 22652 8381 22661 8415
rect 22661 8381 22695 8415
rect 22695 8381 22704 8415
rect 22652 8372 22704 8381
rect 18604 8304 18656 8356
rect 21088 8304 21140 8356
rect 23112 8372 23164 8424
rect 26148 8483 26200 8492
rect 24492 8372 24544 8424
rect 25688 8372 25740 8424
rect 26148 8449 26157 8483
rect 26157 8449 26191 8483
rect 26191 8449 26200 8483
rect 26148 8440 26200 8449
rect 27160 8440 27212 8492
rect 27252 8483 27304 8492
rect 27252 8449 27261 8483
rect 27261 8449 27295 8483
rect 27295 8449 27304 8483
rect 27252 8440 27304 8449
rect 27988 8483 28040 8492
rect 27988 8449 27997 8483
rect 27997 8449 28031 8483
rect 28031 8449 28040 8483
rect 27988 8440 28040 8449
rect 28724 8483 28776 8492
rect 28724 8449 28733 8483
rect 28733 8449 28767 8483
rect 28767 8449 28776 8483
rect 28724 8440 28776 8449
rect 29552 8483 29604 8492
rect 29552 8449 29561 8483
rect 29561 8449 29595 8483
rect 29595 8449 29604 8483
rect 29552 8440 29604 8449
rect 30840 8483 30892 8492
rect 30840 8449 30849 8483
rect 30849 8449 30883 8483
rect 30883 8449 30892 8483
rect 30840 8440 30892 8449
rect 32864 8483 32916 8492
rect 32864 8449 32873 8483
rect 32873 8449 32907 8483
rect 32907 8449 32916 8483
rect 32864 8440 32916 8449
rect 31944 8372 31996 8424
rect 33692 8483 33744 8492
rect 33692 8449 33701 8483
rect 33701 8449 33735 8483
rect 33735 8449 33744 8483
rect 33692 8440 33744 8449
rect 54668 8483 54720 8492
rect 54668 8449 54677 8483
rect 54677 8449 54711 8483
rect 54711 8449 54720 8483
rect 54668 8440 54720 8449
rect 55588 8483 55640 8492
rect 55588 8449 55597 8483
rect 55597 8449 55631 8483
rect 55631 8449 55640 8483
rect 55588 8440 55640 8449
rect 55680 8483 55732 8492
rect 55680 8449 55689 8483
rect 55689 8449 55723 8483
rect 55723 8449 55732 8483
rect 55680 8440 55732 8449
rect 57152 8483 57204 8492
rect 57152 8449 57161 8483
rect 57161 8449 57195 8483
rect 57195 8449 57204 8483
rect 57152 8440 57204 8449
rect 54392 8372 54444 8424
rect 56416 8372 56468 8424
rect 57336 8440 57388 8492
rect 65984 8508 66036 8560
rect 67088 8508 67140 8560
rect 87512 8576 87564 8628
rect 90824 8619 90876 8628
rect 90824 8585 90833 8619
rect 90833 8585 90867 8619
rect 90867 8585 90876 8619
rect 90824 8576 90876 8585
rect 91560 8576 91612 8628
rect 92572 8576 92624 8628
rect 94596 8619 94648 8628
rect 94596 8585 94605 8619
rect 94605 8585 94639 8619
rect 94639 8585 94648 8619
rect 94596 8576 94648 8585
rect 95056 8619 95108 8628
rect 95056 8585 95065 8619
rect 95065 8585 95099 8619
rect 95099 8585 95108 8619
rect 95056 8576 95108 8585
rect 95424 8619 95476 8628
rect 95424 8585 95433 8619
rect 95433 8585 95467 8619
rect 95467 8585 95476 8619
rect 95424 8576 95476 8585
rect 96160 8619 96212 8628
rect 96160 8585 96169 8619
rect 96169 8585 96203 8619
rect 96203 8585 96212 8619
rect 96160 8576 96212 8585
rect 96896 8619 96948 8628
rect 96896 8585 96905 8619
rect 96905 8585 96939 8619
rect 96939 8585 96948 8619
rect 96896 8576 96948 8585
rect 97264 8576 97316 8628
rect 58256 8440 58308 8492
rect 59360 8483 59412 8492
rect 59360 8449 59369 8483
rect 59369 8449 59403 8483
rect 59403 8449 59412 8483
rect 59360 8440 59412 8449
rect 60096 8483 60148 8492
rect 60096 8449 60105 8483
rect 60105 8449 60139 8483
rect 60139 8449 60148 8483
rect 60096 8440 60148 8449
rect 60832 8483 60884 8492
rect 60832 8449 60841 8483
rect 60841 8449 60875 8483
rect 60875 8449 60884 8483
rect 60832 8440 60884 8449
rect 62028 8440 62080 8492
rect 62488 8440 62540 8492
rect 63776 8483 63828 8492
rect 63776 8449 63785 8483
rect 63785 8449 63819 8483
rect 63819 8449 63828 8483
rect 63776 8440 63828 8449
rect 64512 8483 64564 8492
rect 64512 8449 64521 8483
rect 64521 8449 64555 8483
rect 64555 8449 64564 8483
rect 64512 8440 64564 8449
rect 65340 8483 65392 8492
rect 65340 8449 65349 8483
rect 65349 8449 65383 8483
rect 65383 8449 65392 8483
rect 65340 8440 65392 8449
rect 66076 8483 66128 8492
rect 66076 8449 66085 8483
rect 66085 8449 66119 8483
rect 66119 8449 66128 8483
rect 66076 8440 66128 8449
rect 89628 8508 89680 8560
rect 74264 8483 74316 8492
rect 74264 8449 74273 8483
rect 74273 8449 74307 8483
rect 74307 8449 74316 8483
rect 74264 8440 74316 8449
rect 74540 8483 74592 8492
rect 74540 8449 74549 8483
rect 74549 8449 74583 8483
rect 74583 8449 74592 8483
rect 74540 8440 74592 8449
rect 76472 8483 76524 8492
rect 76472 8449 76481 8483
rect 76481 8449 76515 8483
rect 76515 8449 76524 8483
rect 76472 8440 76524 8449
rect 88800 8483 88852 8492
rect 88800 8449 88809 8483
rect 88809 8449 88843 8483
rect 88843 8449 88852 8483
rect 88800 8440 88852 8449
rect 89996 8440 90048 8492
rect 90640 8483 90692 8492
rect 90640 8449 90649 8483
rect 90649 8449 90683 8483
rect 90683 8449 90692 8483
rect 90640 8440 90692 8449
rect 91008 8440 91060 8492
rect 93492 8440 93544 8492
rect 61292 8372 61344 8424
rect 61476 8372 61528 8424
rect 67364 8372 67416 8424
rect 82728 8372 82780 8424
rect 84844 8372 84896 8424
rect 92940 8372 92992 8424
rect 93032 8415 93084 8424
rect 93032 8381 93041 8415
rect 93041 8381 93075 8415
rect 93075 8381 93084 8415
rect 93032 8372 93084 8381
rect 23480 8304 23532 8356
rect 25044 8279 25096 8288
rect 25044 8245 25053 8279
rect 25053 8245 25087 8279
rect 25087 8245 25096 8279
rect 25044 8236 25096 8245
rect 28540 8304 28592 8356
rect 32956 8304 33008 8356
rect 54116 8304 54168 8356
rect 57336 8304 57388 8356
rect 57428 8304 57480 8356
rect 62672 8304 62724 8356
rect 65524 8347 65576 8356
rect 65524 8313 65533 8347
rect 65533 8313 65567 8347
rect 65567 8313 65576 8347
rect 65524 8304 65576 8313
rect 65892 8304 65944 8356
rect 97172 8508 97224 8560
rect 94412 8483 94464 8492
rect 94412 8449 94421 8483
rect 94421 8449 94455 8483
rect 94455 8449 94464 8483
rect 94412 8440 94464 8449
rect 94872 8483 94924 8492
rect 94872 8449 94881 8483
rect 94881 8449 94915 8483
rect 94915 8449 94924 8483
rect 94872 8440 94924 8449
rect 95056 8440 95108 8492
rect 95424 8440 95476 8492
rect 95700 8440 95752 8492
rect 95884 8440 95936 8492
rect 97264 8440 97316 8492
rect 97540 8619 97592 8628
rect 97540 8585 97549 8619
rect 97549 8585 97583 8619
rect 97583 8585 97592 8619
rect 97540 8576 97592 8585
rect 98000 8576 98052 8628
rect 99380 8576 99432 8628
rect 99472 8508 99524 8560
rect 121552 8576 121604 8628
rect 121644 8619 121696 8628
rect 121644 8585 121653 8619
rect 121653 8585 121687 8619
rect 121687 8585 121696 8619
rect 121644 8576 121696 8585
rect 122380 8619 122432 8628
rect 122380 8585 122389 8619
rect 122389 8585 122423 8619
rect 122423 8585 122432 8619
rect 122380 8576 122432 8585
rect 123208 8619 123260 8628
rect 123208 8585 123217 8619
rect 123217 8585 123251 8619
rect 123251 8585 123260 8619
rect 123208 8576 123260 8585
rect 124036 8619 124088 8628
rect 124036 8585 124045 8619
rect 124045 8585 124079 8619
rect 124079 8585 124088 8619
rect 124036 8576 124088 8585
rect 125600 8619 125652 8628
rect 125600 8585 125609 8619
rect 125609 8585 125643 8619
rect 125643 8585 125652 8619
rect 125600 8576 125652 8585
rect 126980 8619 127032 8628
rect 126980 8585 126989 8619
rect 126989 8585 127023 8619
rect 127023 8585 127032 8619
rect 126980 8576 127032 8585
rect 127716 8619 127768 8628
rect 127716 8585 127725 8619
rect 127725 8585 127759 8619
rect 127759 8585 127768 8619
rect 127716 8576 127768 8585
rect 128268 8619 128320 8628
rect 128268 8585 128277 8619
rect 128277 8585 128311 8619
rect 128311 8585 128320 8619
rect 128268 8576 128320 8585
rect 129372 8576 129424 8628
rect 132132 8619 132184 8628
rect 132132 8585 132141 8619
rect 132141 8585 132175 8619
rect 132175 8585 132184 8619
rect 132132 8576 132184 8585
rect 134524 8619 134576 8628
rect 134524 8585 134533 8619
rect 134533 8585 134567 8619
rect 134567 8585 134576 8619
rect 134524 8576 134576 8585
rect 137192 8576 137244 8628
rect 153844 8576 153896 8628
rect 156052 8576 156104 8628
rect 156236 8576 156288 8628
rect 161848 8576 161900 8628
rect 161940 8576 161992 8628
rect 100300 8508 100352 8560
rect 123392 8508 123444 8560
rect 127808 8508 127860 8560
rect 98092 8483 98144 8492
rect 98092 8449 98101 8483
rect 98101 8449 98135 8483
rect 98135 8449 98144 8483
rect 98092 8440 98144 8449
rect 99656 8483 99708 8492
rect 99656 8449 99665 8483
rect 99665 8449 99699 8483
rect 99699 8449 99708 8483
rect 99656 8440 99708 8449
rect 102048 8440 102100 8492
rect 96436 8372 96488 8424
rect 96620 8372 96672 8424
rect 98000 8372 98052 8424
rect 51172 8236 51224 8288
rect 61016 8279 61068 8288
rect 61016 8245 61025 8279
rect 61025 8245 61059 8279
rect 61059 8245 61068 8279
rect 61016 8236 61068 8245
rect 70400 8236 70452 8288
rect 90088 8279 90140 8288
rect 90088 8245 90097 8279
rect 90097 8245 90131 8279
rect 90131 8245 90140 8279
rect 90088 8236 90140 8245
rect 93216 8236 93268 8288
rect 95700 8304 95752 8356
rect 100760 8372 100812 8424
rect 100944 8415 100996 8424
rect 100944 8381 100953 8415
rect 100953 8381 100987 8415
rect 100987 8381 100996 8415
rect 100944 8372 100996 8381
rect 101956 8415 102008 8424
rect 101956 8381 101965 8415
rect 101965 8381 101999 8415
rect 101999 8381 102008 8415
rect 101956 8372 102008 8381
rect 120816 8372 120868 8424
rect 121828 8440 121880 8492
rect 122196 8483 122248 8492
rect 122196 8449 122205 8483
rect 122205 8449 122239 8483
rect 122239 8449 122248 8483
rect 122196 8440 122248 8449
rect 123024 8483 123076 8492
rect 123024 8449 123033 8483
rect 123033 8449 123067 8483
rect 123067 8449 123076 8483
rect 123024 8440 123076 8449
rect 123852 8483 123904 8492
rect 123852 8449 123861 8483
rect 123861 8449 123895 8483
rect 123895 8449 123904 8483
rect 123852 8440 123904 8449
rect 125416 8483 125468 8492
rect 125416 8449 125425 8483
rect 125425 8449 125459 8483
rect 125459 8449 125468 8483
rect 125416 8440 125468 8449
rect 126796 8483 126848 8492
rect 126796 8449 126805 8483
rect 126805 8449 126839 8483
rect 126839 8449 126848 8483
rect 126796 8440 126848 8449
rect 127532 8483 127584 8492
rect 127532 8449 127541 8483
rect 127541 8449 127575 8483
rect 127575 8449 127584 8483
rect 127532 8440 127584 8449
rect 128084 8483 128136 8492
rect 128084 8449 128093 8483
rect 128093 8449 128127 8483
rect 128127 8449 128136 8483
rect 128084 8440 128136 8449
rect 128820 8440 128872 8492
rect 131948 8483 132000 8492
rect 131948 8449 131957 8483
rect 131957 8449 131991 8483
rect 131991 8449 132000 8483
rect 131948 8440 132000 8449
rect 132868 8483 132920 8492
rect 132868 8449 132877 8483
rect 132877 8449 132911 8483
rect 132911 8449 132920 8483
rect 132868 8440 132920 8449
rect 134248 8483 134300 8492
rect 134248 8449 134257 8483
rect 134257 8449 134291 8483
rect 134291 8449 134300 8483
rect 134248 8440 134300 8449
rect 135536 8508 135588 8560
rect 143724 8508 143776 8560
rect 152464 8508 152516 8560
rect 154028 8508 154080 8560
rect 156512 8508 156564 8560
rect 153752 8440 153804 8492
rect 155960 8483 156012 8492
rect 155960 8449 155969 8483
rect 155969 8449 156003 8483
rect 156003 8449 156012 8483
rect 155960 8440 156012 8449
rect 171876 8508 171928 8560
rect 128912 8372 128964 8424
rect 113824 8304 113876 8356
rect 130200 8415 130252 8424
rect 130200 8381 130209 8415
rect 130209 8381 130243 8415
rect 130243 8381 130252 8415
rect 130844 8415 130896 8424
rect 130200 8372 130252 8381
rect 130844 8381 130853 8415
rect 130853 8381 130887 8415
rect 130887 8381 130896 8415
rect 130844 8372 130896 8381
rect 132684 8415 132736 8424
rect 132684 8381 132693 8415
rect 132693 8381 132727 8415
rect 132727 8381 132736 8415
rect 132684 8372 132736 8381
rect 142804 8372 142856 8424
rect 148784 8372 148836 8424
rect 156144 8372 156196 8424
rect 156236 8372 156288 8424
rect 157800 8415 157852 8424
rect 157800 8381 157809 8415
rect 157809 8381 157843 8415
rect 157843 8381 157852 8415
rect 157800 8372 157852 8381
rect 161296 8440 161348 8492
rect 162124 8483 162176 8492
rect 162124 8449 162133 8483
rect 162133 8449 162167 8483
rect 162167 8449 162176 8483
rect 162124 8440 162176 8449
rect 163872 8440 163924 8492
rect 165068 8483 165120 8492
rect 165068 8449 165077 8483
rect 165077 8449 165111 8483
rect 165111 8449 165120 8483
rect 165068 8440 165120 8449
rect 166356 8483 166408 8492
rect 166356 8449 166365 8483
rect 166365 8449 166399 8483
rect 166399 8449 166408 8483
rect 166356 8440 166408 8449
rect 166540 8440 166592 8492
rect 166816 8440 166868 8492
rect 166908 8440 166960 8492
rect 213920 8508 213972 8560
rect 186964 8483 187016 8492
rect 186964 8449 186973 8483
rect 186973 8449 187007 8483
rect 187007 8449 187016 8483
rect 186964 8440 187016 8449
rect 190368 8483 190420 8492
rect 190368 8449 190377 8483
rect 190377 8449 190411 8483
rect 190411 8449 190420 8483
rect 190368 8440 190420 8449
rect 191932 8440 191984 8492
rect 192392 8483 192444 8492
rect 192392 8449 192401 8483
rect 192401 8449 192435 8483
rect 192435 8449 192444 8483
rect 192392 8440 192444 8449
rect 192484 8483 192536 8492
rect 192484 8449 192493 8483
rect 192493 8449 192527 8483
rect 192527 8449 192536 8483
rect 192484 8440 192536 8449
rect 192668 8483 192720 8492
rect 192668 8449 192677 8483
rect 192677 8449 192711 8483
rect 192711 8449 192720 8483
rect 192668 8440 192720 8449
rect 193128 8483 193180 8492
rect 193128 8449 193137 8483
rect 193137 8449 193171 8483
rect 193171 8449 193180 8483
rect 193128 8440 193180 8449
rect 193864 8483 193916 8492
rect 193864 8449 193873 8483
rect 193873 8449 193907 8483
rect 193907 8449 193916 8483
rect 193864 8440 193916 8449
rect 159548 8372 159600 8424
rect 159916 8372 159968 8424
rect 161112 8372 161164 8424
rect 161664 8372 161716 8424
rect 162308 8372 162360 8424
rect 162676 8415 162728 8424
rect 162676 8381 162685 8415
rect 162685 8381 162719 8415
rect 162719 8381 162728 8415
rect 162676 8372 162728 8381
rect 163596 8372 163648 8424
rect 165344 8415 165396 8424
rect 111524 8236 111576 8288
rect 129096 8236 129148 8288
rect 132776 8236 132828 8288
rect 151452 8304 151504 8356
rect 154028 8304 154080 8356
rect 154672 8304 154724 8356
rect 165344 8381 165353 8415
rect 165353 8381 165387 8415
rect 165387 8381 165396 8415
rect 165344 8372 165396 8381
rect 168656 8415 168708 8424
rect 168656 8381 168665 8415
rect 168665 8381 168699 8415
rect 168699 8381 168708 8415
rect 168656 8372 168708 8381
rect 168932 8415 168984 8424
rect 168932 8381 168941 8415
rect 168941 8381 168975 8415
rect 168975 8381 168984 8415
rect 168932 8372 168984 8381
rect 169760 8372 169812 8424
rect 159272 8304 159324 8356
rect 161480 8304 161532 8356
rect 165068 8304 165120 8356
rect 151728 8236 151780 8288
rect 157064 8279 157116 8288
rect 157064 8245 157073 8279
rect 157073 8245 157107 8279
rect 157107 8245 157116 8279
rect 157064 8236 157116 8245
rect 160744 8236 160796 8288
rect 161940 8236 161992 8288
rect 164240 8236 164292 8288
rect 164700 8236 164752 8288
rect 166632 8279 166684 8288
rect 166632 8245 166641 8279
rect 166641 8245 166675 8279
rect 166675 8245 166684 8279
rect 166632 8236 166684 8245
rect 168840 8304 168892 8356
rect 169668 8304 169720 8356
rect 195612 8483 195664 8492
rect 195612 8449 195621 8483
rect 195621 8449 195655 8483
rect 195655 8449 195664 8483
rect 195612 8440 195664 8449
rect 196072 8483 196124 8492
rect 196072 8449 196081 8483
rect 196081 8449 196115 8483
rect 196115 8449 196124 8483
rect 196072 8440 196124 8449
rect 189908 8304 189960 8356
rect 191288 8347 191340 8356
rect 191288 8313 191297 8347
rect 191297 8313 191331 8347
rect 191331 8313 191340 8347
rect 191288 8304 191340 8313
rect 192852 8304 192904 8356
rect 194048 8347 194100 8356
rect 194048 8313 194057 8347
rect 194057 8313 194091 8347
rect 194091 8313 194100 8347
rect 194048 8304 194100 8313
rect 195980 8372 196032 8424
rect 197544 8483 197596 8492
rect 197544 8449 197553 8483
rect 197553 8449 197587 8483
rect 197587 8449 197596 8483
rect 197544 8440 197596 8449
rect 197728 8440 197780 8492
rect 198556 8483 198608 8492
rect 198556 8449 198565 8483
rect 198565 8449 198599 8483
rect 198599 8449 198608 8483
rect 198556 8440 198608 8449
rect 199200 8440 199252 8492
rect 200212 8440 200264 8492
rect 201040 8440 201092 8492
rect 201868 8440 201920 8492
rect 202512 8483 202564 8492
rect 202512 8449 202521 8483
rect 202521 8449 202555 8483
rect 202555 8449 202564 8483
rect 202512 8440 202564 8449
rect 202696 8483 202748 8492
rect 202696 8449 202705 8483
rect 202705 8449 202739 8483
rect 202739 8449 202748 8483
rect 202696 8440 202748 8449
rect 197084 8372 197136 8424
rect 198740 8372 198792 8424
rect 203524 8483 203576 8492
rect 203524 8449 203533 8483
rect 203533 8449 203567 8483
rect 203567 8449 203576 8483
rect 203524 8440 203576 8449
rect 195796 8304 195848 8356
rect 199108 8304 199160 8356
rect 199936 8347 199988 8356
rect 199936 8313 199945 8347
rect 199945 8313 199979 8347
rect 199979 8313 199988 8347
rect 199936 8304 199988 8313
rect 200764 8347 200816 8356
rect 200764 8313 200773 8347
rect 200773 8313 200807 8347
rect 200807 8313 200816 8347
rect 200764 8304 200816 8313
rect 200948 8304 201000 8356
rect 202972 8372 203024 8424
rect 203248 8304 203300 8356
rect 211804 8304 211856 8356
rect 216404 8576 216456 8628
rect 219440 8576 219492 8628
rect 220912 8576 220964 8628
rect 223488 8576 223540 8628
rect 224684 8619 224736 8628
rect 224684 8585 224693 8619
rect 224693 8585 224727 8619
rect 224727 8585 224736 8619
rect 224684 8576 224736 8585
rect 224960 8576 225012 8628
rect 215484 8508 215536 8560
rect 217968 8508 218020 8560
rect 219256 8508 219308 8560
rect 223212 8508 223264 8560
rect 224408 8508 224460 8560
rect 225512 8619 225564 8628
rect 225512 8585 225521 8619
rect 225521 8585 225555 8619
rect 225555 8585 225564 8619
rect 225512 8576 225564 8585
rect 226248 8619 226300 8628
rect 226248 8585 226257 8619
rect 226257 8585 226291 8619
rect 226291 8585 226300 8619
rect 226248 8576 226300 8585
rect 226984 8619 227036 8628
rect 226984 8585 226993 8619
rect 226993 8585 227027 8619
rect 227027 8585 227036 8619
rect 226984 8576 227036 8585
rect 228456 8619 228508 8628
rect 228456 8585 228465 8619
rect 228465 8585 228499 8619
rect 228499 8585 228508 8619
rect 228456 8576 228508 8585
rect 229192 8619 229244 8628
rect 229192 8585 229201 8619
rect 229201 8585 229235 8619
rect 229235 8585 229244 8619
rect 229192 8576 229244 8585
rect 230848 8576 230900 8628
rect 230940 8619 230992 8628
rect 230940 8585 230949 8619
rect 230949 8585 230983 8619
rect 230983 8585 230992 8619
rect 230940 8576 230992 8585
rect 231676 8619 231728 8628
rect 231676 8585 231685 8619
rect 231685 8585 231719 8619
rect 231719 8585 231728 8619
rect 231676 8576 231728 8585
rect 231768 8576 231820 8628
rect 232504 8576 232556 8628
rect 232596 8619 232648 8628
rect 232596 8585 232605 8619
rect 232605 8585 232639 8619
rect 232639 8585 232648 8619
rect 232596 8576 232648 8585
rect 234436 8619 234488 8628
rect 234436 8585 234445 8619
rect 234445 8585 234479 8619
rect 234479 8585 234488 8619
rect 234436 8576 234488 8585
rect 236276 8619 236328 8628
rect 236276 8585 236285 8619
rect 236285 8585 236319 8619
rect 236319 8585 236328 8619
rect 236276 8576 236328 8585
rect 215208 8440 215260 8492
rect 220452 8440 220504 8492
rect 221464 8440 221516 8492
rect 195980 8236 196032 8288
rect 196164 8236 196216 8288
rect 219164 8304 219216 8356
rect 221280 8372 221332 8424
rect 223764 8372 223816 8424
rect 224040 8440 224092 8492
rect 224224 8372 224276 8424
rect 224500 8483 224552 8492
rect 224500 8449 224509 8483
rect 224509 8449 224543 8483
rect 224543 8449 224552 8483
rect 224500 8440 224552 8449
rect 225328 8483 225380 8492
rect 225328 8449 225337 8483
rect 225337 8449 225371 8483
rect 225371 8449 225380 8483
rect 225328 8440 225380 8449
rect 226064 8483 226116 8492
rect 226064 8449 226073 8483
rect 226073 8449 226107 8483
rect 226107 8449 226116 8483
rect 226064 8440 226116 8449
rect 226800 8483 226852 8492
rect 226800 8449 226809 8483
rect 226809 8449 226843 8483
rect 226843 8449 226852 8483
rect 226800 8440 226852 8449
rect 227812 8440 227864 8492
rect 226248 8372 226300 8424
rect 228272 8483 228324 8492
rect 228272 8449 228281 8483
rect 228281 8449 228315 8483
rect 228315 8449 228324 8483
rect 228272 8440 228324 8449
rect 229008 8483 229060 8492
rect 229008 8449 229017 8483
rect 229017 8449 229051 8483
rect 229051 8449 229060 8483
rect 229008 8440 229060 8449
rect 230204 8508 230256 8560
rect 232320 8508 232372 8560
rect 248880 8576 248932 8628
rect 248972 8576 249024 8628
rect 251548 8576 251600 8628
rect 258264 8619 258316 8628
rect 258264 8585 258273 8619
rect 258273 8585 258307 8619
rect 258307 8585 258316 8619
rect 258264 8576 258316 8585
rect 259184 8619 259236 8628
rect 259184 8585 259193 8619
rect 259193 8585 259227 8619
rect 259227 8585 259236 8619
rect 259184 8576 259236 8585
rect 259920 8619 259972 8628
rect 259920 8585 259929 8619
rect 259929 8585 259963 8619
rect 259963 8585 259972 8619
rect 259920 8576 259972 8585
rect 260472 8619 260524 8628
rect 260472 8585 260481 8619
rect 260481 8585 260515 8619
rect 260515 8585 260524 8619
rect 260472 8576 260524 8585
rect 261852 8576 261904 8628
rect 262588 8576 262640 8628
rect 230112 8483 230164 8492
rect 230112 8449 230121 8483
rect 230121 8449 230155 8483
rect 230155 8449 230164 8483
rect 230112 8440 230164 8449
rect 231492 8483 231544 8492
rect 231492 8449 231501 8483
rect 231501 8449 231535 8483
rect 231535 8449 231544 8483
rect 231492 8440 231544 8449
rect 232412 8483 232464 8492
rect 232412 8449 232421 8483
rect 232421 8449 232455 8483
rect 232455 8449 232464 8483
rect 232412 8440 232464 8449
rect 239312 8508 239364 8560
rect 228916 8372 228968 8424
rect 229100 8372 229152 8424
rect 229652 8372 229704 8424
rect 233700 8440 233752 8492
rect 234436 8440 234488 8492
rect 224776 8304 224828 8356
rect 224868 8304 224920 8356
rect 228364 8304 228416 8356
rect 228456 8304 228508 8356
rect 233424 8415 233476 8424
rect 233424 8381 233433 8415
rect 233433 8381 233467 8415
rect 233467 8381 233476 8415
rect 233424 8372 233476 8381
rect 235816 8372 235868 8424
rect 236000 8372 236052 8424
rect 250260 8440 250312 8492
rect 256700 8483 256752 8492
rect 256700 8449 256709 8483
rect 256709 8449 256743 8483
rect 256743 8449 256752 8483
rect 256700 8440 256752 8449
rect 256976 8415 257028 8424
rect 256976 8381 256985 8415
rect 256985 8381 257019 8415
rect 257019 8381 257028 8415
rect 256976 8372 257028 8381
rect 258080 8483 258132 8492
rect 258080 8449 258089 8483
rect 258089 8449 258123 8483
rect 258123 8449 258132 8483
rect 258080 8440 258132 8449
rect 258264 8440 258316 8492
rect 263876 8508 263928 8560
rect 264244 8551 264296 8560
rect 264244 8517 264253 8551
rect 264253 8517 264287 8551
rect 264287 8517 264296 8551
rect 264244 8508 264296 8517
rect 264520 8508 264572 8560
rect 259736 8483 259788 8492
rect 259736 8449 259745 8483
rect 259745 8449 259779 8483
rect 259779 8449 259788 8483
rect 259736 8440 259788 8449
rect 260288 8483 260340 8492
rect 260288 8449 260297 8483
rect 260297 8449 260331 8483
rect 260331 8449 260340 8483
rect 260288 8440 260340 8449
rect 260380 8440 260432 8492
rect 230572 8304 230624 8356
rect 236460 8304 236512 8356
rect 260380 8304 260432 8356
rect 224592 8236 224644 8288
rect 224684 8236 224736 8288
rect 232504 8236 232556 8288
rect 232688 8236 232740 8288
rect 249064 8236 249116 8288
rect 251272 8236 251324 8288
rect 258724 8236 258776 8288
rect 261484 8440 261536 8492
rect 263048 8440 263100 8492
rect 265624 8576 265676 8628
rect 266268 8576 266320 8628
rect 265900 8508 265952 8560
rect 267096 8576 267148 8628
rect 268016 8508 268068 8560
rect 260932 8415 260984 8424
rect 260932 8381 260941 8415
rect 260941 8381 260975 8415
rect 260975 8381 260984 8415
rect 260932 8372 260984 8381
rect 261392 8372 261444 8424
rect 262404 8372 262456 8424
rect 265716 8483 265768 8492
rect 265716 8449 265725 8483
rect 265725 8449 265759 8483
rect 265759 8449 265768 8483
rect 265716 8440 265768 8449
rect 265808 8440 265860 8492
rect 263876 8304 263928 8356
rect 263968 8304 264020 8356
rect 264244 8304 264296 8356
rect 266544 8415 266596 8424
rect 266544 8381 266553 8415
rect 266553 8381 266587 8415
rect 266587 8381 266596 8415
rect 266544 8372 266596 8381
rect 266728 8483 266780 8492
rect 266728 8449 266737 8483
rect 266737 8449 266771 8483
rect 266771 8449 266780 8483
rect 266728 8440 266780 8449
rect 267280 8372 267332 8424
rect 267648 8483 267700 8492
rect 267648 8449 267657 8483
rect 267657 8449 267691 8483
rect 267691 8449 267700 8483
rect 267648 8440 267700 8449
rect 268384 8483 268436 8492
rect 268384 8449 268393 8483
rect 268393 8449 268427 8483
rect 268427 8449 268436 8483
rect 268384 8440 268436 8449
rect 268752 8440 268804 8492
rect 269764 8440 269816 8492
rect 270684 8483 270736 8492
rect 270684 8449 270693 8483
rect 270693 8449 270727 8483
rect 270727 8449 270736 8483
rect 270684 8440 270736 8449
rect 269304 8372 269356 8424
rect 262956 8236 263008 8288
rect 263232 8236 263284 8288
rect 264060 8236 264112 8288
rect 265164 8236 265216 8288
rect 268384 8236 268436 8288
rect 268476 8279 268528 8288
rect 268476 8245 268485 8279
rect 268485 8245 268519 8279
rect 268519 8245 268528 8279
rect 270500 8304 270552 8356
rect 268476 8236 268528 8245
rect 270040 8236 270092 8288
rect 34748 8134 34800 8186
rect 34812 8134 34864 8186
rect 34876 8134 34928 8186
rect 34940 8134 34992 8186
rect 35004 8134 35056 8186
rect 102345 8134 102397 8186
rect 102409 8134 102461 8186
rect 102473 8134 102525 8186
rect 102537 8134 102589 8186
rect 102601 8134 102653 8186
rect 169942 8134 169994 8186
rect 170006 8134 170058 8186
rect 170070 8134 170122 8186
rect 170134 8134 170186 8186
rect 170198 8134 170250 8186
rect 237539 8134 237591 8186
rect 237603 8134 237655 8186
rect 237667 8134 237719 8186
rect 237731 8134 237783 8186
rect 237795 8134 237847 8186
rect 9680 8032 9732 8084
rect 39212 8032 39264 8084
rect 66996 8032 67048 8084
rect 77576 8032 77628 8084
rect 84108 8032 84160 8084
rect 86684 8032 86736 8084
rect 100484 8032 100536 8084
rect 101036 8032 101088 8084
rect 21916 8007 21968 8016
rect 21916 7973 21925 8007
rect 21925 7973 21959 8007
rect 21959 7973 21968 8007
rect 21916 7964 21968 7973
rect 22928 8007 22980 8016
rect 22928 7973 22937 8007
rect 22937 7973 22971 8007
rect 22971 7973 22980 8007
rect 22928 7964 22980 7973
rect 23664 8007 23716 8016
rect 23664 7973 23673 8007
rect 23673 7973 23707 8007
rect 23707 7973 23716 8007
rect 23664 7964 23716 7973
rect 25228 8007 25280 8016
rect 25228 7973 25237 8007
rect 25237 7973 25271 8007
rect 25271 7973 25280 8007
rect 25228 7964 25280 7973
rect 25320 7964 25372 8016
rect 48964 7964 49016 8016
rect 75000 7964 75052 8016
rect 95148 7964 95200 8016
rect 100668 7964 100720 8016
rect 109592 8032 109644 8084
rect 101496 7964 101548 8016
rect 116860 8032 116912 8084
rect 129280 8075 129332 8084
rect 129280 8041 129289 8075
rect 129289 8041 129323 8075
rect 129323 8041 129332 8075
rect 129280 8032 129332 8041
rect 132960 8075 133012 8084
rect 132960 8041 132969 8075
rect 132969 8041 133003 8075
rect 133003 8041 133012 8075
rect 132960 8032 133012 8041
rect 148600 8032 148652 8084
rect 153568 8032 153620 8084
rect 157248 8075 157300 8084
rect 157248 8041 157257 8075
rect 157257 8041 157291 8075
rect 157291 8041 157300 8075
rect 157248 8032 157300 8041
rect 158720 8075 158772 8084
rect 158720 8041 158729 8075
rect 158729 8041 158763 8075
rect 158763 8041 158772 8075
rect 158720 8032 158772 8041
rect 159456 8032 159508 8084
rect 160928 8075 160980 8084
rect 160928 8041 160937 8075
rect 160937 8041 160971 8075
rect 160971 8041 160980 8075
rect 160928 8032 160980 8041
rect 161020 8032 161072 8084
rect 162400 8075 162452 8084
rect 162400 8041 162409 8075
rect 162409 8041 162443 8075
rect 162443 8041 162452 8075
rect 162400 8032 162452 8041
rect 163872 8075 163924 8084
rect 163872 8041 163881 8075
rect 163881 8041 163915 8075
rect 163915 8041 163924 8075
rect 163872 8032 163924 8041
rect 163964 8032 164016 8084
rect 165344 8032 165396 8084
rect 16488 7896 16540 7948
rect 21640 7828 21692 7880
rect 22744 7871 22796 7880
rect 22744 7837 22753 7871
rect 22753 7837 22787 7871
rect 22787 7837 22796 7871
rect 22744 7828 22796 7837
rect 23480 7871 23532 7880
rect 23480 7837 23489 7871
rect 23489 7837 23523 7871
rect 23523 7837 23532 7871
rect 23480 7828 23532 7837
rect 25044 7871 25096 7880
rect 25044 7837 25053 7871
rect 25053 7837 25087 7871
rect 25087 7837 25096 7871
rect 25044 7828 25096 7837
rect 32864 7939 32916 7948
rect 32864 7905 32873 7939
rect 32873 7905 32907 7939
rect 32907 7905 32916 7939
rect 32864 7896 32916 7905
rect 46112 7896 46164 7948
rect 73712 7896 73764 7948
rect 88524 7896 88576 7948
rect 92572 7896 92624 7948
rect 96620 7896 96672 7948
rect 101956 7896 102008 7948
rect 104440 7896 104492 7948
rect 33968 7828 34020 7880
rect 51724 7828 51776 7880
rect 67088 7871 67140 7880
rect 67088 7837 67097 7871
rect 67097 7837 67131 7871
rect 67131 7837 67140 7871
rect 67088 7828 67140 7837
rect 90088 7828 90140 7880
rect 18420 7760 18472 7812
rect 25320 7760 25372 7812
rect 19156 7692 19208 7744
rect 27620 7692 27672 7744
rect 33968 7692 34020 7744
rect 51632 7760 51684 7812
rect 83280 7760 83332 7812
rect 91928 7828 91980 7880
rect 99288 7828 99340 7880
rect 100944 7828 100996 7880
rect 107752 7828 107804 7880
rect 109316 7871 109368 7880
rect 109316 7837 109325 7871
rect 109325 7837 109359 7871
rect 109359 7837 109368 7871
rect 109316 7828 109368 7837
rect 109592 7828 109644 7880
rect 117872 7964 117924 8016
rect 156604 7964 156656 8016
rect 164700 7964 164752 8016
rect 112812 7896 112864 7948
rect 120908 7896 120960 7948
rect 134248 7939 134300 7948
rect 134248 7905 134257 7939
rect 134257 7905 134291 7939
rect 134291 7905 134300 7939
rect 134248 7896 134300 7905
rect 144000 7896 144052 7948
rect 161940 7896 161992 7948
rect 177672 8032 177724 8084
rect 197176 8032 197228 8084
rect 219072 8032 219124 8084
rect 221096 8032 221148 8084
rect 249800 8032 249852 8084
rect 259552 8075 259604 8084
rect 259552 8041 259561 8075
rect 259561 8041 259595 8075
rect 259595 8041 259604 8075
rect 259552 8032 259604 8041
rect 259736 8032 259788 8084
rect 261760 8075 261812 8084
rect 261760 8041 261769 8075
rect 261769 8041 261803 8075
rect 261803 8041 261812 8075
rect 261760 8032 261812 8041
rect 262496 8075 262548 8084
rect 262496 8041 262505 8075
rect 262505 8041 262539 8075
rect 262539 8041 262548 8075
rect 262496 8032 262548 8041
rect 263324 8075 263376 8084
rect 263324 8041 263333 8075
rect 263333 8041 263367 8075
rect 263367 8041 263376 8075
rect 263324 8032 263376 8041
rect 110052 7871 110104 7880
rect 110052 7837 110061 7871
rect 110061 7837 110095 7871
rect 110095 7837 110104 7871
rect 110052 7828 110104 7837
rect 115388 7828 115440 7880
rect 117504 7828 117556 7880
rect 129096 7871 129148 7880
rect 129096 7837 129105 7871
rect 129105 7837 129139 7871
rect 129139 7837 129148 7871
rect 129096 7828 129148 7837
rect 132776 7871 132828 7880
rect 132776 7837 132785 7871
rect 132785 7837 132819 7871
rect 132819 7837 132828 7871
rect 132776 7828 132828 7837
rect 146484 7828 146536 7880
rect 154580 7828 154632 7880
rect 157064 7871 157116 7880
rect 157064 7837 157073 7871
rect 157073 7837 157107 7871
rect 157107 7837 157116 7871
rect 157064 7828 157116 7837
rect 158536 7871 158588 7880
rect 158536 7837 158545 7871
rect 158545 7837 158579 7871
rect 158579 7837 158588 7871
rect 158536 7828 158588 7837
rect 159272 7871 159324 7880
rect 159272 7837 159281 7871
rect 159281 7837 159315 7871
rect 159315 7837 159324 7871
rect 159272 7828 159324 7837
rect 160008 7871 160060 7880
rect 160008 7837 160017 7871
rect 160017 7837 160051 7871
rect 160051 7837 160060 7871
rect 160008 7828 160060 7837
rect 160744 7871 160796 7880
rect 160744 7837 160753 7871
rect 160753 7837 160787 7871
rect 160787 7837 160796 7871
rect 160744 7828 160796 7837
rect 161480 7871 161532 7880
rect 161480 7837 161489 7871
rect 161489 7837 161523 7871
rect 161523 7837 161532 7871
rect 161480 7828 161532 7837
rect 104164 7760 104216 7812
rect 115296 7803 115348 7812
rect 115296 7769 115305 7803
rect 115305 7769 115339 7803
rect 115339 7769 115348 7803
rect 115296 7760 115348 7769
rect 115756 7760 115808 7812
rect 152004 7760 152056 7812
rect 162216 7871 162268 7880
rect 162216 7837 162225 7871
rect 162225 7837 162259 7871
rect 162259 7837 162268 7871
rect 162216 7828 162268 7837
rect 163688 7871 163740 7880
rect 163688 7837 163697 7871
rect 163697 7837 163731 7871
rect 163731 7837 163740 7871
rect 163688 7828 163740 7837
rect 164424 7871 164476 7880
rect 164424 7837 164433 7871
rect 164433 7837 164467 7871
rect 164467 7837 164476 7871
rect 164424 7828 164476 7837
rect 165160 7871 165212 7880
rect 165160 7837 165169 7871
rect 165169 7837 165203 7871
rect 165203 7837 165212 7871
rect 165160 7828 165212 7837
rect 165896 7871 165948 7880
rect 165896 7837 165905 7871
rect 165905 7837 165939 7871
rect 165939 7837 165948 7871
rect 165896 7828 165948 7837
rect 166632 7964 166684 8016
rect 169024 7964 169076 8016
rect 169208 8007 169260 8016
rect 169208 7973 169217 8007
rect 169217 7973 169251 8007
rect 169251 7973 169260 8007
rect 169208 7964 169260 7973
rect 169668 7964 169720 8016
rect 166816 7896 166868 7948
rect 167828 7871 167880 7880
rect 167828 7837 167837 7871
rect 167837 7837 167871 7871
rect 167871 7837 167880 7871
rect 167828 7828 167880 7837
rect 169760 7896 169812 7948
rect 171784 7964 171836 8016
rect 182088 7964 182140 8016
rect 198740 7964 198792 8016
rect 199384 7964 199436 8016
rect 211252 7964 211304 8016
rect 218980 7964 219032 8016
rect 226064 7964 226116 8016
rect 226340 7964 226392 8016
rect 256884 7964 256936 8016
rect 258724 7964 258776 8016
rect 263232 7964 263284 8016
rect 213552 7896 213604 7948
rect 223856 7896 223908 7948
rect 255320 7896 255372 7948
rect 264888 8032 264940 8084
rect 265256 8032 265308 8084
rect 266360 8032 266412 8084
rect 267004 7964 267056 8016
rect 268016 7964 268068 8016
rect 268844 8075 268896 8084
rect 268844 8041 268853 8075
rect 268853 8041 268887 8075
rect 268887 8041 268896 8075
rect 268844 8032 268896 8041
rect 269580 8032 269632 8084
rect 270040 8032 270092 8084
rect 271052 8032 271104 8084
rect 271144 8032 271196 8084
rect 272156 8032 272208 8084
rect 270316 7964 270368 8016
rect 168932 7828 168984 7880
rect 170588 7828 170640 7880
rect 172612 7828 172664 7880
rect 202972 7871 203024 7880
rect 202972 7837 202981 7871
rect 202981 7837 203015 7871
rect 203015 7837 203024 7871
rect 202972 7828 203024 7837
rect 211160 7828 211212 7880
rect 219256 7828 219308 7880
rect 224040 7828 224092 7880
rect 162124 7760 162176 7812
rect 210332 7760 210384 7812
rect 213828 7760 213880 7812
rect 89720 7735 89772 7744
rect 89720 7701 89729 7735
rect 89729 7701 89763 7735
rect 89763 7701 89772 7735
rect 89720 7692 89772 7701
rect 95976 7692 96028 7744
rect 98000 7692 98052 7744
rect 109040 7692 109092 7744
rect 109500 7692 109552 7744
rect 114928 7692 114980 7744
rect 115112 7735 115164 7744
rect 115112 7701 115121 7735
rect 115121 7701 115155 7735
rect 115155 7701 115164 7735
rect 115112 7692 115164 7701
rect 115204 7735 115256 7744
rect 115204 7701 115213 7735
rect 115213 7701 115247 7735
rect 115247 7701 115256 7735
rect 115204 7692 115256 7701
rect 115480 7735 115532 7744
rect 115480 7701 115489 7735
rect 115489 7701 115523 7735
rect 115523 7701 115532 7735
rect 115480 7692 115532 7701
rect 151820 7692 151872 7744
rect 158076 7692 158128 7744
rect 159364 7692 159416 7744
rect 165252 7692 165304 7744
rect 166540 7692 166592 7744
rect 169668 7692 169720 7744
rect 189724 7692 189776 7744
rect 210424 7692 210476 7744
rect 220820 7692 220872 7744
rect 223672 7760 223724 7812
rect 224776 7760 224828 7812
rect 225512 7871 225564 7880
rect 225512 7837 225521 7871
rect 225521 7837 225555 7871
rect 225555 7837 225564 7871
rect 225512 7828 225564 7837
rect 227352 7828 227404 7880
rect 234528 7828 234580 7880
rect 234712 7871 234764 7880
rect 234712 7837 234721 7871
rect 234721 7837 234755 7871
rect 234755 7837 234764 7871
rect 234712 7828 234764 7837
rect 234804 7828 234856 7880
rect 253112 7828 253164 7880
rect 234436 7760 234488 7812
rect 236644 7760 236696 7812
rect 256976 7760 257028 7812
rect 261576 7871 261628 7880
rect 261576 7837 261585 7871
rect 261585 7837 261619 7871
rect 261619 7837 261628 7871
rect 261576 7828 261628 7837
rect 262312 7871 262364 7880
rect 262312 7837 262321 7871
rect 262321 7837 262355 7871
rect 262355 7837 262364 7871
rect 262312 7828 262364 7837
rect 263140 7871 263192 7880
rect 263140 7837 263149 7871
rect 263149 7837 263183 7871
rect 263183 7837 263192 7871
rect 263140 7828 263192 7837
rect 263876 7828 263928 7880
rect 265624 7871 265676 7880
rect 265624 7837 265633 7871
rect 265633 7837 265667 7871
rect 265667 7837 265676 7871
rect 265624 7828 265676 7837
rect 267740 7896 267792 7948
rect 267556 7828 267608 7880
rect 264888 7760 264940 7812
rect 268200 7828 268252 7880
rect 268384 7828 268436 7880
rect 268476 7828 268528 7880
rect 268936 7828 268988 7880
rect 224960 7692 225012 7744
rect 225696 7735 225748 7744
rect 225696 7701 225705 7735
rect 225705 7701 225739 7735
rect 225739 7701 225748 7735
rect 225696 7692 225748 7701
rect 234528 7692 234580 7744
rect 234804 7692 234856 7744
rect 234896 7735 234948 7744
rect 234896 7701 234905 7735
rect 234905 7701 234939 7735
rect 234939 7701 234948 7735
rect 234896 7692 234948 7701
rect 235816 7735 235868 7744
rect 235816 7701 235825 7735
rect 235825 7701 235859 7735
rect 235859 7701 235868 7735
rect 235816 7692 235868 7701
rect 237196 7692 237248 7744
rect 240140 7692 240192 7744
rect 248880 7692 248932 7744
rect 249800 7692 249852 7744
rect 262220 7692 262272 7744
rect 262772 7692 262824 7744
rect 265992 7692 266044 7744
rect 268016 7692 268068 7744
rect 269212 7735 269264 7744
rect 269212 7701 269221 7735
rect 269221 7701 269255 7735
rect 269255 7701 269264 7735
rect 269212 7692 269264 7701
rect 269856 7871 269908 7880
rect 269856 7837 269865 7871
rect 269865 7837 269899 7871
rect 269899 7837 269908 7871
rect 269856 7828 269908 7837
rect 270132 7871 270184 7880
rect 270132 7837 270135 7871
rect 270135 7837 270184 7871
rect 270132 7828 270184 7837
rect 270224 7760 270276 7812
rect 270040 7692 270092 7744
rect 68546 7590 68598 7642
rect 68610 7590 68662 7642
rect 68674 7590 68726 7642
rect 68738 7590 68790 7642
rect 68802 7590 68854 7642
rect 136143 7590 136195 7642
rect 136207 7590 136259 7642
rect 136271 7590 136323 7642
rect 136335 7590 136387 7642
rect 136399 7590 136451 7642
rect 203740 7590 203792 7642
rect 203804 7590 203856 7642
rect 203868 7590 203920 7642
rect 203932 7590 203984 7642
rect 203996 7590 204048 7642
rect 271337 7590 271389 7642
rect 271401 7590 271453 7642
rect 271465 7590 271517 7642
rect 271529 7590 271581 7642
rect 271593 7590 271645 7642
rect 4068 7488 4120 7540
rect 24952 7488 25004 7540
rect 76380 7531 76432 7540
rect 76380 7497 76389 7531
rect 76389 7497 76423 7531
rect 76423 7497 76432 7531
rect 76380 7488 76432 7497
rect 88524 7488 88576 7540
rect 95700 7488 95752 7540
rect 95884 7488 95936 7540
rect 100576 7488 100628 7540
rect 100760 7488 100812 7540
rect 107844 7488 107896 7540
rect 111524 7531 111576 7540
rect 111524 7497 111533 7531
rect 111533 7497 111567 7531
rect 111567 7497 111576 7531
rect 111524 7488 111576 7497
rect 111616 7488 111668 7540
rect 113088 7488 113140 7540
rect 24400 7420 24452 7472
rect 42984 7420 43036 7472
rect 97264 7420 97316 7472
rect 99196 7420 99248 7472
rect 99288 7420 99340 7472
rect 104164 7420 104216 7472
rect 108856 7420 108908 7472
rect 115296 7531 115348 7540
rect 115296 7497 115305 7531
rect 115305 7497 115339 7531
rect 115339 7497 115348 7531
rect 115296 7488 115348 7497
rect 115388 7531 115440 7540
rect 115388 7497 115397 7531
rect 115397 7497 115431 7531
rect 115431 7497 115440 7531
rect 115388 7488 115440 7497
rect 117504 7531 117556 7540
rect 117504 7497 117513 7531
rect 117513 7497 117547 7531
rect 117547 7497 117556 7531
rect 117504 7488 117556 7497
rect 121000 7488 121052 7540
rect 76564 7395 76616 7404
rect 76564 7361 76573 7395
rect 76573 7361 76607 7395
rect 76607 7361 76616 7395
rect 76564 7352 76616 7361
rect 78772 7395 78824 7404
rect 78772 7361 78781 7395
rect 78781 7361 78815 7395
rect 78815 7361 78824 7395
rect 78772 7352 78824 7361
rect 84200 7352 84252 7404
rect 95884 7352 95936 7404
rect 97356 7395 97408 7404
rect 97356 7361 97365 7395
rect 97365 7361 97399 7395
rect 97399 7361 97408 7395
rect 97356 7352 97408 7361
rect 97540 7395 97592 7404
rect 97540 7361 97549 7395
rect 97549 7361 97583 7395
rect 97583 7361 97592 7395
rect 97540 7352 97592 7361
rect 93952 7284 94004 7336
rect 33692 7148 33744 7200
rect 93860 7216 93912 7268
rect 96160 7284 96212 7336
rect 96528 7284 96580 7336
rect 98552 7284 98604 7336
rect 98736 7352 98788 7404
rect 101404 7352 101456 7404
rect 101496 7395 101548 7404
rect 101496 7361 101505 7395
rect 101505 7361 101539 7395
rect 101539 7361 101548 7395
rect 101496 7352 101548 7361
rect 107108 7395 107160 7404
rect 107108 7361 107117 7395
rect 107117 7361 107151 7395
rect 107151 7361 107160 7395
rect 107108 7352 107160 7361
rect 99012 7284 99064 7336
rect 109040 7395 109092 7404
rect 109040 7361 109049 7395
rect 109049 7361 109083 7395
rect 109083 7361 109092 7395
rect 109040 7352 109092 7361
rect 110696 7352 110748 7404
rect 111248 7395 111300 7404
rect 111248 7361 111257 7395
rect 111257 7361 111291 7395
rect 111291 7361 111300 7395
rect 111248 7352 111300 7361
rect 111340 7352 111392 7404
rect 116584 7420 116636 7472
rect 118516 7420 118568 7472
rect 151544 7488 151596 7540
rect 152556 7488 152608 7540
rect 162124 7488 162176 7540
rect 162400 7488 162452 7540
rect 166908 7531 166960 7540
rect 166908 7497 166917 7531
rect 166917 7497 166951 7531
rect 166951 7497 166960 7531
rect 166908 7488 166960 7497
rect 112812 7395 112864 7404
rect 112812 7361 112821 7395
rect 112821 7361 112855 7395
rect 112855 7361 112864 7395
rect 112812 7352 112864 7361
rect 113088 7395 113140 7404
rect 113088 7361 113097 7395
rect 113097 7361 113131 7395
rect 113131 7361 113140 7395
rect 113088 7352 113140 7361
rect 115204 7352 115256 7404
rect 115572 7352 115624 7404
rect 116308 7395 116360 7404
rect 116308 7361 116317 7395
rect 116317 7361 116351 7395
rect 116351 7361 116360 7395
rect 116308 7352 116360 7361
rect 116768 7352 116820 7404
rect 118056 7395 118108 7404
rect 118056 7361 118065 7395
rect 118065 7361 118099 7395
rect 118099 7361 118108 7395
rect 118056 7352 118108 7361
rect 120080 7395 120132 7404
rect 120080 7361 120089 7395
rect 120089 7361 120123 7395
rect 120123 7361 120132 7395
rect 120080 7352 120132 7361
rect 124220 7352 124272 7404
rect 124772 7352 124824 7404
rect 154672 7420 154724 7472
rect 168656 7488 168708 7540
rect 179420 7488 179472 7540
rect 210424 7488 210476 7540
rect 221464 7531 221516 7540
rect 221464 7497 221473 7531
rect 221473 7497 221507 7531
rect 221507 7497 221516 7531
rect 221464 7488 221516 7497
rect 221924 7488 221976 7540
rect 224684 7488 224736 7540
rect 109132 7284 109184 7336
rect 99104 7216 99156 7268
rect 99472 7216 99524 7268
rect 109776 7216 109828 7268
rect 112536 7259 112588 7268
rect 112536 7225 112545 7259
rect 112545 7225 112579 7259
rect 112579 7225 112588 7259
rect 112536 7216 112588 7225
rect 115112 7284 115164 7336
rect 115480 7327 115532 7336
rect 115480 7293 115489 7327
rect 115489 7293 115523 7327
rect 115523 7293 115532 7327
rect 115480 7284 115532 7293
rect 117688 7284 117740 7336
rect 139216 7284 139268 7336
rect 151728 7352 151780 7404
rect 151820 7395 151872 7404
rect 151820 7361 151829 7395
rect 151829 7361 151863 7395
rect 151863 7361 151872 7395
rect 151820 7352 151872 7361
rect 152740 7395 152792 7404
rect 152740 7361 152749 7395
rect 152749 7361 152783 7395
rect 152783 7361 152792 7395
rect 152740 7352 152792 7361
rect 151636 7284 151688 7336
rect 97080 7148 97132 7200
rect 97448 7191 97500 7200
rect 97448 7157 97457 7191
rect 97457 7157 97491 7191
rect 97491 7157 97500 7191
rect 97448 7148 97500 7157
rect 97724 7191 97776 7200
rect 97724 7157 97733 7191
rect 97733 7157 97767 7191
rect 97767 7157 97776 7191
rect 97724 7148 97776 7157
rect 97816 7148 97868 7200
rect 99288 7191 99340 7200
rect 99288 7157 99297 7191
rect 99297 7157 99331 7191
rect 99331 7157 99340 7191
rect 99288 7148 99340 7157
rect 99932 7191 99984 7200
rect 99932 7157 99941 7191
rect 99941 7157 99975 7191
rect 99975 7157 99984 7191
rect 99932 7148 99984 7157
rect 100576 7148 100628 7200
rect 103428 7148 103480 7200
rect 103888 7148 103940 7200
rect 109224 7148 109276 7200
rect 111064 7191 111116 7200
rect 111064 7157 111073 7191
rect 111073 7157 111107 7191
rect 111107 7157 111116 7191
rect 111064 7148 111116 7157
rect 113272 7148 113324 7200
rect 113732 7191 113784 7200
rect 113732 7157 113741 7191
rect 113741 7157 113775 7191
rect 113775 7157 113784 7191
rect 113732 7148 113784 7157
rect 115664 7259 115716 7268
rect 115664 7225 115673 7259
rect 115673 7225 115707 7259
rect 115707 7225 115716 7259
rect 115664 7216 115716 7225
rect 118608 7216 118660 7268
rect 149336 7216 149388 7268
rect 160468 7352 160520 7404
rect 161296 7352 161348 7404
rect 162952 7395 163004 7404
rect 162952 7361 162961 7395
rect 162961 7361 162995 7395
rect 162995 7361 163004 7395
rect 162952 7352 163004 7361
rect 166724 7395 166776 7404
rect 166724 7361 166733 7395
rect 166733 7361 166767 7395
rect 166767 7361 166776 7395
rect 166724 7352 166776 7361
rect 169024 7352 169076 7404
rect 154672 7284 154724 7336
rect 171784 7284 171836 7336
rect 153660 7216 153712 7268
rect 210516 7420 210568 7472
rect 211436 7420 211488 7472
rect 219164 7420 219216 7472
rect 219256 7420 219308 7472
rect 223580 7420 223632 7472
rect 227352 7488 227404 7540
rect 227536 7488 227588 7540
rect 256792 7488 256844 7540
rect 213460 7395 213512 7404
rect 213460 7361 213469 7395
rect 213469 7361 213503 7395
rect 213503 7361 213512 7395
rect 213460 7352 213512 7361
rect 216864 7352 216916 7404
rect 225512 7420 225564 7472
rect 229744 7420 229796 7472
rect 249616 7420 249668 7472
rect 252100 7463 252152 7472
rect 252100 7429 252109 7463
rect 252109 7429 252143 7463
rect 252143 7429 252152 7463
rect 252100 7420 252152 7429
rect 213368 7284 213420 7336
rect 217968 7284 218020 7336
rect 224592 7395 224644 7404
rect 224592 7361 224601 7395
rect 224601 7361 224635 7395
rect 224635 7361 224644 7395
rect 224592 7352 224644 7361
rect 234436 7352 234488 7404
rect 236644 7352 236696 7404
rect 251456 7352 251508 7404
rect 252836 7395 252888 7404
rect 252836 7361 252845 7395
rect 252845 7361 252879 7395
rect 252879 7361 252888 7395
rect 252836 7352 252888 7361
rect 253112 7463 253164 7472
rect 253112 7429 253121 7463
rect 253121 7429 253155 7463
rect 253155 7429 253164 7463
rect 253112 7420 253164 7429
rect 262404 7488 262456 7540
rect 262772 7531 262824 7540
rect 262772 7497 262781 7531
rect 262781 7497 262815 7531
rect 262815 7497 262824 7531
rect 262772 7488 262824 7497
rect 263416 7531 263468 7540
rect 263416 7497 263425 7531
rect 263425 7497 263459 7531
rect 263459 7497 263468 7531
rect 263416 7488 263468 7497
rect 264336 7531 264388 7540
rect 264336 7497 264345 7531
rect 264345 7497 264379 7531
rect 264379 7497 264388 7531
rect 264336 7488 264388 7497
rect 265348 7488 265400 7540
rect 266176 7531 266228 7540
rect 266176 7497 266185 7531
rect 266185 7497 266219 7531
rect 266219 7497 266228 7531
rect 266176 7488 266228 7497
rect 253204 7352 253256 7404
rect 116400 7148 116452 7200
rect 116584 7191 116636 7200
rect 116584 7157 116593 7191
rect 116593 7157 116627 7191
rect 116627 7157 116636 7191
rect 116584 7148 116636 7157
rect 117136 7148 117188 7200
rect 118148 7191 118200 7200
rect 118148 7157 118157 7191
rect 118157 7157 118191 7191
rect 118191 7157 118200 7191
rect 118148 7148 118200 7157
rect 119436 7148 119488 7200
rect 146300 7148 146352 7200
rect 146392 7148 146444 7200
rect 151452 7148 151504 7200
rect 152188 7148 152240 7200
rect 172520 7148 172572 7200
rect 214288 7216 214340 7268
rect 210424 7148 210476 7200
rect 215300 7148 215352 7200
rect 219440 7216 219492 7268
rect 225052 7327 225104 7336
rect 225052 7293 225061 7327
rect 225061 7293 225095 7327
rect 225095 7293 225104 7327
rect 225052 7284 225104 7293
rect 249984 7327 250036 7336
rect 249984 7293 249993 7327
rect 249993 7293 250027 7327
rect 250027 7293 250036 7327
rect 249984 7284 250036 7293
rect 251180 7327 251232 7336
rect 251180 7293 251189 7327
rect 251189 7293 251223 7327
rect 251223 7293 251232 7327
rect 251180 7284 251232 7293
rect 261576 7352 261628 7404
rect 261668 7395 261720 7404
rect 261668 7361 261677 7395
rect 261677 7361 261711 7395
rect 261711 7361 261720 7395
rect 261668 7352 261720 7361
rect 262312 7395 262364 7404
rect 262312 7361 262321 7395
rect 262321 7361 262355 7395
rect 262355 7361 262364 7395
rect 262312 7352 262364 7361
rect 251640 7216 251692 7268
rect 267924 7420 267976 7472
rect 264060 7352 264112 7404
rect 264152 7395 264204 7404
rect 264152 7361 264161 7395
rect 264161 7361 264195 7395
rect 264195 7361 264204 7395
rect 264152 7352 264204 7361
rect 264336 7352 264388 7404
rect 264796 7352 264848 7404
rect 265256 7395 265308 7404
rect 265256 7361 265265 7395
rect 265265 7361 265299 7395
rect 265299 7361 265308 7395
rect 265256 7352 265308 7361
rect 265992 7395 266044 7404
rect 265992 7361 266007 7395
rect 266007 7361 266041 7395
rect 266041 7361 266044 7395
rect 265992 7352 266044 7361
rect 267280 7395 267332 7404
rect 267280 7361 267289 7395
rect 267289 7361 267323 7395
rect 267323 7361 267332 7395
rect 267280 7352 267332 7361
rect 267096 7327 267148 7336
rect 267096 7293 267105 7327
rect 267105 7293 267139 7327
rect 267139 7293 267148 7327
rect 267096 7284 267148 7293
rect 268200 7352 268252 7404
rect 268476 7488 268528 7540
rect 270316 7488 270368 7540
rect 270684 7488 270736 7540
rect 271144 7488 271196 7540
rect 272156 7488 272208 7540
rect 268844 7420 268896 7472
rect 269580 7395 269632 7404
rect 269580 7361 269611 7395
rect 269611 7361 269632 7395
rect 269580 7352 269632 7361
rect 270408 7420 270460 7472
rect 269764 7352 269816 7404
rect 223672 7148 223724 7200
rect 224592 7148 224644 7200
rect 226984 7148 227036 7200
rect 248420 7148 248472 7200
rect 252836 7148 252888 7200
rect 270776 7216 270828 7268
rect 266268 7148 266320 7200
rect 266912 7148 266964 7200
rect 267832 7148 267884 7200
rect 269120 7148 269172 7200
rect 34748 7046 34800 7098
rect 34812 7046 34864 7098
rect 34876 7046 34928 7098
rect 34940 7046 34992 7098
rect 35004 7046 35056 7098
rect 102345 7046 102397 7098
rect 102409 7046 102461 7098
rect 102473 7046 102525 7098
rect 102537 7046 102589 7098
rect 102601 7046 102653 7098
rect 169942 7046 169994 7098
rect 170006 7046 170058 7098
rect 170070 7046 170122 7098
rect 170134 7046 170186 7098
rect 170198 7046 170250 7098
rect 237539 7046 237591 7098
rect 237603 7046 237655 7098
rect 237667 7046 237719 7098
rect 237731 7046 237783 7098
rect 237795 7046 237847 7098
rect 93584 6944 93636 6996
rect 96528 6944 96580 6996
rect 95516 6876 95568 6928
rect 96160 6876 96212 6928
rect 19248 6808 19300 6860
rect 24768 6808 24820 6860
rect 30472 6808 30524 6860
rect 40868 6808 40920 6860
rect 95240 6808 95292 6860
rect 97172 6876 97224 6928
rect 98000 6944 98052 6996
rect 100944 6944 100996 6996
rect 106372 6944 106424 6996
rect 108396 6944 108448 6996
rect 108764 6987 108816 6996
rect 108764 6953 108773 6987
rect 108773 6953 108807 6987
rect 108807 6953 108816 6987
rect 108764 6944 108816 6953
rect 109040 6944 109092 6996
rect 110236 6944 110288 6996
rect 97908 6876 97960 6928
rect 96988 6808 97040 6860
rect 97540 6851 97592 6860
rect 97540 6817 97549 6851
rect 97549 6817 97583 6851
rect 97583 6817 97592 6851
rect 97540 6808 97592 6817
rect 24584 6740 24636 6792
rect 38844 6740 38896 6792
rect 39120 6740 39172 6792
rect 55864 6740 55916 6792
rect 20812 6672 20864 6724
rect 43996 6672 44048 6724
rect 46664 6672 46716 6724
rect 94504 6740 94556 6792
rect 96160 6783 96212 6792
rect 96160 6749 96169 6783
rect 96169 6749 96203 6783
rect 96203 6749 96212 6783
rect 96160 6740 96212 6749
rect 83188 6672 83240 6724
rect 93768 6672 93820 6724
rect 94688 6672 94740 6724
rect 97356 6740 97408 6792
rect 98276 6783 98328 6792
rect 98276 6749 98285 6783
rect 98285 6749 98319 6783
rect 98319 6749 98328 6783
rect 98276 6740 98328 6749
rect 98460 6783 98512 6792
rect 98460 6749 98469 6783
rect 98469 6749 98503 6783
rect 98503 6749 98512 6783
rect 98460 6740 98512 6749
rect 99196 6808 99248 6860
rect 100024 6808 100076 6860
rect 99380 6740 99432 6792
rect 99840 6783 99892 6792
rect 99840 6749 99849 6783
rect 99849 6749 99883 6783
rect 99883 6749 99892 6783
rect 99840 6740 99892 6749
rect 20720 6604 20772 6656
rect 45100 6604 45152 6656
rect 82820 6604 82872 6656
rect 94228 6604 94280 6656
rect 95976 6647 96028 6656
rect 95976 6613 95985 6647
rect 95985 6613 96019 6647
rect 96019 6613 96028 6647
rect 95976 6604 96028 6613
rect 96712 6647 96764 6656
rect 96712 6613 96721 6647
rect 96721 6613 96755 6647
rect 96755 6613 96764 6647
rect 96712 6604 96764 6613
rect 98092 6672 98144 6724
rect 98644 6647 98696 6656
rect 98644 6613 98653 6647
rect 98653 6613 98687 6647
rect 98687 6613 98696 6647
rect 98644 6604 98696 6613
rect 99656 6647 99708 6656
rect 99656 6613 99665 6647
rect 99665 6613 99699 6647
rect 99699 6613 99708 6647
rect 99656 6604 99708 6613
rect 99840 6604 99892 6656
rect 101220 6672 101272 6724
rect 101680 6740 101732 6792
rect 102232 6808 102284 6860
rect 107200 6876 107252 6928
rect 106280 6808 106332 6860
rect 110972 6876 111024 6928
rect 102324 6672 102376 6724
rect 102692 6783 102744 6792
rect 102692 6749 102701 6783
rect 102701 6749 102735 6783
rect 102735 6749 102744 6783
rect 102692 6740 102744 6749
rect 106188 6740 106240 6792
rect 107568 6740 107620 6792
rect 107016 6672 107068 6724
rect 110144 6808 110196 6860
rect 112536 6876 112588 6928
rect 113548 6876 113600 6928
rect 113732 6851 113784 6860
rect 113732 6817 113741 6851
rect 113741 6817 113775 6851
rect 113775 6817 113784 6851
rect 113732 6808 113784 6817
rect 114652 6876 114704 6928
rect 116584 6876 116636 6928
rect 116860 6876 116912 6928
rect 118608 6944 118660 6996
rect 144920 6944 144972 6996
rect 150900 6944 150952 6996
rect 151544 6944 151596 6996
rect 152096 6944 152148 6996
rect 114560 6851 114612 6860
rect 114560 6817 114569 6851
rect 114569 6817 114603 6851
rect 114603 6817 114612 6851
rect 114560 6808 114612 6817
rect 118148 6808 118200 6860
rect 145012 6876 145064 6928
rect 148968 6876 149020 6928
rect 150440 6876 150492 6928
rect 133236 6808 133288 6860
rect 151084 6808 151136 6860
rect 151820 6808 151872 6860
rect 152280 6808 152332 6860
rect 108580 6783 108632 6792
rect 108580 6749 108589 6783
rect 108589 6749 108623 6783
rect 108623 6749 108632 6783
rect 108580 6740 108632 6749
rect 108672 6783 108724 6792
rect 108672 6749 108681 6783
rect 108681 6749 108715 6783
rect 108715 6749 108724 6783
rect 108672 6740 108724 6749
rect 109960 6740 110012 6792
rect 110420 6783 110472 6792
rect 110420 6749 110429 6783
rect 110429 6749 110463 6783
rect 110463 6749 110472 6783
rect 110420 6740 110472 6749
rect 110972 6740 111024 6792
rect 112352 6783 112404 6792
rect 112352 6749 112361 6783
rect 112361 6749 112395 6783
rect 112395 6749 112404 6783
rect 112352 6740 112404 6749
rect 112996 6783 113048 6792
rect 112996 6749 113005 6783
rect 113005 6749 113039 6783
rect 113039 6749 113048 6783
rect 112996 6740 113048 6749
rect 115664 6740 115716 6792
rect 116216 6740 116268 6792
rect 109408 6672 109460 6724
rect 113088 6672 113140 6724
rect 113916 6715 113968 6724
rect 113916 6681 113925 6715
rect 113925 6681 113959 6715
rect 113959 6681 113968 6715
rect 113916 6672 113968 6681
rect 101128 6647 101180 6656
rect 101128 6613 101137 6647
rect 101137 6613 101171 6647
rect 101171 6613 101180 6647
rect 101128 6604 101180 6613
rect 101588 6604 101640 6656
rect 102140 6604 102192 6656
rect 103336 6604 103388 6656
rect 107476 6604 107528 6656
rect 107936 6647 107988 6656
rect 107936 6613 107945 6647
rect 107945 6613 107979 6647
rect 107979 6613 107988 6647
rect 107936 6604 107988 6613
rect 108028 6604 108080 6656
rect 109960 6604 110012 6656
rect 110972 6604 111024 6656
rect 111340 6604 111392 6656
rect 112536 6604 112588 6656
rect 112812 6647 112864 6656
rect 112812 6613 112821 6647
rect 112821 6613 112855 6647
rect 112855 6613 112864 6647
rect 112812 6604 112864 6613
rect 115112 6604 115164 6656
rect 115388 6604 115440 6656
rect 118424 6740 118476 6792
rect 150624 6740 150676 6792
rect 151544 6740 151596 6792
rect 152096 6740 152148 6792
rect 153384 6808 153436 6860
rect 153844 6808 153896 6860
rect 161296 6876 161348 6928
rect 161388 6876 161440 6928
rect 190184 6919 190236 6928
rect 190184 6885 190193 6919
rect 190193 6885 190227 6919
rect 190227 6885 190236 6919
rect 190184 6876 190236 6885
rect 213920 6944 213972 6996
rect 220820 6944 220872 6996
rect 221280 6944 221332 6996
rect 229744 6944 229796 6996
rect 249984 6944 250036 6996
rect 259736 6944 259788 6996
rect 261576 6944 261628 6996
rect 210424 6876 210476 6928
rect 210516 6876 210568 6928
rect 155040 6808 155092 6860
rect 157248 6808 157300 6860
rect 116860 6672 116912 6724
rect 117780 6672 117832 6724
rect 118148 6672 118200 6724
rect 142804 6672 142856 6724
rect 152464 6715 152516 6724
rect 152464 6681 152473 6715
rect 152473 6681 152507 6715
rect 152507 6681 152516 6715
rect 152464 6672 152516 6681
rect 153752 6740 153804 6792
rect 188804 6740 188856 6792
rect 189724 6740 189776 6792
rect 213184 6783 213236 6792
rect 213184 6749 213193 6783
rect 213193 6749 213227 6783
rect 213227 6749 213236 6783
rect 213184 6740 213236 6749
rect 213552 6740 213604 6792
rect 116676 6604 116728 6656
rect 117596 6604 117648 6656
rect 118056 6604 118108 6656
rect 119988 6604 120040 6656
rect 128084 6604 128136 6656
rect 140320 6604 140372 6656
rect 148968 6604 149020 6656
rect 151452 6604 151504 6656
rect 151728 6604 151780 6656
rect 153844 6672 153896 6724
rect 189356 6672 189408 6724
rect 189816 6672 189868 6724
rect 167736 6604 167788 6656
rect 168840 6604 168892 6656
rect 213644 6672 213696 6724
rect 210332 6604 210384 6656
rect 213920 6604 213972 6656
rect 216864 6851 216916 6860
rect 216864 6817 216873 6851
rect 216873 6817 216907 6851
rect 216907 6817 216916 6851
rect 216864 6808 216916 6817
rect 216128 6740 216180 6792
rect 217324 6783 217376 6792
rect 217324 6749 217333 6783
rect 217333 6749 217367 6783
rect 217367 6749 217376 6783
rect 217324 6740 217376 6749
rect 217876 6808 217928 6860
rect 218244 6808 218296 6860
rect 219624 6808 219676 6860
rect 224868 6876 224920 6928
rect 227628 6876 227680 6928
rect 236460 6876 236512 6928
rect 224316 6808 224368 6860
rect 226616 6808 226668 6860
rect 226984 6851 227036 6860
rect 226984 6817 226993 6851
rect 226993 6817 227027 6851
rect 227027 6817 227036 6851
rect 226984 6808 227036 6817
rect 219164 6740 219216 6792
rect 224224 6740 224276 6792
rect 224776 6740 224828 6792
rect 224960 6740 225012 6792
rect 241244 6808 241296 6860
rect 264612 6944 264664 6996
rect 267648 6944 267700 6996
rect 267740 6944 267792 6996
rect 270500 6944 270552 6996
rect 250076 6808 250128 6860
rect 251640 6808 251692 6860
rect 268292 6876 268344 6928
rect 216312 6715 216364 6724
rect 216312 6681 216321 6715
rect 216321 6681 216355 6715
rect 216355 6681 216364 6715
rect 216312 6672 216364 6681
rect 219256 6672 219308 6724
rect 224132 6715 224184 6724
rect 216496 6647 216548 6656
rect 216496 6613 216505 6647
rect 216505 6613 216539 6647
rect 216539 6613 216548 6647
rect 216496 6604 216548 6613
rect 217048 6604 217100 6656
rect 218704 6604 218756 6656
rect 224132 6681 224141 6715
rect 224141 6681 224175 6715
rect 224175 6681 224184 6715
rect 224132 6672 224184 6681
rect 219532 6604 219584 6656
rect 221096 6604 221148 6656
rect 223488 6604 223540 6656
rect 225788 6672 225840 6724
rect 233056 6672 233108 6724
rect 239036 6715 239088 6724
rect 239036 6681 239045 6715
rect 239045 6681 239079 6715
rect 239079 6681 239088 6715
rect 239036 6672 239088 6681
rect 241336 6740 241388 6792
rect 248420 6740 248472 6792
rect 248512 6740 248564 6792
rect 249340 6783 249392 6792
rect 249340 6749 249349 6783
rect 249349 6749 249383 6783
rect 249383 6749 249392 6783
rect 249340 6740 249392 6749
rect 251364 6783 251416 6792
rect 251364 6749 251373 6783
rect 251373 6749 251407 6783
rect 251407 6749 251416 6783
rect 251364 6740 251416 6749
rect 251456 6783 251508 6792
rect 251456 6749 251465 6783
rect 251465 6749 251499 6783
rect 251499 6749 251508 6783
rect 251456 6740 251508 6749
rect 253020 6783 253072 6792
rect 253020 6749 253029 6783
rect 253029 6749 253063 6783
rect 253063 6749 253072 6783
rect 253020 6740 253072 6749
rect 253204 6740 253256 6792
rect 256700 6740 256752 6792
rect 261944 6783 261996 6792
rect 261944 6749 261953 6783
rect 261953 6749 261987 6783
rect 261987 6749 261996 6783
rect 261944 6740 261996 6749
rect 263968 6808 264020 6860
rect 264060 6808 264112 6860
rect 267924 6808 267976 6860
rect 263232 6783 263284 6792
rect 263232 6749 263241 6783
rect 263241 6749 263275 6783
rect 263275 6749 263284 6783
rect 263232 6740 263284 6749
rect 263692 6783 263744 6792
rect 263692 6749 263701 6783
rect 263701 6749 263735 6783
rect 263735 6749 263744 6783
rect 263692 6740 263744 6749
rect 226156 6604 226208 6656
rect 226800 6604 226852 6656
rect 253112 6672 253164 6724
rect 248880 6604 248932 6656
rect 249248 6604 249300 6656
rect 251640 6647 251692 6656
rect 251640 6613 251649 6647
rect 251649 6613 251683 6647
rect 251683 6613 251692 6647
rect 251640 6604 251692 6613
rect 251732 6604 251784 6656
rect 260840 6672 260892 6724
rect 253848 6604 253900 6656
rect 255596 6604 255648 6656
rect 255780 6647 255832 6656
rect 255780 6613 255789 6647
rect 255789 6613 255823 6647
rect 255823 6613 255832 6647
rect 255780 6604 255832 6613
rect 256608 6604 256660 6656
rect 263048 6647 263100 6656
rect 263048 6613 263057 6647
rect 263057 6613 263091 6647
rect 263091 6613 263100 6647
rect 263048 6604 263100 6613
rect 263784 6647 263836 6656
rect 263784 6613 263793 6647
rect 263793 6613 263827 6647
rect 263827 6613 263836 6647
rect 263784 6604 263836 6613
rect 264888 6715 264940 6724
rect 264888 6681 264897 6715
rect 264897 6681 264931 6715
rect 264931 6681 264940 6715
rect 264888 6672 264940 6681
rect 265900 6783 265952 6792
rect 265900 6749 265909 6783
rect 265909 6749 265943 6783
rect 265943 6749 265952 6783
rect 265900 6740 265952 6749
rect 266820 6783 266872 6792
rect 266820 6749 266829 6783
rect 266829 6749 266863 6783
rect 266863 6749 266872 6783
rect 266820 6740 266872 6749
rect 267280 6740 267332 6792
rect 267556 6740 267608 6792
rect 267740 6672 267792 6724
rect 268016 6783 268068 6792
rect 268016 6749 268025 6783
rect 268025 6749 268059 6783
rect 268059 6749 268068 6783
rect 268016 6740 268068 6749
rect 268752 6808 268804 6860
rect 270224 6808 270276 6860
rect 269212 6783 269264 6792
rect 269212 6749 269221 6783
rect 269221 6749 269255 6783
rect 269255 6749 269264 6783
rect 269212 6740 269264 6749
rect 269856 6783 269908 6792
rect 269856 6749 269865 6783
rect 269865 6749 269899 6783
rect 269899 6749 269908 6783
rect 269856 6740 269908 6749
rect 270040 6783 270092 6792
rect 270040 6749 270049 6783
rect 270049 6749 270083 6783
rect 270083 6749 270092 6783
rect 270040 6740 270092 6749
rect 265992 6604 266044 6656
rect 266360 6604 266412 6656
rect 266636 6604 266688 6656
rect 267648 6604 267700 6656
rect 270132 6604 270184 6656
rect 68546 6502 68598 6554
rect 68610 6502 68662 6554
rect 68674 6502 68726 6554
rect 68738 6502 68790 6554
rect 68802 6502 68854 6554
rect 136143 6502 136195 6554
rect 136207 6502 136259 6554
rect 136271 6502 136323 6554
rect 136335 6502 136387 6554
rect 136399 6502 136451 6554
rect 203740 6502 203792 6554
rect 203804 6502 203856 6554
rect 203868 6502 203920 6554
rect 203932 6502 203984 6554
rect 203996 6502 204048 6554
rect 271337 6502 271389 6554
rect 271401 6502 271453 6554
rect 271465 6502 271517 6554
rect 271529 6502 271581 6554
rect 271593 6502 271645 6554
rect 12900 6400 12952 6452
rect 42708 6400 42760 6452
rect 72332 6400 72384 6452
rect 93952 6400 94004 6452
rect 95332 6400 95384 6452
rect 97724 6400 97776 6452
rect 98368 6400 98420 6452
rect 98736 6443 98788 6452
rect 98736 6409 98745 6443
rect 98745 6409 98779 6443
rect 98779 6409 98788 6443
rect 98736 6400 98788 6409
rect 8484 6332 8536 6384
rect 38752 6332 38804 6384
rect 15568 6264 15620 6316
rect 49516 6264 49568 6316
rect 13636 6196 13688 6248
rect 47492 6196 47544 6248
rect 13728 6128 13780 6180
rect 48872 6196 48924 6248
rect 48044 6128 48096 6180
rect 55772 6332 55824 6384
rect 96712 6332 96764 6384
rect 96804 6332 96856 6384
rect 98552 6332 98604 6384
rect 101036 6400 101088 6452
rect 101864 6400 101916 6452
rect 102324 6443 102376 6452
rect 102324 6409 102333 6443
rect 102333 6409 102367 6443
rect 102367 6409 102376 6443
rect 102324 6400 102376 6409
rect 108028 6400 108080 6452
rect 109316 6400 109368 6452
rect 51448 6264 51500 6316
rect 52368 6264 52420 6316
rect 80244 6264 80296 6316
rect 92940 6307 92992 6316
rect 92940 6273 92949 6307
rect 92949 6273 92983 6307
rect 92983 6273 92992 6307
rect 92940 6264 92992 6273
rect 95240 6264 95292 6316
rect 97908 6307 97960 6316
rect 97908 6273 97917 6307
rect 97917 6273 97951 6307
rect 97951 6273 97960 6307
rect 97908 6264 97960 6273
rect 98276 6264 98328 6316
rect 106004 6332 106056 6384
rect 110420 6400 110472 6452
rect 113916 6400 113968 6452
rect 115204 6400 115256 6452
rect 115480 6400 115532 6452
rect 116860 6400 116912 6452
rect 117872 6400 117924 6452
rect 118056 6400 118108 6452
rect 118148 6443 118200 6452
rect 118148 6409 118157 6443
rect 118157 6409 118191 6443
rect 118191 6409 118200 6443
rect 118148 6400 118200 6409
rect 118240 6400 118292 6452
rect 120080 6400 120132 6452
rect 130384 6400 130436 6452
rect 148140 6400 148192 6452
rect 149060 6400 149112 6452
rect 150256 6400 150308 6452
rect 150992 6400 151044 6452
rect 151268 6400 151320 6452
rect 151452 6400 151504 6452
rect 152372 6400 152424 6452
rect 153568 6400 153620 6452
rect 156328 6400 156380 6452
rect 159456 6400 159508 6452
rect 184848 6400 184900 6452
rect 188804 6443 188856 6452
rect 188804 6409 188813 6443
rect 188813 6409 188847 6443
rect 188847 6409 188856 6443
rect 188804 6400 188856 6409
rect 99564 6264 99616 6316
rect 100392 6264 100444 6316
rect 100668 6307 100720 6316
rect 100668 6273 100677 6307
rect 100677 6273 100711 6307
rect 100711 6273 100720 6307
rect 100668 6264 100720 6273
rect 101036 6264 101088 6316
rect 101496 6264 101548 6316
rect 101864 6264 101916 6316
rect 102048 6307 102100 6316
rect 102048 6273 102057 6307
rect 102057 6273 102091 6307
rect 102091 6273 102100 6307
rect 102048 6264 102100 6273
rect 104624 6307 104676 6316
rect 104624 6273 104633 6307
rect 104633 6273 104667 6307
rect 104667 6273 104676 6307
rect 104624 6264 104676 6273
rect 105636 6307 105688 6316
rect 105636 6273 105645 6307
rect 105645 6273 105679 6307
rect 105679 6273 105688 6307
rect 105636 6264 105688 6273
rect 106464 6264 106516 6316
rect 53104 6239 53156 6248
rect 53104 6205 53113 6239
rect 53113 6205 53147 6239
rect 53147 6205 53156 6239
rect 53104 6196 53156 6205
rect 91100 6196 91152 6248
rect 92664 6239 92716 6248
rect 92664 6205 92673 6239
rect 92673 6205 92707 6239
rect 92707 6205 92716 6239
rect 92664 6196 92716 6205
rect 53748 6171 53800 6180
rect 53748 6137 53757 6171
rect 53757 6137 53791 6171
rect 53791 6137 53800 6171
rect 53748 6128 53800 6137
rect 96896 6239 96948 6248
rect 96896 6205 96905 6239
rect 96905 6205 96939 6239
rect 96939 6205 96948 6239
rect 96896 6196 96948 6205
rect 97356 6196 97408 6248
rect 98460 6239 98512 6248
rect 98460 6205 98469 6239
rect 98469 6205 98503 6239
rect 98503 6205 98512 6239
rect 98460 6196 98512 6205
rect 99380 6196 99432 6248
rect 109776 6375 109828 6384
rect 109776 6341 109785 6375
rect 109785 6341 109819 6375
rect 109819 6341 109828 6375
rect 109776 6332 109828 6341
rect 113272 6332 113324 6384
rect 113548 6332 113600 6384
rect 108580 6307 108632 6316
rect 108580 6273 108589 6307
rect 108589 6273 108623 6307
rect 108623 6273 108632 6307
rect 108580 6264 108632 6273
rect 109592 6307 109644 6316
rect 109592 6273 109601 6307
rect 109601 6273 109635 6307
rect 109635 6273 109644 6307
rect 109592 6264 109644 6273
rect 18696 6060 18748 6112
rect 51540 6060 51592 6112
rect 92204 6060 92256 6112
rect 93860 6060 93912 6112
rect 94136 6060 94188 6112
rect 94780 6060 94832 6112
rect 96068 6060 96120 6112
rect 97448 6060 97500 6112
rect 97724 6103 97776 6112
rect 97724 6069 97733 6103
rect 97733 6069 97767 6103
rect 97767 6069 97776 6103
rect 97724 6060 97776 6069
rect 98000 6060 98052 6112
rect 99472 6060 99524 6112
rect 99748 6060 99800 6112
rect 100944 6060 100996 6112
rect 101680 6128 101732 6180
rect 104532 6128 104584 6180
rect 108672 6239 108724 6248
rect 108672 6205 108681 6239
rect 108681 6205 108715 6239
rect 108715 6205 108724 6239
rect 108672 6196 108724 6205
rect 109316 6196 109368 6248
rect 113456 6307 113508 6316
rect 113456 6273 113465 6307
rect 113465 6273 113499 6307
rect 113499 6273 113508 6307
rect 113456 6264 113508 6273
rect 113732 6307 113784 6316
rect 113732 6273 113741 6307
rect 113741 6273 113775 6307
rect 113775 6273 113784 6307
rect 113732 6264 113784 6273
rect 115020 6307 115072 6316
rect 115020 6273 115029 6307
rect 115029 6273 115063 6307
rect 115063 6273 115072 6307
rect 115020 6264 115072 6273
rect 115940 6307 115992 6316
rect 115940 6273 115949 6307
rect 115949 6273 115983 6307
rect 115983 6273 115992 6307
rect 115940 6264 115992 6273
rect 107384 6128 107436 6180
rect 108212 6128 108264 6180
rect 113456 6128 113508 6180
rect 115020 6128 115072 6180
rect 101864 6060 101916 6112
rect 103520 6060 103572 6112
rect 103796 6060 103848 6112
rect 105912 6060 105964 6112
rect 108764 6103 108816 6112
rect 108764 6069 108773 6103
rect 108773 6069 108807 6103
rect 108807 6069 108816 6103
rect 108764 6060 108816 6069
rect 108948 6103 109000 6112
rect 108948 6069 108957 6103
rect 108957 6069 108991 6103
rect 108991 6069 109000 6103
rect 108948 6060 109000 6069
rect 112260 6060 112312 6112
rect 112720 6060 112772 6112
rect 114652 6060 114704 6112
rect 116124 6196 116176 6248
rect 116400 6196 116452 6248
rect 116584 6196 116636 6248
rect 116860 6196 116912 6248
rect 117872 6239 117924 6248
rect 117872 6205 117881 6239
rect 117881 6205 117915 6239
rect 117915 6205 117924 6239
rect 117872 6196 117924 6205
rect 118424 6196 118476 6248
rect 118700 6196 118752 6248
rect 116216 6060 116268 6112
rect 116400 6060 116452 6112
rect 117320 6060 117372 6112
rect 118148 6060 118200 6112
rect 118884 6307 118936 6316
rect 118884 6273 118893 6307
rect 118893 6273 118927 6307
rect 118927 6273 118936 6307
rect 132868 6332 132920 6384
rect 162124 6332 162176 6384
rect 168012 6332 168064 6384
rect 189356 6443 189408 6452
rect 189356 6409 189365 6443
rect 189365 6409 189399 6443
rect 189399 6409 189408 6443
rect 189356 6400 189408 6409
rect 189448 6443 189500 6452
rect 189448 6409 189457 6443
rect 189457 6409 189491 6443
rect 189491 6409 189500 6443
rect 189448 6400 189500 6409
rect 189724 6443 189776 6452
rect 189724 6409 189733 6443
rect 189733 6409 189767 6443
rect 189767 6409 189776 6443
rect 189724 6400 189776 6409
rect 189816 6400 189868 6452
rect 216496 6400 216548 6452
rect 216588 6400 216640 6452
rect 222200 6400 222252 6452
rect 226156 6400 226208 6452
rect 226248 6400 226300 6452
rect 248328 6400 248380 6452
rect 249340 6443 249392 6452
rect 249340 6409 249349 6443
rect 249349 6409 249383 6443
rect 249383 6409 249392 6443
rect 249340 6400 249392 6409
rect 253112 6443 253164 6452
rect 253112 6409 253121 6443
rect 253121 6409 253155 6443
rect 253155 6409 253164 6443
rect 253112 6400 253164 6409
rect 255320 6400 255372 6452
rect 255596 6400 255648 6452
rect 256700 6443 256752 6452
rect 256700 6409 256709 6443
rect 256709 6409 256743 6443
rect 256743 6409 256752 6443
rect 256700 6400 256752 6409
rect 261944 6400 261996 6452
rect 264796 6400 264848 6452
rect 266820 6400 266872 6452
rect 269120 6400 269172 6452
rect 190000 6375 190052 6384
rect 190000 6341 190009 6375
rect 190009 6341 190043 6375
rect 190043 6341 190052 6375
rect 190000 6332 190052 6341
rect 216036 6332 216088 6384
rect 217324 6332 217376 6384
rect 221556 6332 221608 6384
rect 224408 6332 224460 6384
rect 231400 6332 231452 6384
rect 245108 6332 245160 6384
rect 118884 6264 118936 6273
rect 119068 6196 119120 6248
rect 130384 6196 130436 6248
rect 135536 6239 135588 6248
rect 135536 6205 135545 6239
rect 135545 6205 135579 6239
rect 135579 6205 135588 6239
rect 135536 6196 135588 6205
rect 137008 6307 137060 6316
rect 137008 6273 137017 6307
rect 137017 6273 137051 6307
rect 137051 6273 137060 6307
rect 137008 6264 137060 6273
rect 138664 6264 138716 6316
rect 140044 6264 140096 6316
rect 137192 6239 137244 6248
rect 137192 6205 137201 6239
rect 137201 6205 137235 6239
rect 137235 6205 137244 6239
rect 137192 6196 137244 6205
rect 139584 6196 139636 6248
rect 150164 6196 150216 6248
rect 120540 6128 120592 6180
rect 119896 6060 119948 6112
rect 142804 6128 142856 6180
rect 150624 6264 150676 6316
rect 150992 6196 151044 6248
rect 151544 6196 151596 6248
rect 152556 6264 152608 6316
rect 153752 6264 153804 6316
rect 152280 6196 152332 6248
rect 154856 6307 154908 6316
rect 154856 6273 154865 6307
rect 154865 6273 154899 6307
rect 154899 6273 154908 6307
rect 154856 6264 154908 6273
rect 156144 6307 156196 6316
rect 156144 6273 156153 6307
rect 156153 6273 156187 6307
rect 156187 6273 156196 6307
rect 156144 6264 156196 6273
rect 154948 6196 155000 6248
rect 155868 6196 155920 6248
rect 161204 6264 161256 6316
rect 161296 6264 161348 6316
rect 156328 6196 156380 6248
rect 161664 6196 161716 6248
rect 162860 6196 162912 6248
rect 165712 6196 165764 6248
rect 168656 6239 168708 6248
rect 168656 6205 168665 6239
rect 168665 6205 168699 6239
rect 168699 6205 168708 6239
rect 168656 6196 168708 6205
rect 153752 6128 153804 6180
rect 137008 6060 137060 6112
rect 139952 6060 140004 6112
rect 142252 6060 142304 6112
rect 143172 6060 143224 6112
rect 149060 6060 149112 6112
rect 150072 6103 150124 6112
rect 150072 6069 150081 6103
rect 150081 6069 150115 6103
rect 150115 6069 150124 6103
rect 150072 6060 150124 6069
rect 150900 6103 150952 6112
rect 150900 6069 150909 6103
rect 150909 6069 150943 6103
rect 150943 6069 150952 6103
rect 150900 6060 150952 6069
rect 152740 6060 152792 6112
rect 155776 6060 155828 6112
rect 158444 6128 158496 6180
rect 167736 6171 167788 6180
rect 167736 6137 167745 6171
rect 167745 6137 167779 6171
rect 167779 6137 167788 6171
rect 167736 6128 167788 6137
rect 169024 6171 169076 6180
rect 169024 6137 169033 6171
rect 169033 6137 169067 6171
rect 169067 6137 169076 6171
rect 169024 6128 169076 6137
rect 156328 6060 156380 6112
rect 156420 6060 156472 6112
rect 156788 6060 156840 6112
rect 159824 6060 159876 6112
rect 169760 6264 169812 6316
rect 171232 6264 171284 6316
rect 189540 6307 189592 6316
rect 189540 6273 189549 6307
rect 189549 6273 189583 6307
rect 189583 6273 189592 6307
rect 189540 6264 189592 6273
rect 207480 6264 207532 6316
rect 209136 6307 209188 6316
rect 209136 6273 209145 6307
rect 209145 6273 209179 6307
rect 209179 6273 209188 6307
rect 209136 6264 209188 6273
rect 209320 6264 209372 6316
rect 213092 6307 213144 6316
rect 213092 6273 213101 6307
rect 213101 6273 213135 6307
rect 213135 6273 213144 6307
rect 213092 6264 213144 6273
rect 216312 6264 216364 6316
rect 217876 6307 217928 6316
rect 217876 6273 217885 6307
rect 217885 6273 217919 6307
rect 217919 6273 217928 6307
rect 217876 6264 217928 6273
rect 185492 6128 185544 6180
rect 208492 6196 208544 6248
rect 209412 6239 209464 6248
rect 209412 6205 209421 6239
rect 209421 6205 209455 6239
rect 209455 6205 209464 6239
rect 209412 6196 209464 6205
rect 207756 6128 207808 6180
rect 212816 6196 212868 6248
rect 213460 6128 213512 6180
rect 200764 6060 200816 6112
rect 207296 6060 207348 6112
rect 215852 6103 215904 6112
rect 215852 6069 215861 6103
rect 215861 6069 215895 6103
rect 215895 6069 215904 6103
rect 217048 6196 217100 6248
rect 218060 6307 218112 6316
rect 218060 6273 218069 6307
rect 218069 6273 218103 6307
rect 218103 6273 218112 6307
rect 218060 6264 218112 6273
rect 218428 6264 218480 6316
rect 221372 6264 221424 6316
rect 221740 6307 221792 6316
rect 221740 6273 221749 6307
rect 221749 6273 221783 6307
rect 221783 6273 221792 6307
rect 221740 6264 221792 6273
rect 221832 6307 221884 6316
rect 221832 6273 221841 6307
rect 221841 6273 221875 6307
rect 221875 6273 221884 6307
rect 221832 6264 221884 6273
rect 224592 6307 224644 6316
rect 224592 6273 224601 6307
rect 224601 6273 224635 6307
rect 224635 6273 224644 6307
rect 224592 6264 224644 6273
rect 226156 6307 226208 6316
rect 226156 6273 226165 6307
rect 226165 6273 226199 6307
rect 226199 6273 226208 6307
rect 226156 6264 226208 6273
rect 226432 6307 226484 6316
rect 226432 6273 226441 6307
rect 226441 6273 226475 6307
rect 226475 6273 226484 6307
rect 226432 6264 226484 6273
rect 244648 6264 244700 6316
rect 248236 6264 248288 6316
rect 248328 6264 248380 6316
rect 218336 6196 218388 6248
rect 218980 6239 219032 6248
rect 218980 6205 218989 6239
rect 218989 6205 219023 6239
rect 219023 6205 219032 6239
rect 218980 6196 219032 6205
rect 219532 6196 219584 6248
rect 219900 6196 219952 6248
rect 220728 6196 220780 6248
rect 222292 6196 222344 6248
rect 222752 6239 222804 6248
rect 222752 6205 222761 6239
rect 222761 6205 222795 6239
rect 222795 6205 222804 6239
rect 222752 6196 222804 6205
rect 223304 6196 223356 6248
rect 225236 6239 225288 6248
rect 225236 6205 225245 6239
rect 225245 6205 225279 6239
rect 225279 6205 225288 6239
rect 225236 6196 225288 6205
rect 225420 6239 225472 6248
rect 225420 6205 225429 6239
rect 225429 6205 225463 6239
rect 225463 6205 225472 6239
rect 225420 6196 225472 6205
rect 226248 6239 226300 6248
rect 226248 6205 226282 6239
rect 226282 6205 226300 6239
rect 226248 6196 226300 6205
rect 226800 6196 226852 6248
rect 241520 6196 241572 6248
rect 216772 6171 216824 6180
rect 216772 6137 216781 6171
rect 216781 6137 216815 6171
rect 216815 6137 216824 6171
rect 216772 6128 216824 6137
rect 217140 6128 217192 6180
rect 215852 6060 215904 6069
rect 218152 6060 218204 6112
rect 218612 6128 218664 6180
rect 218704 6060 218756 6112
rect 220452 6128 220504 6180
rect 221648 6128 221700 6180
rect 222844 6128 222896 6180
rect 224776 6128 224828 6180
rect 225880 6171 225932 6180
rect 225880 6137 225889 6171
rect 225889 6137 225923 6171
rect 225923 6137 225932 6171
rect 225880 6128 225932 6137
rect 219808 6060 219860 6112
rect 220176 6060 220228 6112
rect 223120 6060 223172 6112
rect 223212 6060 223264 6112
rect 224868 6060 224920 6112
rect 226156 6060 226208 6112
rect 227076 6103 227128 6112
rect 227076 6069 227085 6103
rect 227085 6069 227119 6103
rect 227119 6069 227128 6103
rect 227076 6060 227128 6069
rect 227444 6128 227496 6180
rect 248696 6196 248748 6248
rect 249156 6307 249208 6316
rect 249156 6273 249165 6307
rect 249165 6273 249199 6307
rect 249199 6273 249208 6307
rect 249156 6264 249208 6273
rect 249340 6196 249392 6248
rect 248144 6128 248196 6180
rect 251364 6264 251416 6316
rect 255228 6332 255280 6384
rect 256332 6332 256384 6384
rect 259644 6332 259696 6384
rect 261760 6332 261812 6384
rect 263784 6332 263836 6384
rect 270224 6332 270276 6384
rect 239496 6060 239548 6112
rect 242900 6060 242952 6112
rect 247408 6060 247460 6112
rect 248604 6060 248656 6112
rect 248788 6060 248840 6112
rect 249064 6060 249116 6112
rect 249892 6060 249944 6112
rect 251456 6060 251508 6112
rect 253204 6264 253256 6316
rect 254032 6264 254084 6316
rect 255412 6264 255464 6316
rect 256792 6264 256844 6316
rect 258908 6264 258960 6316
rect 261576 6264 261628 6316
rect 262496 6264 262548 6316
rect 263140 6264 263192 6316
rect 265256 6264 265308 6316
rect 266544 6264 266596 6316
rect 266636 6307 266688 6316
rect 266636 6273 266645 6307
rect 266645 6273 266679 6307
rect 266679 6273 266688 6307
rect 266636 6264 266688 6273
rect 267188 6307 267240 6316
rect 267188 6273 267197 6307
rect 267197 6273 267231 6307
rect 267231 6273 267240 6307
rect 267188 6264 267240 6273
rect 267832 6307 267884 6316
rect 267832 6273 267841 6307
rect 267841 6273 267875 6307
rect 267875 6273 267884 6307
rect 267832 6264 267884 6273
rect 268936 6264 268988 6316
rect 269396 6307 269448 6316
rect 269396 6273 269405 6307
rect 269405 6273 269439 6307
rect 269439 6273 269448 6307
rect 269396 6264 269448 6273
rect 254584 6196 254636 6248
rect 256700 6196 256752 6248
rect 258816 6128 258868 6180
rect 262128 6196 262180 6248
rect 263232 6239 263284 6248
rect 263232 6205 263241 6239
rect 263241 6205 263275 6239
rect 263275 6205 263284 6239
rect 263232 6196 263284 6205
rect 264520 6239 264572 6248
rect 264520 6205 264529 6239
rect 264529 6205 264563 6239
rect 264563 6205 264572 6239
rect 264520 6196 264572 6205
rect 265716 6239 265768 6248
rect 265716 6205 265725 6239
rect 265725 6205 265759 6239
rect 265759 6205 265768 6239
rect 265716 6196 265768 6205
rect 270868 6400 270920 6452
rect 270500 6332 270552 6384
rect 261760 6128 261812 6180
rect 263048 6128 263100 6180
rect 268844 6128 268896 6180
rect 254400 6060 254452 6112
rect 255780 6060 255832 6112
rect 256424 6103 256476 6112
rect 256424 6069 256433 6103
rect 256433 6069 256467 6103
rect 256467 6069 256476 6103
rect 256424 6060 256476 6069
rect 256516 6060 256568 6112
rect 260380 6060 260432 6112
rect 261668 6060 261720 6112
rect 267648 6060 267700 6112
rect 270500 6239 270552 6248
rect 270500 6205 270509 6239
rect 270509 6205 270543 6239
rect 270543 6205 270552 6239
rect 270500 6196 270552 6205
rect 270868 6103 270920 6112
rect 270868 6069 270877 6103
rect 270877 6069 270911 6103
rect 270911 6069 270920 6103
rect 270868 6060 270920 6069
rect 34748 5958 34800 6010
rect 34812 5958 34864 6010
rect 34876 5958 34928 6010
rect 34940 5958 34992 6010
rect 35004 5958 35056 6010
rect 102345 5958 102397 6010
rect 102409 5958 102461 6010
rect 102473 5958 102525 6010
rect 102537 5958 102589 6010
rect 102601 5958 102653 6010
rect 169942 5958 169994 6010
rect 170006 5958 170058 6010
rect 170070 5958 170122 6010
rect 170134 5958 170186 6010
rect 170198 5958 170250 6010
rect 237539 5958 237591 6010
rect 237603 5958 237655 6010
rect 237667 5958 237719 6010
rect 237731 5958 237783 6010
rect 237795 5958 237847 6010
rect 46664 5899 46716 5908
rect 46664 5865 46673 5899
rect 46673 5865 46707 5899
rect 46707 5865 46716 5899
rect 46664 5856 46716 5865
rect 55772 5856 55824 5908
rect 94504 5856 94556 5908
rect 96068 5856 96120 5908
rect 96160 5899 96212 5908
rect 96160 5865 96169 5899
rect 96169 5865 96203 5899
rect 96203 5865 96212 5899
rect 96160 5856 96212 5865
rect 96436 5856 96488 5908
rect 100116 5899 100168 5908
rect 100116 5865 100125 5899
rect 100125 5865 100159 5899
rect 100159 5865 100168 5899
rect 100116 5856 100168 5865
rect 100944 5899 100996 5908
rect 100944 5865 100953 5899
rect 100953 5865 100987 5899
rect 100987 5865 100996 5899
rect 100944 5856 100996 5865
rect 101772 5856 101824 5908
rect 103428 5856 103480 5908
rect 106924 5856 106976 5908
rect 107200 5899 107252 5908
rect 107200 5865 107209 5899
rect 107209 5865 107243 5899
rect 107243 5865 107252 5899
rect 107200 5856 107252 5865
rect 107292 5856 107344 5908
rect 112168 5856 112220 5908
rect 112720 5856 112772 5908
rect 46480 5720 46532 5772
rect 53104 5720 53156 5772
rect 45652 5695 45704 5704
rect 45652 5661 45661 5695
rect 45661 5661 45695 5695
rect 45695 5661 45704 5695
rect 45652 5652 45704 5661
rect 46112 5695 46164 5704
rect 46112 5661 46121 5695
rect 46121 5661 46155 5695
rect 46155 5661 46164 5695
rect 46112 5652 46164 5661
rect 46940 5652 46992 5704
rect 47952 5652 48004 5704
rect 51540 5695 51592 5704
rect 51540 5661 51549 5695
rect 51549 5661 51583 5695
rect 51583 5661 51592 5695
rect 51540 5652 51592 5661
rect 35532 5584 35584 5636
rect 45376 5559 45428 5568
rect 45376 5525 45385 5559
rect 45385 5525 45419 5559
rect 45419 5525 45428 5559
rect 45376 5516 45428 5525
rect 45744 5627 45796 5636
rect 45744 5593 45753 5627
rect 45753 5593 45787 5627
rect 45787 5593 45796 5627
rect 45744 5584 45796 5593
rect 47216 5584 47268 5636
rect 52276 5695 52328 5704
rect 52276 5661 52285 5695
rect 52285 5661 52319 5695
rect 52319 5661 52328 5695
rect 52276 5652 52328 5661
rect 52368 5695 52420 5704
rect 52368 5661 52377 5695
rect 52377 5661 52411 5695
rect 52411 5661 52420 5695
rect 52368 5652 52420 5661
rect 55864 5652 55916 5704
rect 92664 5788 92716 5840
rect 94044 5788 94096 5840
rect 96620 5788 96672 5840
rect 97632 5788 97684 5840
rect 97908 5788 97960 5840
rect 101680 5788 101732 5840
rect 94596 5652 94648 5704
rect 94688 5695 94740 5704
rect 94688 5661 94697 5695
rect 94697 5661 94731 5695
rect 94731 5661 94740 5695
rect 94688 5652 94740 5661
rect 77484 5584 77536 5636
rect 48320 5559 48372 5568
rect 48320 5525 48329 5559
rect 48329 5525 48363 5559
rect 48363 5525 48372 5559
rect 48320 5516 48372 5525
rect 51448 5516 51500 5568
rect 52000 5559 52052 5568
rect 52000 5525 52009 5559
rect 52009 5525 52043 5559
rect 52043 5525 52052 5559
rect 52000 5516 52052 5525
rect 52552 5516 52604 5568
rect 53288 5559 53340 5568
rect 53288 5525 53297 5559
rect 53297 5525 53331 5559
rect 53331 5525 53340 5559
rect 53288 5516 53340 5525
rect 92388 5584 92440 5636
rect 95240 5584 95292 5636
rect 96068 5652 96120 5704
rect 96988 5720 97040 5772
rect 97080 5720 97132 5772
rect 97724 5763 97776 5772
rect 97724 5729 97733 5763
rect 97733 5729 97767 5763
rect 97767 5729 97776 5763
rect 97724 5720 97776 5729
rect 98460 5763 98512 5772
rect 98460 5729 98469 5763
rect 98469 5729 98503 5763
rect 98503 5729 98512 5763
rect 98460 5720 98512 5729
rect 98552 5720 98604 5772
rect 101496 5720 101548 5772
rect 102416 5720 102468 5772
rect 102968 5831 103020 5840
rect 102968 5797 102977 5831
rect 102977 5797 103011 5831
rect 103011 5797 103020 5831
rect 102968 5788 103020 5797
rect 104532 5788 104584 5840
rect 104900 5788 104952 5840
rect 108212 5788 108264 5840
rect 108764 5788 108816 5840
rect 96804 5652 96856 5704
rect 97356 5652 97408 5704
rect 99380 5652 99432 5704
rect 99564 5652 99616 5704
rect 98644 5584 98696 5636
rect 100392 5652 100444 5704
rect 100944 5695 100996 5704
rect 100944 5661 100953 5695
rect 100953 5661 100987 5695
rect 100987 5661 100996 5695
rect 100944 5652 100996 5661
rect 102324 5652 102376 5704
rect 102968 5652 103020 5704
rect 104532 5695 104584 5704
rect 104532 5661 104541 5695
rect 104541 5661 104575 5695
rect 104575 5661 104584 5695
rect 104532 5652 104584 5661
rect 105268 5652 105320 5704
rect 106372 5652 106424 5704
rect 108948 5720 109000 5772
rect 109040 5763 109092 5772
rect 109040 5729 109049 5763
rect 109049 5729 109083 5763
rect 109083 5729 109092 5763
rect 109040 5720 109092 5729
rect 109224 5763 109276 5772
rect 109224 5729 109233 5763
rect 109233 5729 109267 5763
rect 109267 5729 109276 5763
rect 109224 5720 109276 5729
rect 109960 5788 110012 5840
rect 112904 5788 112956 5840
rect 114836 5856 114888 5908
rect 116032 5856 116084 5908
rect 116584 5899 116636 5908
rect 116584 5865 116593 5899
rect 116593 5865 116627 5899
rect 116627 5865 116636 5899
rect 116584 5856 116636 5865
rect 116768 5899 116820 5908
rect 116768 5865 116777 5899
rect 116777 5865 116811 5899
rect 116811 5865 116820 5899
rect 116768 5856 116820 5865
rect 148324 5899 148376 5908
rect 113364 5788 113416 5840
rect 114652 5831 114704 5840
rect 114652 5797 114661 5831
rect 114661 5797 114695 5831
rect 114695 5797 114704 5831
rect 114652 5788 114704 5797
rect 114744 5788 114796 5840
rect 148324 5865 148333 5899
rect 148333 5865 148367 5899
rect 148367 5865 148376 5899
rect 148324 5856 148376 5865
rect 149796 5856 149848 5908
rect 107200 5652 107252 5704
rect 107384 5695 107436 5704
rect 107384 5661 107393 5695
rect 107393 5661 107427 5695
rect 107427 5661 107436 5695
rect 107384 5652 107436 5661
rect 110420 5652 110472 5704
rect 112168 5652 112220 5704
rect 113732 5720 113784 5772
rect 115204 5720 115256 5772
rect 115756 5720 115808 5772
rect 116492 5763 116544 5772
rect 116492 5729 116501 5763
rect 116501 5729 116535 5763
rect 116535 5729 116544 5763
rect 116492 5720 116544 5729
rect 100300 5584 100352 5636
rect 100668 5584 100720 5636
rect 101956 5584 102008 5636
rect 94412 5516 94464 5568
rect 96160 5516 96212 5568
rect 96436 5516 96488 5568
rect 97448 5516 97500 5568
rect 99012 5516 99064 5568
rect 100024 5516 100076 5568
rect 100116 5516 100168 5568
rect 107292 5584 107344 5636
rect 107660 5584 107712 5636
rect 110236 5584 110288 5636
rect 110880 5627 110932 5636
rect 110880 5593 110889 5627
rect 110889 5593 110923 5627
rect 110923 5593 110932 5627
rect 110880 5584 110932 5593
rect 111432 5627 111484 5636
rect 111432 5593 111441 5627
rect 111441 5593 111475 5627
rect 111475 5593 111484 5627
rect 111432 5584 111484 5593
rect 102968 5516 103020 5568
rect 104808 5516 104860 5568
rect 105452 5516 105504 5568
rect 108120 5516 108172 5568
rect 108672 5516 108724 5568
rect 114192 5652 114244 5704
rect 115112 5695 115164 5704
rect 115112 5661 115121 5695
rect 115121 5661 115155 5695
rect 115155 5661 115164 5695
rect 115112 5652 115164 5661
rect 115664 5652 115716 5704
rect 116400 5695 116452 5704
rect 116400 5661 116409 5695
rect 116409 5661 116443 5695
rect 116443 5661 116452 5695
rect 116400 5652 116452 5661
rect 114468 5584 114520 5636
rect 117320 5763 117372 5772
rect 117320 5729 117329 5763
rect 117329 5729 117363 5763
rect 117363 5729 117372 5763
rect 117320 5720 117372 5729
rect 117596 5720 117648 5772
rect 119068 5720 119120 5772
rect 119252 5652 119304 5704
rect 117504 5627 117556 5636
rect 117504 5593 117513 5627
rect 117513 5593 117547 5627
rect 117547 5593 117556 5627
rect 117504 5584 117556 5593
rect 118240 5584 118292 5636
rect 121460 5720 121512 5772
rect 121644 5788 121696 5840
rect 135536 5788 135588 5840
rect 113640 5516 113692 5568
rect 114008 5516 114060 5568
rect 116032 5516 116084 5568
rect 117596 5516 117648 5568
rect 118700 5516 118752 5568
rect 119896 5627 119948 5636
rect 119896 5593 119905 5627
rect 119905 5593 119939 5627
rect 119939 5593 119948 5627
rect 119896 5584 119948 5593
rect 120540 5584 120592 5636
rect 121920 5695 121972 5704
rect 121920 5661 121929 5695
rect 121929 5661 121963 5695
rect 121963 5661 121972 5695
rect 121920 5652 121972 5661
rect 127716 5695 127768 5704
rect 127716 5661 127725 5695
rect 127725 5661 127759 5695
rect 127759 5661 127768 5695
rect 127716 5652 127768 5661
rect 128084 5695 128136 5704
rect 128084 5661 128093 5695
rect 128093 5661 128127 5695
rect 128127 5661 128136 5695
rect 128084 5652 128136 5661
rect 137192 5720 137244 5772
rect 138756 5720 138808 5772
rect 140044 5763 140096 5772
rect 140044 5729 140053 5763
rect 140053 5729 140087 5763
rect 140087 5729 140096 5763
rect 140044 5720 140096 5729
rect 140688 5788 140740 5840
rect 120724 5584 120776 5636
rect 136088 5695 136140 5704
rect 136088 5661 136097 5695
rect 136097 5661 136131 5695
rect 136131 5661 136140 5695
rect 136088 5652 136140 5661
rect 138112 5652 138164 5704
rect 139768 5695 139820 5704
rect 139768 5661 139777 5695
rect 139777 5661 139811 5695
rect 139811 5661 139820 5695
rect 139768 5652 139820 5661
rect 132868 5627 132920 5636
rect 132868 5593 132877 5627
rect 132877 5593 132911 5627
rect 132911 5593 132920 5627
rect 132868 5584 132920 5593
rect 133236 5627 133288 5636
rect 133236 5593 133245 5627
rect 133245 5593 133279 5627
rect 133279 5593 133288 5627
rect 145104 5720 145156 5772
rect 154856 5856 154908 5908
rect 156420 5856 156472 5908
rect 157708 5899 157760 5908
rect 157708 5865 157717 5899
rect 157717 5865 157751 5899
rect 157751 5865 157760 5899
rect 157708 5856 157760 5865
rect 162124 5856 162176 5908
rect 142436 5695 142488 5704
rect 142436 5661 142445 5695
rect 142445 5661 142479 5695
rect 142479 5661 142488 5695
rect 142436 5652 142488 5661
rect 143264 5695 143316 5704
rect 143264 5661 143273 5695
rect 143273 5661 143307 5695
rect 143307 5661 143316 5695
rect 143264 5652 143316 5661
rect 143540 5652 143592 5704
rect 144828 5695 144880 5704
rect 144828 5661 144837 5695
rect 144837 5661 144871 5695
rect 144871 5661 144880 5695
rect 144828 5652 144880 5661
rect 147128 5720 147180 5772
rect 148508 5763 148560 5772
rect 148508 5729 148517 5763
rect 148517 5729 148551 5763
rect 148551 5729 148560 5763
rect 148508 5720 148560 5729
rect 133236 5584 133288 5593
rect 121184 5516 121236 5568
rect 135904 5516 135956 5568
rect 140320 5516 140372 5568
rect 143356 5516 143408 5568
rect 145564 5584 145616 5636
rect 147956 5652 148008 5704
rect 148140 5652 148192 5704
rect 151268 5720 151320 5772
rect 151360 5720 151412 5772
rect 151636 5763 151688 5772
rect 151636 5729 151645 5763
rect 151645 5729 151679 5763
rect 151679 5729 151688 5763
rect 151636 5720 151688 5729
rect 154488 5788 154540 5840
rect 188804 5831 188856 5840
rect 188804 5797 188813 5831
rect 188813 5797 188847 5831
rect 188847 5797 188856 5831
rect 188804 5788 188856 5797
rect 190460 5788 190512 5840
rect 210424 5856 210476 5908
rect 216680 5856 216732 5908
rect 217968 5856 218020 5908
rect 218428 5856 218480 5908
rect 218796 5856 218848 5908
rect 218980 5856 219032 5908
rect 222660 5856 222712 5908
rect 222752 5856 222804 5908
rect 225052 5856 225104 5908
rect 226892 5856 226944 5908
rect 245568 5856 245620 5908
rect 248052 5899 248104 5908
rect 248052 5865 248061 5899
rect 248061 5865 248095 5899
rect 248095 5865 248104 5899
rect 248052 5856 248104 5865
rect 248236 5899 248288 5908
rect 248236 5865 248245 5899
rect 248245 5865 248279 5899
rect 248279 5865 248288 5899
rect 248236 5856 248288 5865
rect 248788 5856 248840 5908
rect 251732 5856 251784 5908
rect 213368 5788 213420 5840
rect 213460 5788 213512 5840
rect 223212 5788 223264 5840
rect 223304 5788 223356 5840
rect 224776 5788 224828 5840
rect 153292 5720 153344 5772
rect 153844 5720 153896 5772
rect 154672 5763 154724 5772
rect 154672 5729 154681 5763
rect 154681 5729 154715 5763
rect 154715 5729 154724 5763
rect 154672 5720 154724 5729
rect 155868 5720 155920 5772
rect 158812 5720 158864 5772
rect 150256 5695 150308 5704
rect 150256 5661 150265 5695
rect 150265 5661 150299 5695
rect 150299 5661 150308 5695
rect 150256 5652 150308 5661
rect 150348 5652 150400 5704
rect 151176 5695 151228 5704
rect 151176 5661 151185 5695
rect 151185 5661 151219 5695
rect 151219 5661 151228 5695
rect 151176 5652 151228 5661
rect 151912 5695 151964 5704
rect 151912 5661 151921 5695
rect 151921 5661 151955 5695
rect 151955 5661 151964 5695
rect 151912 5652 151964 5661
rect 152096 5652 152148 5704
rect 152188 5695 152240 5704
rect 152188 5661 152197 5695
rect 152197 5661 152231 5695
rect 152231 5661 152240 5695
rect 152188 5652 152240 5661
rect 149704 5584 149756 5636
rect 149796 5584 149848 5636
rect 150900 5584 150952 5636
rect 152648 5516 152700 5568
rect 152832 5559 152884 5568
rect 152832 5525 152841 5559
rect 152841 5525 152875 5559
rect 152875 5525 152884 5559
rect 152832 5516 152884 5525
rect 154948 5695 155000 5704
rect 154948 5661 154957 5695
rect 154957 5661 154991 5695
rect 154991 5661 155000 5695
rect 154948 5652 155000 5661
rect 155960 5584 156012 5636
rect 156236 5584 156288 5636
rect 154856 5516 154908 5568
rect 156880 5618 156932 5670
rect 159732 5652 159784 5704
rect 159824 5652 159876 5704
rect 169668 5720 169720 5772
rect 185492 5720 185544 5772
rect 215852 5720 215904 5772
rect 217048 5763 217100 5772
rect 217048 5729 217057 5763
rect 217057 5729 217091 5763
rect 217091 5729 217100 5763
rect 217048 5720 217100 5729
rect 168288 5652 168340 5704
rect 168840 5695 168892 5704
rect 168840 5661 168849 5695
rect 168849 5661 168883 5695
rect 168883 5661 168892 5695
rect 168840 5652 168892 5661
rect 169208 5695 169260 5704
rect 169208 5661 169217 5695
rect 169217 5661 169251 5695
rect 169251 5661 169260 5695
rect 169208 5652 169260 5661
rect 169852 5695 169904 5704
rect 169852 5661 169861 5695
rect 169861 5661 169895 5695
rect 169895 5661 169904 5695
rect 169852 5652 169904 5661
rect 188804 5652 188856 5704
rect 207296 5695 207348 5704
rect 207296 5661 207305 5695
rect 207305 5661 207339 5695
rect 207339 5661 207348 5695
rect 207296 5652 207348 5661
rect 212816 5695 212868 5704
rect 212816 5661 212825 5695
rect 212825 5661 212859 5695
rect 212859 5661 212868 5695
rect 212816 5652 212868 5661
rect 157248 5584 157300 5636
rect 158628 5584 158680 5636
rect 168656 5584 168708 5636
rect 189540 5584 189592 5636
rect 206744 5584 206796 5636
rect 207112 5584 207164 5636
rect 207480 5627 207532 5636
rect 207480 5593 207489 5627
rect 207489 5593 207523 5627
rect 207523 5593 207532 5627
rect 207480 5584 207532 5593
rect 209136 5627 209188 5636
rect 209136 5593 209145 5627
rect 209145 5593 209179 5627
rect 209179 5593 209188 5627
rect 213368 5695 213420 5704
rect 213368 5661 213377 5695
rect 213377 5661 213411 5695
rect 213411 5661 213420 5695
rect 213368 5652 213420 5661
rect 213644 5695 213696 5704
rect 213644 5661 213653 5695
rect 213653 5661 213687 5695
rect 213687 5661 213696 5695
rect 213644 5652 213696 5661
rect 215208 5652 215260 5704
rect 216496 5652 216548 5704
rect 220820 5763 220872 5772
rect 220820 5729 220829 5763
rect 220829 5729 220863 5763
rect 220863 5729 220872 5763
rect 220820 5720 220872 5729
rect 222936 5720 222988 5772
rect 223488 5720 223540 5772
rect 224040 5763 224092 5772
rect 224040 5729 224049 5763
rect 224049 5729 224083 5763
rect 224083 5729 224092 5763
rect 224040 5720 224092 5729
rect 226064 5720 226116 5772
rect 226432 5788 226484 5840
rect 226616 5788 226668 5840
rect 227628 5788 227680 5840
rect 236460 5788 236512 5840
rect 247684 5788 247736 5840
rect 248420 5788 248472 5840
rect 248512 5788 248564 5840
rect 249432 5788 249484 5840
rect 250628 5788 250680 5840
rect 250996 5788 251048 5840
rect 256332 5856 256384 5908
rect 260840 5856 260892 5908
rect 263140 5899 263192 5908
rect 263140 5865 263149 5899
rect 263149 5865 263183 5899
rect 263183 5865 263192 5899
rect 263140 5856 263192 5865
rect 254584 5831 254636 5840
rect 254584 5797 254593 5831
rect 254593 5797 254627 5831
rect 254627 5797 254636 5831
rect 254584 5788 254636 5797
rect 254676 5788 254728 5840
rect 256792 5788 256844 5840
rect 239036 5720 239088 5772
rect 245568 5720 245620 5772
rect 247040 5720 247092 5772
rect 217876 5652 217928 5704
rect 209136 5584 209188 5593
rect 156788 5516 156840 5568
rect 167460 5516 167512 5568
rect 169392 5559 169444 5568
rect 169392 5525 169401 5559
rect 169401 5525 169435 5559
rect 169435 5525 169444 5559
rect 169392 5516 169444 5525
rect 171048 5516 171100 5568
rect 172612 5516 172664 5568
rect 189356 5516 189408 5568
rect 200764 5516 200816 5568
rect 210424 5516 210476 5568
rect 216036 5584 216088 5636
rect 216680 5584 216732 5636
rect 217232 5627 217284 5636
rect 217232 5593 217266 5627
rect 217266 5593 217284 5627
rect 217232 5584 217284 5593
rect 215116 5516 215168 5568
rect 216220 5516 216272 5568
rect 217140 5559 217192 5568
rect 217140 5525 217149 5559
rect 217149 5525 217183 5559
rect 217183 5525 217192 5559
rect 217140 5516 217192 5525
rect 218336 5695 218388 5704
rect 218336 5661 218345 5695
rect 218345 5661 218379 5695
rect 218379 5661 218388 5695
rect 218336 5652 218388 5661
rect 218060 5584 218112 5636
rect 218796 5652 218848 5704
rect 219532 5652 219584 5704
rect 220084 5584 220136 5636
rect 223212 5652 223264 5704
rect 223304 5695 223356 5704
rect 223304 5661 223313 5695
rect 223313 5661 223347 5695
rect 223347 5661 223356 5695
rect 223304 5652 223356 5661
rect 224316 5695 224368 5704
rect 224316 5661 224325 5695
rect 224325 5661 224359 5695
rect 224359 5661 224368 5695
rect 224316 5652 224368 5661
rect 224960 5652 225012 5704
rect 225696 5652 225748 5704
rect 246856 5652 246908 5704
rect 247960 5720 248012 5772
rect 248328 5720 248380 5772
rect 249800 5763 249852 5772
rect 249800 5729 249809 5763
rect 249809 5729 249843 5763
rect 249843 5729 249852 5763
rect 249800 5720 249852 5729
rect 249984 5720 250036 5772
rect 253296 5720 253348 5772
rect 259552 5788 259604 5840
rect 264888 5856 264940 5908
rect 265256 5899 265308 5908
rect 265256 5865 265265 5899
rect 265265 5865 265299 5899
rect 265299 5865 265308 5899
rect 265256 5856 265308 5865
rect 265440 5856 265492 5908
rect 265900 5856 265952 5908
rect 266176 5856 266228 5908
rect 269028 5856 269080 5908
rect 219716 5516 219768 5568
rect 227076 5584 227128 5636
rect 227720 5584 227772 5636
rect 243084 5584 243136 5636
rect 247040 5584 247092 5636
rect 247776 5627 247828 5636
rect 247776 5593 247785 5627
rect 247785 5593 247819 5627
rect 247819 5593 247828 5627
rect 247776 5584 247828 5593
rect 248236 5652 248288 5704
rect 248420 5652 248472 5704
rect 249156 5652 249208 5704
rect 250536 5652 250588 5704
rect 250720 5695 250772 5704
rect 250720 5661 250729 5695
rect 250729 5661 250763 5695
rect 250763 5661 250772 5695
rect 250720 5652 250772 5661
rect 238760 5516 238812 5568
rect 242992 5516 243044 5568
rect 248512 5516 248564 5568
rect 249340 5584 249392 5636
rect 249984 5516 250036 5568
rect 250444 5516 250496 5568
rect 253848 5695 253900 5704
rect 253848 5661 253857 5695
rect 253857 5661 253891 5695
rect 253891 5661 253900 5695
rect 253848 5652 253900 5661
rect 255412 5652 255464 5704
rect 256332 5652 256384 5704
rect 256792 5652 256844 5704
rect 257620 5652 257672 5704
rect 259184 5652 259236 5704
rect 260932 5720 260984 5772
rect 259644 5652 259696 5704
rect 260380 5695 260432 5704
rect 260380 5661 260389 5695
rect 260389 5661 260423 5695
rect 260423 5661 260432 5695
rect 260380 5652 260432 5661
rect 261576 5720 261628 5772
rect 251272 5584 251324 5636
rect 254308 5584 254360 5636
rect 254400 5627 254452 5636
rect 254400 5593 254409 5627
rect 254409 5593 254443 5627
rect 254443 5593 254452 5627
rect 254400 5584 254452 5593
rect 259460 5584 259512 5636
rect 261668 5695 261720 5704
rect 261668 5661 261677 5695
rect 261677 5661 261711 5695
rect 261711 5661 261720 5695
rect 261668 5652 261720 5661
rect 254216 5516 254268 5568
rect 255688 5516 255740 5568
rect 257804 5516 257856 5568
rect 260748 5627 260800 5636
rect 260748 5593 260757 5627
rect 260757 5593 260791 5627
rect 260791 5593 260800 5627
rect 260748 5584 260800 5593
rect 261024 5584 261076 5636
rect 259828 5516 259880 5568
rect 268384 5788 268436 5840
rect 268936 5788 268988 5840
rect 264428 5652 264480 5704
rect 264980 5720 265032 5772
rect 265256 5720 265308 5772
rect 268292 5720 268344 5772
rect 264888 5695 264940 5704
rect 264888 5661 264897 5695
rect 264897 5661 264931 5695
rect 264931 5661 264940 5695
rect 264888 5652 264940 5661
rect 265716 5652 265768 5704
rect 266912 5695 266964 5704
rect 266912 5661 266921 5695
rect 266921 5661 266955 5695
rect 266955 5661 266964 5695
rect 266912 5652 266964 5661
rect 269580 5695 269632 5704
rect 269580 5661 269589 5695
rect 269589 5661 269623 5695
rect 269623 5661 269632 5695
rect 269580 5652 269632 5661
rect 266360 5584 266412 5636
rect 268016 5584 268068 5636
rect 269948 5652 270000 5704
rect 269856 5584 269908 5636
rect 265716 5559 265768 5568
rect 265716 5525 265725 5559
rect 265725 5525 265759 5559
rect 265759 5525 265768 5559
rect 265716 5516 265768 5525
rect 265992 5516 266044 5568
rect 267096 5516 267148 5568
rect 271236 5584 271288 5636
rect 271144 5516 271196 5568
rect 271788 5516 271840 5568
rect 68546 5414 68598 5466
rect 68610 5414 68662 5466
rect 68674 5414 68726 5466
rect 68738 5414 68790 5466
rect 68802 5414 68854 5466
rect 136143 5414 136195 5466
rect 136207 5414 136259 5466
rect 136271 5414 136323 5466
rect 136335 5414 136387 5466
rect 136399 5414 136451 5466
rect 203740 5414 203792 5466
rect 203804 5414 203856 5466
rect 203868 5414 203920 5466
rect 203932 5414 203984 5466
rect 203996 5414 204048 5466
rect 271337 5414 271389 5466
rect 271401 5414 271453 5466
rect 271465 5414 271517 5466
rect 271529 5414 271581 5466
rect 271593 5414 271645 5466
rect 36084 5312 36136 5364
rect 37004 5312 37056 5364
rect 35808 5287 35860 5296
rect 35808 5253 35817 5287
rect 35817 5253 35851 5287
rect 35851 5253 35860 5287
rect 35808 5244 35860 5253
rect 36268 5287 36320 5296
rect 36268 5253 36277 5287
rect 36277 5253 36311 5287
rect 36311 5253 36320 5287
rect 36268 5244 36320 5253
rect 35900 5219 35952 5228
rect 35900 5185 35909 5219
rect 35909 5185 35943 5219
rect 35943 5185 35952 5219
rect 35900 5176 35952 5185
rect 35992 5176 36044 5228
rect 45836 5287 45888 5296
rect 45836 5253 45845 5287
rect 45845 5253 45879 5287
rect 45879 5253 45888 5287
rect 45836 5244 45888 5253
rect 46020 5244 46072 5296
rect 46664 5244 46716 5296
rect 36728 5176 36780 5228
rect 44088 5176 44140 5228
rect 46204 5219 46256 5228
rect 46204 5185 46213 5219
rect 46213 5185 46247 5219
rect 46247 5185 46256 5219
rect 46204 5176 46256 5185
rect 46572 5219 46624 5228
rect 46572 5185 46581 5219
rect 46581 5185 46615 5219
rect 46615 5185 46624 5219
rect 46572 5176 46624 5185
rect 46756 5176 46808 5228
rect 50988 5287 51040 5296
rect 50988 5253 50997 5287
rect 50997 5253 51031 5287
rect 51031 5253 51040 5287
rect 50988 5244 51040 5253
rect 51264 5219 51316 5228
rect 51264 5185 51273 5219
rect 51273 5185 51307 5219
rect 51307 5185 51316 5219
rect 51264 5176 51316 5185
rect 51356 5219 51408 5228
rect 51356 5185 51365 5219
rect 51365 5185 51399 5219
rect 51399 5185 51408 5219
rect 51356 5176 51408 5185
rect 51724 5219 51776 5228
rect 51724 5185 51733 5219
rect 51733 5185 51767 5219
rect 51767 5185 51776 5219
rect 51724 5176 51776 5185
rect 92388 5176 92440 5228
rect 95148 5312 95200 5364
rect 96068 5312 96120 5364
rect 96160 5312 96212 5364
rect 96436 5312 96488 5364
rect 96620 5312 96672 5364
rect 96988 5312 97040 5364
rect 98000 5312 98052 5364
rect 98092 5312 98144 5364
rect 100024 5312 100076 5364
rect 101404 5312 101456 5364
rect 95240 5244 95292 5296
rect 37096 5108 37148 5160
rect 46480 5108 46532 5160
rect 52092 5108 52144 5160
rect 53012 5108 53064 5160
rect 98460 5219 98512 5228
rect 98460 5185 98469 5219
rect 98469 5185 98503 5219
rect 98503 5185 98512 5219
rect 98460 5176 98512 5185
rect 99380 5176 99432 5228
rect 99564 5244 99616 5296
rect 100392 5244 100444 5296
rect 38752 5040 38804 5092
rect 40960 5040 41012 5092
rect 42248 5040 42300 5092
rect 47124 5083 47176 5092
rect 47124 5049 47133 5083
rect 47133 5049 47167 5083
rect 47167 5049 47176 5083
rect 47124 5040 47176 5049
rect 52184 5040 52236 5092
rect 52368 5040 52420 5092
rect 55864 5040 55916 5092
rect 94320 5040 94372 5092
rect 95976 5108 96028 5160
rect 95332 5040 95384 5092
rect 96620 5151 96672 5160
rect 96620 5117 96629 5151
rect 96629 5117 96663 5151
rect 96663 5117 96672 5151
rect 96620 5108 96672 5117
rect 97448 5108 97500 5160
rect 97724 5108 97776 5160
rect 98828 5108 98880 5160
rect 99564 5151 99616 5160
rect 99564 5117 99573 5151
rect 99573 5117 99607 5151
rect 99607 5117 99616 5151
rect 99564 5108 99616 5117
rect 100300 5219 100352 5228
rect 100300 5185 100309 5219
rect 100309 5185 100343 5219
rect 100343 5185 100352 5219
rect 100300 5176 100352 5185
rect 101312 5219 101364 5228
rect 101312 5185 101321 5219
rect 101321 5185 101355 5219
rect 101355 5185 101364 5219
rect 101312 5176 101364 5185
rect 101680 5219 101732 5228
rect 101680 5185 101689 5219
rect 101689 5185 101723 5219
rect 101723 5185 101732 5219
rect 101680 5176 101732 5185
rect 101864 5176 101916 5228
rect 102324 5219 102376 5228
rect 102324 5185 102333 5219
rect 102333 5185 102367 5219
rect 102367 5185 102376 5219
rect 102324 5176 102376 5185
rect 100576 5151 100628 5160
rect 100576 5117 100585 5151
rect 100585 5117 100619 5151
rect 100619 5117 100628 5151
rect 100576 5108 100628 5117
rect 102416 5151 102468 5160
rect 102416 5117 102425 5151
rect 102425 5117 102459 5151
rect 102459 5117 102468 5151
rect 102416 5108 102468 5117
rect 108856 5312 108908 5364
rect 115204 5312 115256 5364
rect 108028 5244 108080 5296
rect 110972 5287 111024 5296
rect 110972 5253 110981 5287
rect 110981 5253 111015 5287
rect 111015 5253 111024 5287
rect 110972 5244 111024 5253
rect 113548 5244 113600 5296
rect 113732 5244 113784 5296
rect 114284 5244 114336 5296
rect 107016 5219 107068 5228
rect 107016 5185 107025 5219
rect 107025 5185 107059 5219
rect 107059 5185 107068 5219
rect 107016 5176 107068 5185
rect 107660 5176 107712 5228
rect 108580 5219 108632 5228
rect 108580 5185 108589 5219
rect 108589 5185 108623 5219
rect 108623 5185 108632 5219
rect 108580 5176 108632 5185
rect 108672 5219 108724 5228
rect 108672 5185 108681 5219
rect 108681 5185 108715 5219
rect 108715 5185 108724 5219
rect 108672 5176 108724 5185
rect 105820 5108 105872 5160
rect 107200 5108 107252 5160
rect 110512 5176 110564 5228
rect 110788 5219 110840 5228
rect 110788 5185 110797 5219
rect 110797 5185 110831 5219
rect 110831 5185 110840 5219
rect 110788 5176 110840 5185
rect 110236 5108 110288 5160
rect 96896 5040 96948 5092
rect 99840 5040 99892 5092
rect 100024 5040 100076 5092
rect 111432 5040 111484 5092
rect 114192 5176 114244 5228
rect 114928 5244 114980 5296
rect 117320 5312 117372 5364
rect 122472 5312 122524 5364
rect 113732 5108 113784 5160
rect 116216 5219 116268 5228
rect 116216 5185 116225 5219
rect 116225 5185 116259 5219
rect 116259 5185 116268 5219
rect 116216 5176 116268 5185
rect 116032 5108 116084 5160
rect 117504 5244 117556 5296
rect 117596 5244 117648 5296
rect 143448 5244 143500 5296
rect 116952 5219 117004 5228
rect 116952 5185 116961 5219
rect 116961 5185 116995 5219
rect 116995 5185 117004 5219
rect 116952 5176 117004 5185
rect 119252 5176 119304 5228
rect 119988 5176 120040 5228
rect 116676 5108 116728 5160
rect 117412 5108 117464 5160
rect 121000 5219 121052 5228
rect 121000 5185 121009 5219
rect 121009 5185 121043 5219
rect 121043 5185 121052 5219
rect 121000 5176 121052 5185
rect 121828 5219 121880 5228
rect 121828 5185 121837 5219
rect 121837 5185 121871 5219
rect 121871 5185 121880 5219
rect 121828 5176 121880 5185
rect 121920 5176 121972 5228
rect 137468 5219 137520 5228
rect 137468 5185 137477 5219
rect 137477 5185 137511 5219
rect 137511 5185 137520 5219
rect 137468 5176 137520 5185
rect 138756 5219 138808 5228
rect 138756 5185 138765 5219
rect 138765 5185 138799 5219
rect 138799 5185 138808 5219
rect 138756 5176 138808 5185
rect 139400 5219 139452 5228
rect 139400 5185 139409 5219
rect 139409 5185 139443 5219
rect 139443 5185 139452 5219
rect 139400 5176 139452 5185
rect 121276 5108 121328 5160
rect 122748 5108 122800 5160
rect 114468 5040 114520 5092
rect 115112 5083 115164 5092
rect 115112 5049 115121 5083
rect 115121 5049 115155 5083
rect 115155 5049 115164 5083
rect 115112 5040 115164 5049
rect 120172 5040 120224 5092
rect 122380 5040 122432 5092
rect 137284 5040 137336 5092
rect 12072 4972 12124 5024
rect 35532 4972 35584 5024
rect 36820 5015 36872 5024
rect 36820 4981 36829 5015
rect 36829 4981 36863 5015
rect 36863 4981 36872 5015
rect 36820 4972 36872 4981
rect 36912 4972 36964 5024
rect 42616 4972 42668 5024
rect 92296 4972 92348 5024
rect 93308 4972 93360 5024
rect 94504 4972 94556 5024
rect 94688 4972 94740 5024
rect 99196 4972 99248 5024
rect 100116 4972 100168 5024
rect 100392 5015 100444 5024
rect 100392 4981 100401 5015
rect 100401 4981 100435 5015
rect 100435 4981 100444 5015
rect 101404 5015 101456 5024
rect 100392 4972 100444 4981
rect 101404 4981 101413 5015
rect 101413 4981 101447 5015
rect 101447 4981 101456 5015
rect 101404 4972 101456 4981
rect 101772 4972 101824 5024
rect 103152 5015 103204 5024
rect 103152 4981 103161 5015
rect 103161 4981 103195 5015
rect 103195 4981 103204 5015
rect 103152 4972 103204 4981
rect 103244 4972 103296 5024
rect 105728 4972 105780 5024
rect 106004 4972 106056 5024
rect 106924 4972 106976 5024
rect 108764 5015 108816 5024
rect 108764 4981 108773 5015
rect 108773 4981 108807 5015
rect 108807 4981 108816 5015
rect 108764 4972 108816 4981
rect 109776 4972 109828 5024
rect 109960 4972 110012 5024
rect 113364 4972 113416 5024
rect 114008 4972 114060 5024
rect 114192 5015 114244 5024
rect 114192 4981 114201 5015
rect 114201 4981 114235 5015
rect 114235 4981 114244 5015
rect 114192 4972 114244 4981
rect 114376 4972 114428 5024
rect 116032 4972 116084 5024
rect 116308 5015 116360 5024
rect 116308 4981 116317 5015
rect 116317 4981 116351 5015
rect 116351 4981 116360 5015
rect 116308 4972 116360 4981
rect 117136 4972 117188 5024
rect 118148 4972 118200 5024
rect 120908 5015 120960 5024
rect 120908 4981 120917 5015
rect 120917 4981 120951 5015
rect 120951 4981 120960 5015
rect 120908 4972 120960 4981
rect 121644 5015 121696 5024
rect 121644 4981 121653 5015
rect 121653 4981 121687 5015
rect 121687 4981 121696 5015
rect 121644 4972 121696 4981
rect 122288 5015 122340 5024
rect 122288 4981 122297 5015
rect 122297 4981 122331 5015
rect 122331 4981 122340 5015
rect 122288 4972 122340 4981
rect 135904 4972 135956 5024
rect 138112 5040 138164 5092
rect 139032 5040 139084 5092
rect 139584 5108 139636 5160
rect 139768 5108 139820 5160
rect 140320 5176 140372 5228
rect 141884 5176 141936 5228
rect 140044 5040 140096 5092
rect 145564 5312 145616 5364
rect 165620 5312 165672 5364
rect 143632 5176 143684 5228
rect 147496 5244 147548 5296
rect 148140 5176 148192 5228
rect 148508 5219 148560 5228
rect 148508 5185 148517 5219
rect 148517 5185 148551 5219
rect 148551 5185 148560 5219
rect 148508 5176 148560 5185
rect 149704 5219 149756 5228
rect 149704 5185 149718 5219
rect 149718 5185 149752 5219
rect 149752 5185 149756 5219
rect 150624 5244 150676 5296
rect 152648 5244 152700 5296
rect 153384 5244 153436 5296
rect 156420 5244 156472 5296
rect 149704 5176 149756 5185
rect 150532 5176 150584 5228
rect 145564 5108 145616 5160
rect 142528 5040 142580 5092
rect 146392 5151 146444 5160
rect 146392 5117 146401 5151
rect 146401 5117 146435 5151
rect 146435 5117 146444 5151
rect 146392 5108 146444 5117
rect 151728 5219 151780 5226
rect 151728 5185 151737 5219
rect 151737 5185 151771 5219
rect 151771 5185 151780 5219
rect 151728 5174 151780 5185
rect 150992 5151 151044 5160
rect 150992 5117 151001 5151
rect 151001 5117 151035 5151
rect 151035 5117 151044 5151
rect 150992 5108 151044 5117
rect 151912 5108 151964 5160
rect 152740 5176 152792 5228
rect 155960 5219 156012 5228
rect 155960 5185 155969 5219
rect 155969 5185 156003 5219
rect 156003 5185 156012 5219
rect 155960 5176 156012 5185
rect 159732 5176 159784 5228
rect 167460 5176 167512 5228
rect 167920 5312 167972 5364
rect 171048 5312 171100 5364
rect 206744 5312 206796 5364
rect 207480 5312 207532 5364
rect 169576 5176 169628 5228
rect 205640 5176 205692 5228
rect 206652 5219 206704 5228
rect 206652 5185 206661 5219
rect 206661 5185 206695 5219
rect 206695 5185 206704 5219
rect 206652 5176 206704 5185
rect 148140 5040 148192 5092
rect 139492 5015 139544 5024
rect 139492 4981 139501 5015
rect 139501 4981 139535 5015
rect 139535 4981 139544 5015
rect 139492 4972 139544 4981
rect 142252 5015 142304 5024
rect 142252 4981 142261 5015
rect 142261 4981 142295 5015
rect 142295 4981 142304 5015
rect 142252 4972 142304 4981
rect 142712 5015 142764 5024
rect 142712 4981 142721 5015
rect 142721 4981 142755 5015
rect 142755 4981 142764 5015
rect 142712 4972 142764 4981
rect 143448 5015 143500 5024
rect 143448 4981 143457 5015
rect 143457 4981 143491 5015
rect 143491 4981 143500 5015
rect 143448 4972 143500 4981
rect 145656 4972 145708 5024
rect 148324 5015 148376 5024
rect 148324 4981 148333 5015
rect 148333 4981 148367 5015
rect 148367 4981 148376 5015
rect 148324 4972 148376 4981
rect 148784 5083 148836 5092
rect 148784 5049 148793 5083
rect 148793 5049 148827 5083
rect 148827 5049 148836 5083
rect 148784 5040 148836 5049
rect 149244 4972 149296 5024
rect 149796 5015 149848 5024
rect 149796 4981 149805 5015
rect 149805 4981 149839 5015
rect 149839 4981 149848 5015
rect 149796 4972 149848 4981
rect 150440 5040 150492 5092
rect 150624 5040 150676 5092
rect 151268 5040 151320 5092
rect 151452 5083 151504 5092
rect 151452 5049 151461 5083
rect 151461 5049 151495 5083
rect 151495 5049 151504 5083
rect 151452 5040 151504 5049
rect 150348 4972 150400 5024
rect 154764 5151 154816 5160
rect 154764 5117 154773 5151
rect 154773 5117 154807 5151
rect 154807 5117 154816 5151
rect 154764 5108 154816 5117
rect 154948 5108 155000 5160
rect 156880 5108 156932 5160
rect 157800 5151 157852 5160
rect 157800 5117 157809 5151
rect 157809 5117 157843 5151
rect 157843 5117 157852 5151
rect 157800 5108 157852 5117
rect 167920 5108 167972 5160
rect 168104 5151 168156 5160
rect 168104 5117 168113 5151
rect 168113 5117 168147 5151
rect 168147 5117 168156 5151
rect 168104 5108 168156 5117
rect 168288 5151 168340 5160
rect 168288 5117 168297 5151
rect 168297 5117 168331 5151
rect 168331 5117 168340 5151
rect 168288 5108 168340 5117
rect 169852 5108 169904 5160
rect 205824 5108 205876 5160
rect 206836 5176 206888 5228
rect 214104 5312 214156 5364
rect 217140 5312 217192 5364
rect 210332 5176 210384 5228
rect 213184 5219 213236 5228
rect 213184 5185 213193 5219
rect 213193 5185 213227 5219
rect 213227 5185 213236 5219
rect 213184 5176 213236 5185
rect 213276 5176 213328 5228
rect 214380 5219 214432 5228
rect 214380 5185 214389 5219
rect 214389 5185 214423 5219
rect 214423 5185 214432 5219
rect 214380 5176 214432 5185
rect 214472 5219 214524 5228
rect 214472 5185 214506 5219
rect 214506 5185 214524 5219
rect 214472 5176 214524 5185
rect 207112 5108 207164 5160
rect 208400 5151 208452 5160
rect 208400 5117 208409 5151
rect 208409 5117 208443 5151
rect 208443 5117 208452 5151
rect 208400 5108 208452 5117
rect 208584 5108 208636 5160
rect 209228 5108 209280 5160
rect 213552 5108 213604 5160
rect 214104 5151 214156 5160
rect 214104 5117 214113 5151
rect 214113 5117 214147 5151
rect 214147 5117 214156 5151
rect 214104 5108 214156 5117
rect 152924 5040 152976 5092
rect 207572 5040 207624 5092
rect 207756 5040 207808 5092
rect 213460 5040 213512 5092
rect 153292 4972 153344 5024
rect 153936 4972 153988 5024
rect 154028 4972 154080 5024
rect 155316 4972 155368 5024
rect 165620 4972 165672 5024
rect 168288 4972 168340 5024
rect 172520 4972 172572 5024
rect 184572 4972 184624 5024
rect 206468 4972 206520 5024
rect 209964 5015 210016 5024
rect 209964 4981 209973 5015
rect 209973 4981 210007 5015
rect 210007 4981 210016 5015
rect 209964 4972 210016 4981
rect 214012 4972 214064 5024
rect 216128 5244 216180 5296
rect 216496 5287 216548 5296
rect 216496 5253 216505 5287
rect 216505 5253 216539 5287
rect 216539 5253 216548 5287
rect 216496 5244 216548 5253
rect 215576 5176 215628 5228
rect 215944 5219 215996 5228
rect 215944 5185 215953 5219
rect 215953 5185 215987 5219
rect 215987 5185 215996 5219
rect 215944 5176 215996 5185
rect 216312 5219 216364 5228
rect 216312 5185 216321 5219
rect 216321 5185 216355 5219
rect 216355 5185 216364 5219
rect 216312 5176 216364 5185
rect 217140 5219 217192 5228
rect 217140 5185 217149 5219
rect 217149 5185 217183 5219
rect 217183 5185 217192 5219
rect 217140 5176 217192 5185
rect 217784 5176 217836 5228
rect 219900 5312 219952 5364
rect 219716 5244 219768 5296
rect 221372 5312 221424 5364
rect 220084 5244 220136 5296
rect 220636 5244 220688 5296
rect 223120 5287 223172 5296
rect 223120 5253 223129 5287
rect 223129 5253 223163 5287
rect 223163 5253 223172 5287
rect 223120 5244 223172 5253
rect 223764 5312 223816 5364
rect 246212 5312 246264 5364
rect 224960 5244 225012 5296
rect 218796 5219 218848 5228
rect 218796 5185 218805 5219
rect 218805 5185 218839 5219
rect 218839 5185 218848 5219
rect 218796 5176 218848 5185
rect 215392 5108 215444 5160
rect 218428 5108 218480 5160
rect 218612 5108 218664 5160
rect 218980 5108 219032 5160
rect 220176 5219 220228 5228
rect 220176 5185 220185 5219
rect 220185 5185 220219 5219
rect 220219 5185 220228 5219
rect 220176 5176 220228 5185
rect 224408 5176 224460 5228
rect 242992 5244 243044 5296
rect 245016 5244 245068 5296
rect 246580 5244 246632 5296
rect 246948 5244 247000 5296
rect 247684 5287 247736 5296
rect 247684 5253 247693 5287
rect 247693 5253 247727 5287
rect 247727 5253 247736 5287
rect 247684 5244 247736 5253
rect 248144 5355 248196 5364
rect 248144 5321 248153 5355
rect 248153 5321 248187 5355
rect 248187 5321 248196 5355
rect 248144 5312 248196 5321
rect 248880 5287 248932 5296
rect 248880 5253 248889 5287
rect 248889 5253 248923 5287
rect 248923 5253 248932 5287
rect 248880 5244 248932 5253
rect 251732 5244 251784 5296
rect 220728 5108 220780 5160
rect 220820 5151 220872 5160
rect 220820 5117 220829 5151
rect 220829 5117 220863 5151
rect 220863 5117 220872 5151
rect 220820 5108 220872 5117
rect 221740 5108 221792 5160
rect 215116 5040 215168 5092
rect 216312 5040 216364 5092
rect 219532 5040 219584 5092
rect 215300 5015 215352 5024
rect 215300 4981 215309 5015
rect 215309 4981 215343 5015
rect 215343 4981 215352 5015
rect 215300 4972 215352 4981
rect 216956 5015 217008 5024
rect 216956 4981 216965 5015
rect 216965 4981 216999 5015
rect 216999 4981 217008 5015
rect 216956 4972 217008 4981
rect 217968 4972 218020 5024
rect 220912 5040 220964 5092
rect 222384 5040 222436 5092
rect 222936 5151 222988 5160
rect 222936 5117 222945 5151
rect 222945 5117 222979 5151
rect 222979 5117 222988 5151
rect 222936 5108 222988 5117
rect 223764 5151 223816 5160
rect 223764 5117 223773 5151
rect 223773 5117 223807 5151
rect 223807 5117 223816 5151
rect 223764 5108 223816 5117
rect 225144 5108 225196 5160
rect 225236 5151 225288 5160
rect 225236 5117 225245 5151
rect 225245 5117 225279 5151
rect 225279 5117 225288 5151
rect 225236 5108 225288 5117
rect 228640 5176 228692 5228
rect 246672 5176 246724 5228
rect 247040 5219 247092 5228
rect 247040 5185 247049 5219
rect 247049 5185 247083 5219
rect 247083 5185 247092 5219
rect 247040 5176 247092 5185
rect 247224 5176 247276 5228
rect 247868 5219 247920 5228
rect 247868 5185 247877 5219
rect 247877 5185 247911 5219
rect 247911 5185 247920 5219
rect 247868 5176 247920 5185
rect 223488 5040 223540 5092
rect 223580 5040 223632 5092
rect 227444 5108 227496 5160
rect 227628 5108 227680 5160
rect 237288 5108 237340 5160
rect 246856 5151 246908 5160
rect 246856 5117 246865 5151
rect 246865 5117 246899 5151
rect 246899 5117 246908 5151
rect 246856 5108 246908 5117
rect 248696 5219 248748 5228
rect 248696 5185 248705 5219
rect 248705 5185 248739 5219
rect 248739 5185 248748 5219
rect 248696 5176 248748 5185
rect 254492 5312 254544 5364
rect 256424 5312 256476 5364
rect 261576 5312 261628 5364
rect 262312 5312 262364 5364
rect 262496 5355 262548 5364
rect 262496 5321 262505 5355
rect 262505 5321 262539 5355
rect 262539 5321 262548 5355
rect 262496 5312 262548 5321
rect 263692 5312 263744 5364
rect 264980 5312 265032 5364
rect 266544 5312 266596 5364
rect 267740 5355 267792 5364
rect 267740 5321 267749 5355
rect 267749 5321 267783 5355
rect 267783 5321 267792 5355
rect 267740 5312 267792 5321
rect 268384 5312 268436 5364
rect 269396 5312 269448 5364
rect 254124 5244 254176 5296
rect 249156 5108 249208 5160
rect 252652 5108 252704 5160
rect 226064 5040 226116 5092
rect 247040 5040 247092 5092
rect 248328 5040 248380 5092
rect 251272 5040 251324 5092
rect 254676 5176 254728 5228
rect 253848 5108 253900 5160
rect 254584 5108 254636 5160
rect 255320 5287 255372 5296
rect 255320 5253 255329 5287
rect 255329 5253 255363 5287
rect 255363 5253 255372 5287
rect 255320 5244 255372 5253
rect 255412 5244 255464 5296
rect 255136 5219 255188 5228
rect 255136 5185 255145 5219
rect 255145 5185 255179 5219
rect 255179 5185 255188 5219
rect 255136 5176 255188 5185
rect 260288 5244 260340 5296
rect 257344 5176 257396 5228
rect 257620 5176 257672 5228
rect 259368 5176 259420 5228
rect 261024 5219 261076 5228
rect 261024 5185 261033 5219
rect 261033 5185 261067 5219
rect 261067 5185 261076 5219
rect 261024 5176 261076 5185
rect 262312 5219 262364 5228
rect 262312 5185 262321 5219
rect 262321 5185 262355 5219
rect 262355 5185 262364 5219
rect 262312 5176 262364 5185
rect 263600 5219 263652 5228
rect 263600 5185 263609 5219
rect 263609 5185 263643 5219
rect 263643 5185 263652 5219
rect 263600 5176 263652 5185
rect 264612 5219 264664 5228
rect 264612 5185 264621 5219
rect 264621 5185 264655 5219
rect 264655 5185 264664 5219
rect 264612 5176 264664 5185
rect 265256 5219 265308 5228
rect 265256 5185 265265 5219
rect 265265 5185 265299 5219
rect 265299 5185 265308 5219
rect 265256 5176 265308 5185
rect 265992 5244 266044 5296
rect 266452 5176 266504 5228
rect 266544 5219 266596 5228
rect 266544 5185 266553 5219
rect 266553 5185 266587 5219
rect 266587 5185 266596 5219
rect 266544 5176 266596 5185
rect 266912 5244 266964 5296
rect 267280 5176 267332 5228
rect 255412 5108 255464 5160
rect 256700 5108 256752 5160
rect 257528 5151 257580 5160
rect 257528 5117 257537 5151
rect 257537 5117 257571 5151
rect 257571 5117 257580 5151
rect 257528 5108 257580 5117
rect 258724 5108 258776 5160
rect 260104 5151 260156 5160
rect 260104 5117 260113 5151
rect 260113 5117 260147 5151
rect 260147 5117 260156 5151
rect 260104 5108 260156 5117
rect 261392 5151 261444 5160
rect 261392 5117 261401 5151
rect 261401 5117 261435 5151
rect 261435 5117 261444 5151
rect 261392 5108 261444 5117
rect 262588 5108 262640 5160
rect 267556 5219 267608 5228
rect 267556 5185 267565 5219
rect 267565 5185 267599 5219
rect 267599 5185 267608 5219
rect 267556 5176 267608 5185
rect 268292 5176 268344 5228
rect 267832 5108 267884 5160
rect 268200 5151 268252 5160
rect 268200 5117 268209 5151
rect 268209 5117 268243 5151
rect 268243 5117 268252 5151
rect 268200 5108 268252 5117
rect 268476 5176 268528 5228
rect 269856 5108 269908 5160
rect 244924 4972 244976 5024
rect 245108 4972 245160 5024
rect 246948 5015 247000 5024
rect 246948 4981 246957 5015
rect 246957 4981 246991 5015
rect 246991 4981 247000 5015
rect 246948 4972 247000 4981
rect 248788 4972 248840 5024
rect 251180 5015 251232 5024
rect 251180 4981 251189 5015
rect 251189 4981 251223 5015
rect 251223 4981 251232 5015
rect 251180 4972 251232 4981
rect 251732 5015 251784 5024
rect 251732 4981 251741 5015
rect 251741 4981 251775 5015
rect 251775 4981 251784 5015
rect 251732 4972 251784 4981
rect 253940 4972 253992 5024
rect 254492 5015 254544 5024
rect 254492 4981 254501 5015
rect 254501 4981 254535 5015
rect 254535 4981 254544 5015
rect 254492 4972 254544 4981
rect 255872 4972 255924 5024
rect 256424 4972 256476 5024
rect 258632 5040 258684 5092
rect 258816 4972 258868 5024
rect 265348 5040 265400 5092
rect 264980 4972 265032 5024
rect 265716 4972 265768 5024
rect 267096 4972 267148 5024
rect 267556 4972 267608 5024
rect 34748 4870 34800 4922
rect 34812 4870 34864 4922
rect 34876 4870 34928 4922
rect 34940 4870 34992 4922
rect 35004 4870 35056 4922
rect 102345 4870 102397 4922
rect 102409 4870 102461 4922
rect 102473 4870 102525 4922
rect 102537 4870 102589 4922
rect 102601 4870 102653 4922
rect 169942 4870 169994 4922
rect 170006 4870 170058 4922
rect 170070 4870 170122 4922
rect 170134 4870 170186 4922
rect 170198 4870 170250 4922
rect 237539 4870 237591 4922
rect 237603 4870 237655 4922
rect 237667 4870 237719 4922
rect 237731 4870 237783 4922
rect 237795 4870 237847 4922
rect 3332 4768 3384 4820
rect 29000 4768 29052 4820
rect 37004 4811 37056 4820
rect 37004 4777 37013 4811
rect 37013 4777 37047 4811
rect 37047 4777 37056 4811
rect 37004 4768 37056 4777
rect 40960 4811 41012 4820
rect 40960 4777 40969 4811
rect 40969 4777 41003 4811
rect 41003 4777 41012 4811
rect 40960 4768 41012 4777
rect 42800 4811 42852 4820
rect 42800 4777 42809 4811
rect 42809 4777 42843 4811
rect 42843 4777 42852 4811
rect 42800 4768 42852 4777
rect 44088 4768 44140 4820
rect 46756 4768 46808 4820
rect 48044 4811 48096 4820
rect 48044 4777 48053 4811
rect 48053 4777 48087 4811
rect 48087 4777 48096 4811
rect 48044 4768 48096 4777
rect 48136 4768 48188 4820
rect 55864 4768 55916 4820
rect 86960 4768 87012 4820
rect 99472 4768 99524 4820
rect 100116 4811 100168 4820
rect 100116 4777 100125 4811
rect 100125 4777 100159 4811
rect 100159 4777 100168 4811
rect 100116 4768 100168 4777
rect 100392 4768 100444 4820
rect 101220 4768 101272 4820
rect 102784 4768 102836 4820
rect 103980 4768 104032 4820
rect 106004 4811 106056 4820
rect 106004 4777 106013 4811
rect 106013 4777 106047 4811
rect 106047 4777 106056 4811
rect 106004 4768 106056 4777
rect 106096 4768 106148 4820
rect 45468 4700 45520 4752
rect 46388 4700 46440 4752
rect 36820 4632 36872 4684
rect 37096 4632 37148 4684
rect 42524 4632 42576 4684
rect 42708 4632 42760 4684
rect 46480 4632 46532 4684
rect 50896 4700 50948 4752
rect 51356 4700 51408 4752
rect 52368 4700 52420 4752
rect 92204 4743 92256 4752
rect 92204 4709 92213 4743
rect 92213 4709 92247 4743
rect 92247 4709 92256 4743
rect 92204 4700 92256 4709
rect 50988 4632 51040 4684
rect 51908 4632 51960 4684
rect 88340 4632 88392 4684
rect 92296 4632 92348 4684
rect 94504 4675 94556 4684
rect 94504 4641 94513 4675
rect 94513 4641 94547 4675
rect 94547 4641 94556 4675
rect 94504 4632 94556 4641
rect 94596 4632 94648 4684
rect 98368 4632 98420 4684
rect 98644 4675 98696 4684
rect 98644 4641 98653 4675
rect 98653 4641 98687 4675
rect 98687 4641 98696 4675
rect 98644 4632 98696 4641
rect 103796 4700 103848 4752
rect 105176 4700 105228 4752
rect 100852 4632 100904 4684
rect 103152 4632 103204 4684
rect 35624 4564 35676 4616
rect 21272 4428 21324 4480
rect 35440 4428 35492 4480
rect 35900 4496 35952 4548
rect 37280 4564 37332 4616
rect 38016 4564 38068 4616
rect 41788 4607 41840 4616
rect 41788 4573 41797 4607
rect 41797 4573 41831 4607
rect 41831 4573 41840 4607
rect 41788 4564 41840 4573
rect 42248 4607 42300 4616
rect 42248 4573 42257 4607
rect 42257 4573 42291 4607
rect 42291 4573 42300 4607
rect 42248 4564 42300 4573
rect 44364 4564 44416 4616
rect 46940 4564 46992 4616
rect 47032 4607 47084 4616
rect 47032 4573 47041 4607
rect 47041 4573 47075 4607
rect 47075 4573 47084 4607
rect 47032 4564 47084 4573
rect 47492 4607 47544 4616
rect 47492 4573 47501 4607
rect 47501 4573 47535 4607
rect 47535 4573 47544 4607
rect 47492 4564 47544 4573
rect 81440 4564 81492 4616
rect 92756 4607 92808 4616
rect 92756 4573 92765 4607
rect 92765 4573 92799 4607
rect 92799 4573 92808 4607
rect 92756 4564 92808 4573
rect 94320 4607 94372 4616
rect 94320 4573 94329 4607
rect 94329 4573 94363 4607
rect 94363 4573 94372 4607
rect 94320 4564 94372 4573
rect 96436 4564 96488 4616
rect 99380 4564 99432 4616
rect 36452 4539 36504 4548
rect 36452 4505 36461 4539
rect 36461 4505 36495 4539
rect 36495 4505 36504 4539
rect 36452 4496 36504 4505
rect 36544 4496 36596 4548
rect 41604 4428 41656 4480
rect 41880 4539 41932 4548
rect 41880 4505 41889 4539
rect 41889 4505 41923 4539
rect 41923 4505 41932 4539
rect 41880 4496 41932 4505
rect 45744 4496 45796 4548
rect 46204 4496 46256 4548
rect 48320 4496 48372 4548
rect 48504 4496 48556 4548
rect 49792 4496 49844 4548
rect 55864 4496 55916 4548
rect 93492 4496 93544 4548
rect 94688 4496 94740 4548
rect 96160 4539 96212 4548
rect 96160 4505 96169 4539
rect 96169 4505 96203 4539
rect 96203 4505 96212 4539
rect 96160 4496 96212 4505
rect 97172 4496 97224 4548
rect 44456 4428 44508 4480
rect 45284 4428 45336 4480
rect 47032 4428 47084 4480
rect 47860 4471 47912 4480
rect 47860 4437 47869 4471
rect 47869 4437 47903 4471
rect 47903 4437 47912 4471
rect 47860 4428 47912 4437
rect 47952 4428 48004 4480
rect 48688 4428 48740 4480
rect 49056 4428 49108 4480
rect 92388 4428 92440 4480
rect 93032 4428 93084 4480
rect 94596 4428 94648 4480
rect 95332 4428 95384 4480
rect 95608 4428 95660 4480
rect 97540 4428 97592 4480
rect 99564 4496 99616 4548
rect 100300 4564 100352 4616
rect 100576 4496 100628 4548
rect 104900 4564 104952 4616
rect 106096 4632 106148 4684
rect 106464 4743 106516 4752
rect 106464 4709 106473 4743
rect 106473 4709 106507 4743
rect 106507 4709 106516 4743
rect 106464 4700 106516 4709
rect 106924 4768 106976 4820
rect 108212 4768 108264 4820
rect 107384 4632 107436 4684
rect 113824 4768 113876 4820
rect 114008 4768 114060 4820
rect 114376 4768 114428 4820
rect 114468 4811 114520 4820
rect 114468 4777 114477 4811
rect 114477 4777 114511 4811
rect 114511 4777 114520 4811
rect 114468 4768 114520 4777
rect 117412 4768 117464 4820
rect 113364 4700 113416 4752
rect 114836 4700 114888 4752
rect 116308 4700 116360 4752
rect 118976 4768 119028 4820
rect 120908 4768 120960 4820
rect 118056 4700 118108 4752
rect 118700 4743 118752 4752
rect 118700 4709 118709 4743
rect 118709 4709 118743 4743
rect 118743 4709 118752 4743
rect 118700 4700 118752 4709
rect 105544 4564 105596 4616
rect 107200 4564 107252 4616
rect 108120 4564 108172 4616
rect 110880 4632 110932 4684
rect 111984 4632 112036 4684
rect 108764 4564 108816 4616
rect 109132 4607 109184 4616
rect 109132 4573 109141 4607
rect 109141 4573 109175 4607
rect 109175 4573 109184 4607
rect 109132 4564 109184 4573
rect 111616 4607 111668 4616
rect 111616 4573 111625 4607
rect 111625 4573 111659 4607
rect 111659 4573 111668 4607
rect 111616 4564 111668 4573
rect 113548 4632 113600 4684
rect 113088 4564 113140 4616
rect 115112 4632 115164 4684
rect 117872 4675 117924 4684
rect 117872 4641 117881 4675
rect 117881 4641 117915 4675
rect 117915 4641 117924 4675
rect 117872 4632 117924 4641
rect 118424 4632 118476 4684
rect 121828 4811 121880 4820
rect 121828 4777 121837 4811
rect 121837 4777 121871 4811
rect 121871 4777 121880 4811
rect 121828 4768 121880 4777
rect 137468 4768 137520 4820
rect 138848 4768 138900 4820
rect 114100 4607 114152 4616
rect 114100 4573 114109 4607
rect 114109 4573 114143 4607
rect 114143 4573 114152 4607
rect 114100 4564 114152 4573
rect 114284 4607 114336 4616
rect 114284 4573 114293 4607
rect 114293 4573 114327 4607
rect 114327 4573 114336 4607
rect 114284 4564 114336 4573
rect 114928 4607 114980 4616
rect 114928 4573 114937 4607
rect 114937 4573 114971 4607
rect 114971 4573 114980 4607
rect 114928 4564 114980 4573
rect 117320 4607 117372 4616
rect 117320 4573 117329 4607
rect 117329 4573 117363 4607
rect 117363 4573 117372 4607
rect 117320 4564 117372 4573
rect 118516 4564 118568 4616
rect 121000 4632 121052 4684
rect 122748 4675 122800 4684
rect 122748 4641 122757 4675
rect 122757 4641 122791 4675
rect 122791 4641 122800 4675
rect 122748 4632 122800 4641
rect 138572 4632 138624 4684
rect 138848 4675 138900 4684
rect 138848 4641 138857 4675
rect 138857 4641 138891 4675
rect 138891 4641 138900 4675
rect 138848 4632 138900 4641
rect 139124 4768 139176 4820
rect 140044 4768 140096 4820
rect 139860 4700 139912 4752
rect 119436 4607 119488 4616
rect 119436 4573 119445 4607
rect 119445 4573 119479 4607
rect 119479 4573 119488 4607
rect 119436 4564 119488 4573
rect 106556 4496 106608 4548
rect 101404 4428 101456 4480
rect 104348 4428 104400 4480
rect 104716 4428 104768 4480
rect 106234 4428 106286 4480
rect 107476 4428 107528 4480
rect 111800 4428 111852 4480
rect 113364 4496 113416 4548
rect 120080 4496 120132 4548
rect 121276 4607 121328 4616
rect 121276 4573 121285 4607
rect 121285 4573 121319 4607
rect 121319 4573 121328 4607
rect 122472 4607 122524 4616
rect 121276 4564 121328 4573
rect 122472 4573 122481 4607
rect 122481 4573 122515 4607
rect 122515 4573 122524 4607
rect 122472 4564 122524 4573
rect 138388 4607 138440 4616
rect 138388 4573 138397 4607
rect 138397 4573 138431 4607
rect 138431 4573 138440 4607
rect 138388 4564 138440 4573
rect 139216 4675 139268 4684
rect 139216 4641 139250 4675
rect 139250 4641 139268 4675
rect 139216 4632 139268 4641
rect 139952 4632 140004 4684
rect 140412 4632 140464 4684
rect 141148 4743 141200 4752
rect 141148 4709 141157 4743
rect 141157 4709 141191 4743
rect 141191 4709 141200 4743
rect 141148 4700 141200 4709
rect 142252 4768 142304 4820
rect 143448 4768 143500 4820
rect 143632 4811 143684 4820
rect 143632 4777 143641 4811
rect 143641 4777 143675 4811
rect 143675 4777 143684 4811
rect 143632 4768 143684 4777
rect 141424 4675 141476 4684
rect 141424 4641 141433 4675
rect 141433 4641 141467 4675
rect 141467 4641 141476 4675
rect 141424 4632 141476 4641
rect 141700 4675 141752 4684
rect 141700 4641 141709 4675
rect 141709 4641 141743 4675
rect 141743 4641 141752 4675
rect 141700 4632 141752 4641
rect 120448 4496 120500 4548
rect 121368 4496 121420 4548
rect 113732 4428 113784 4480
rect 118240 4428 118292 4480
rect 119988 4428 120040 4480
rect 122380 4428 122432 4480
rect 123024 4471 123076 4480
rect 123024 4437 123033 4471
rect 123033 4437 123067 4471
rect 123067 4437 123076 4471
rect 123024 4428 123076 4437
rect 135904 4428 135956 4480
rect 139676 4428 139728 4480
rect 141608 4564 141660 4616
rect 141700 4428 141752 4480
rect 142160 4428 142212 4480
rect 143172 4632 143224 4684
rect 144368 4632 144420 4684
rect 145012 4632 145064 4684
rect 145104 4675 145156 4684
rect 145104 4641 145113 4675
rect 145113 4641 145147 4675
rect 145147 4641 145156 4675
rect 145104 4632 145156 4641
rect 145380 4675 145432 4684
rect 145380 4641 145389 4675
rect 145389 4641 145423 4675
rect 145423 4641 145432 4675
rect 145380 4632 145432 4641
rect 146852 4632 146904 4684
rect 142988 4564 143040 4616
rect 145564 4564 145616 4616
rect 147128 4607 147180 4616
rect 147128 4573 147137 4607
rect 147137 4573 147171 4607
rect 147171 4573 147180 4607
rect 147128 4564 147180 4573
rect 148140 4564 148192 4616
rect 148416 4607 148468 4616
rect 148416 4573 148425 4607
rect 148425 4573 148459 4607
rect 148459 4573 148468 4607
rect 148416 4564 148468 4573
rect 148876 4632 148928 4684
rect 149888 4675 149940 4684
rect 149888 4641 149897 4675
rect 149897 4641 149931 4675
rect 149931 4641 149940 4675
rect 149888 4632 149940 4641
rect 150164 4675 150216 4684
rect 150164 4641 150173 4675
rect 150173 4641 150207 4675
rect 150207 4641 150216 4675
rect 150164 4632 150216 4641
rect 150348 4632 150400 4684
rect 150900 4768 150952 4820
rect 153108 4768 153160 4820
rect 154764 4768 154816 4820
rect 155868 4768 155920 4820
rect 161388 4768 161440 4820
rect 167184 4768 167236 4820
rect 153752 4700 153804 4752
rect 151360 4632 151412 4684
rect 152556 4675 152608 4684
rect 152556 4641 152565 4675
rect 152565 4641 152599 4675
rect 152599 4641 152608 4675
rect 152556 4632 152608 4641
rect 152832 4632 152884 4684
rect 153568 4675 153620 4684
rect 153568 4641 153577 4675
rect 153577 4641 153611 4675
rect 153611 4641 153620 4675
rect 153568 4632 153620 4641
rect 154580 4675 154632 4684
rect 154580 4641 154589 4675
rect 154589 4641 154623 4675
rect 154623 4641 154632 4675
rect 154580 4632 154632 4641
rect 156328 4700 156380 4752
rect 168104 4811 168156 4820
rect 168104 4777 168113 4811
rect 168113 4777 168147 4811
rect 168147 4777 168156 4811
rect 168104 4768 168156 4777
rect 186320 4768 186372 4820
rect 208584 4768 208636 4820
rect 216772 4768 216824 4820
rect 217232 4768 217284 4820
rect 222844 4768 222896 4820
rect 222936 4811 222988 4820
rect 222936 4777 222945 4811
rect 222945 4777 222979 4811
rect 222979 4777 222988 4811
rect 222936 4768 222988 4777
rect 223120 4768 223172 4820
rect 224316 4768 224368 4820
rect 169852 4700 169904 4752
rect 170864 4700 170916 4752
rect 205640 4700 205692 4752
rect 156052 4632 156104 4684
rect 156420 4632 156472 4684
rect 156512 4632 156564 4684
rect 158812 4632 158864 4684
rect 147312 4539 147364 4548
rect 147312 4505 147321 4539
rect 147321 4505 147355 4539
rect 147355 4505 147364 4539
rect 147312 4496 147364 4505
rect 148324 4496 148376 4548
rect 150072 4564 150124 4616
rect 151268 4607 151320 4616
rect 151268 4573 151277 4607
rect 151277 4573 151311 4607
rect 151311 4573 151320 4607
rect 151268 4564 151320 4573
rect 151544 4607 151596 4616
rect 151544 4573 151553 4607
rect 151553 4573 151587 4607
rect 151587 4573 151596 4607
rect 151544 4564 151596 4573
rect 155684 4607 155736 4616
rect 155684 4573 155693 4607
rect 155693 4573 155727 4607
rect 155727 4573 155736 4607
rect 155684 4564 155736 4573
rect 146300 4471 146352 4480
rect 146300 4437 146309 4471
rect 146309 4437 146343 4471
rect 146343 4437 146352 4471
rect 146300 4428 146352 4437
rect 148784 4428 148836 4480
rect 150808 4471 150860 4480
rect 150808 4437 150817 4471
rect 150817 4437 150851 4471
rect 150851 4437 150860 4471
rect 150808 4428 150860 4437
rect 152556 4428 152608 4480
rect 152832 4471 152884 4480
rect 152832 4437 152841 4471
rect 152841 4437 152875 4471
rect 152875 4437 152884 4471
rect 152832 4428 152884 4437
rect 152924 4428 152976 4480
rect 155868 4496 155920 4548
rect 155132 4428 155184 4480
rect 159456 4607 159508 4616
rect 159456 4573 159465 4607
rect 159465 4573 159499 4607
rect 159499 4573 159508 4607
rect 159456 4564 159508 4573
rect 159640 4564 159692 4616
rect 159732 4607 159784 4616
rect 159732 4573 159741 4607
rect 159741 4573 159775 4607
rect 159775 4573 159784 4607
rect 159732 4564 159784 4573
rect 164240 4632 164292 4684
rect 164332 4564 164384 4616
rect 167301 4675 167353 4684
rect 167301 4641 167331 4675
rect 167331 4641 167353 4675
rect 167301 4632 167353 4641
rect 168288 4632 168340 4684
rect 167184 4607 167236 4616
rect 167184 4573 167193 4607
rect 167193 4573 167227 4607
rect 167227 4573 167236 4607
rect 167184 4564 167236 4573
rect 167460 4607 167512 4616
rect 167460 4573 167469 4607
rect 167469 4573 167503 4607
rect 167503 4573 167512 4607
rect 167460 4564 167512 4573
rect 169392 4564 169444 4616
rect 205640 4607 205692 4616
rect 205640 4573 205649 4607
rect 205649 4573 205683 4607
rect 205683 4573 205692 4607
rect 205640 4564 205692 4573
rect 160376 4471 160428 4480
rect 160376 4437 160385 4471
rect 160385 4437 160419 4471
rect 160419 4437 160428 4471
rect 160376 4428 160428 4437
rect 165988 4471 166040 4480
rect 165988 4437 165997 4471
rect 165997 4437 166031 4471
rect 166031 4437 166040 4471
rect 165988 4428 166040 4437
rect 169852 4496 169904 4548
rect 205824 4607 205876 4616
rect 205824 4573 205833 4607
rect 205833 4573 205867 4607
rect 205867 4573 205876 4607
rect 205824 4564 205876 4573
rect 206652 4700 206704 4752
rect 210148 4700 210200 4752
rect 212172 4743 212224 4752
rect 212172 4709 212181 4743
rect 212181 4709 212215 4743
rect 212215 4709 212224 4743
rect 212172 4700 212224 4709
rect 206468 4675 206520 4684
rect 206468 4641 206477 4675
rect 206477 4641 206511 4675
rect 206511 4641 206520 4675
rect 206468 4632 206520 4641
rect 207940 4564 207992 4616
rect 211436 4632 211488 4684
rect 212632 4632 212684 4684
rect 213460 4675 213512 4684
rect 213460 4641 213469 4675
rect 213469 4641 213503 4675
rect 213503 4641 213512 4675
rect 213460 4632 213512 4641
rect 214564 4700 214616 4752
rect 219992 4700 220044 4752
rect 220820 4700 220872 4752
rect 208676 4564 208728 4616
rect 207572 4496 207624 4548
rect 208584 4496 208636 4548
rect 209044 4607 209096 4616
rect 209044 4573 209053 4607
rect 209053 4573 209087 4607
rect 209087 4573 209096 4607
rect 209044 4564 209096 4573
rect 209964 4564 210016 4616
rect 210516 4564 210568 4616
rect 211344 4564 211396 4616
rect 211620 4607 211672 4616
rect 211620 4573 211629 4607
rect 211629 4573 211663 4607
rect 211663 4573 211672 4607
rect 211620 4564 211672 4573
rect 211712 4564 211764 4616
rect 213000 4607 213052 4616
rect 213000 4573 213009 4607
rect 213009 4573 213043 4607
rect 213043 4573 213052 4607
rect 213000 4564 213052 4573
rect 213736 4607 213788 4616
rect 213736 4573 213745 4607
rect 213745 4573 213779 4607
rect 213779 4573 213788 4607
rect 213736 4564 213788 4573
rect 214012 4607 214064 4616
rect 214012 4573 214021 4607
rect 214021 4573 214055 4607
rect 214055 4573 214064 4607
rect 214012 4564 214064 4573
rect 167184 4428 167236 4480
rect 167276 4428 167328 4480
rect 187608 4428 187660 4480
rect 208860 4428 208912 4480
rect 209964 4428 210016 4480
rect 210148 4539 210200 4548
rect 210148 4505 210157 4539
rect 210157 4505 210191 4539
rect 210191 4505 210200 4539
rect 210148 4496 210200 4505
rect 214748 4632 214800 4684
rect 217968 4675 218020 4684
rect 217968 4641 217977 4675
rect 217977 4641 218011 4675
rect 218011 4641 218020 4675
rect 217968 4632 218020 4641
rect 218152 4675 218204 4684
rect 218152 4641 218161 4675
rect 218161 4641 218195 4675
rect 218195 4641 218204 4675
rect 218152 4632 218204 4641
rect 218428 4632 218480 4684
rect 219072 4632 219124 4684
rect 219440 4675 219492 4684
rect 219440 4641 219449 4675
rect 219449 4641 219483 4675
rect 219483 4641 219492 4675
rect 219440 4632 219492 4641
rect 220360 4632 220412 4684
rect 221740 4675 221792 4684
rect 216404 4496 216456 4548
rect 217048 4539 217100 4548
rect 217048 4505 217057 4539
rect 217057 4505 217091 4539
rect 217091 4505 217100 4539
rect 217048 4496 217100 4505
rect 217968 4496 218020 4548
rect 218336 4496 218388 4548
rect 218428 4496 218480 4548
rect 218704 4496 218756 4548
rect 218888 4496 218940 4548
rect 220728 4564 220780 4616
rect 221740 4641 221749 4675
rect 221749 4641 221783 4675
rect 221783 4641 221792 4675
rect 221740 4632 221792 4641
rect 223764 4700 223816 4752
rect 224132 4700 224184 4752
rect 224684 4700 224736 4752
rect 224960 4768 225012 4820
rect 228088 4768 228140 4820
rect 228272 4768 228324 4820
rect 245568 4768 245620 4820
rect 246488 4768 246540 4820
rect 246948 4811 247000 4820
rect 246948 4777 246957 4811
rect 246957 4777 246991 4811
rect 246991 4777 247000 4811
rect 246948 4768 247000 4777
rect 248052 4768 248104 4820
rect 251180 4768 251232 4820
rect 252468 4768 252520 4820
rect 253020 4768 253072 4820
rect 253204 4768 253256 4820
rect 225420 4700 225472 4752
rect 227812 4700 227864 4752
rect 247500 4700 247552 4752
rect 248236 4700 248288 4752
rect 219532 4496 219584 4548
rect 220636 4496 220688 4548
rect 210240 4471 210292 4480
rect 210240 4437 210249 4471
rect 210249 4437 210283 4471
rect 210283 4437 210292 4471
rect 210240 4428 210292 4437
rect 210332 4428 210384 4480
rect 215116 4428 215168 4480
rect 216220 4428 216272 4480
rect 220176 4428 220228 4480
rect 220268 4428 220320 4480
rect 222016 4607 222068 4616
rect 222016 4573 222025 4607
rect 222025 4573 222059 4607
rect 222059 4573 222068 4607
rect 222016 4564 222068 4573
rect 222108 4607 222160 4616
rect 222108 4573 222142 4607
rect 222142 4573 222160 4607
rect 222108 4564 222160 4573
rect 222292 4607 222344 4616
rect 222292 4573 222301 4607
rect 222301 4573 222335 4607
rect 222335 4573 222344 4607
rect 222292 4564 222344 4573
rect 223212 4564 223264 4616
rect 223764 4564 223816 4616
rect 222844 4496 222896 4548
rect 223488 4496 223540 4548
rect 224776 4564 224828 4616
rect 227352 4607 227404 4616
rect 227352 4573 227361 4607
rect 227361 4573 227395 4607
rect 227395 4573 227404 4607
rect 227352 4564 227404 4573
rect 227812 4564 227864 4616
rect 224132 4496 224184 4548
rect 244924 4607 244976 4616
rect 244924 4573 244933 4607
rect 244933 4573 244967 4607
rect 244967 4573 244976 4607
rect 244924 4564 244976 4573
rect 245568 4607 245620 4616
rect 245568 4573 245577 4607
rect 245577 4573 245611 4607
rect 245611 4573 245620 4607
rect 245568 4564 245620 4573
rect 247684 4632 247736 4684
rect 249064 4675 249116 4684
rect 249064 4641 249073 4675
rect 249073 4641 249107 4675
rect 249107 4641 249116 4675
rect 249064 4632 249116 4641
rect 246304 4496 246356 4548
rect 246580 4496 246632 4548
rect 246856 4607 246908 4616
rect 246856 4573 246865 4607
rect 246865 4573 246899 4607
rect 246899 4573 246908 4607
rect 246856 4564 246908 4573
rect 246948 4607 247000 4616
rect 246948 4573 246957 4607
rect 246957 4573 246991 4607
rect 246991 4573 247000 4607
rect 246948 4564 247000 4573
rect 247132 4564 247184 4616
rect 247316 4496 247368 4548
rect 247776 4564 247828 4616
rect 248236 4496 248288 4548
rect 248880 4607 248932 4616
rect 248880 4573 248889 4607
rect 248889 4573 248923 4607
rect 248923 4573 248932 4607
rect 248880 4564 248932 4573
rect 253112 4700 253164 4752
rect 251640 4632 251692 4684
rect 253020 4632 253072 4684
rect 251272 4539 251324 4548
rect 251272 4505 251281 4539
rect 251281 4505 251315 4539
rect 251315 4505 251324 4539
rect 251272 4496 251324 4505
rect 251364 4496 251416 4548
rect 222108 4428 222160 4480
rect 222292 4428 222344 4480
rect 223120 4428 223172 4480
rect 224040 4471 224092 4480
rect 224040 4437 224049 4471
rect 224049 4437 224083 4471
rect 224083 4437 224092 4471
rect 224040 4428 224092 4437
rect 224592 4428 224644 4480
rect 227536 4428 227588 4480
rect 245384 4471 245436 4480
rect 245384 4437 245393 4471
rect 245393 4437 245427 4471
rect 245427 4437 245436 4471
rect 245384 4428 245436 4437
rect 247132 4471 247184 4480
rect 247132 4437 247141 4471
rect 247141 4437 247175 4471
rect 247175 4437 247184 4471
rect 247132 4428 247184 4437
rect 249708 4428 249760 4480
rect 252560 4539 252612 4548
rect 252560 4505 252569 4539
rect 252569 4505 252603 4539
rect 252603 4505 252612 4539
rect 252560 4496 252612 4505
rect 252836 4607 252888 4616
rect 252836 4573 252845 4607
rect 252845 4573 252879 4607
rect 252879 4573 252888 4607
rect 254492 4700 254544 4752
rect 258632 4768 258684 4820
rect 259184 4811 259236 4820
rect 259184 4777 259193 4811
rect 259193 4777 259227 4811
rect 259227 4777 259236 4811
rect 259184 4768 259236 4777
rect 260288 4768 260340 4820
rect 265164 4768 265216 4820
rect 265348 4811 265400 4820
rect 265348 4777 265357 4811
rect 265357 4777 265391 4811
rect 265391 4777 265400 4811
rect 265348 4768 265400 4777
rect 265716 4768 265768 4820
rect 266912 4768 266964 4820
rect 269028 4768 269080 4820
rect 270316 4768 270368 4820
rect 256608 4675 256660 4684
rect 256608 4641 256617 4675
rect 256617 4641 256651 4675
rect 256651 4641 256660 4675
rect 256608 4632 256660 4641
rect 257344 4632 257396 4684
rect 252836 4564 252888 4573
rect 252744 4428 252796 4480
rect 252928 4539 252980 4548
rect 252928 4505 252937 4539
rect 252937 4505 252971 4539
rect 252971 4505 252980 4539
rect 252928 4496 252980 4505
rect 255872 4607 255924 4616
rect 255872 4573 255881 4607
rect 255881 4573 255915 4607
rect 255915 4573 255924 4607
rect 255872 4564 255924 4573
rect 256424 4607 256476 4616
rect 256424 4573 256433 4607
rect 256433 4573 256467 4607
rect 256467 4573 256476 4607
rect 256424 4564 256476 4573
rect 258724 4632 258776 4684
rect 258264 4539 258316 4548
rect 258264 4505 258273 4539
rect 258273 4505 258307 4539
rect 258307 4505 258316 4539
rect 258264 4496 258316 4505
rect 259368 4564 259420 4616
rect 259828 4607 259880 4616
rect 259828 4573 259837 4607
rect 259837 4573 259871 4607
rect 259871 4573 259880 4607
rect 259828 4564 259880 4573
rect 272156 4700 272208 4752
rect 264336 4564 264388 4616
rect 265072 4564 265124 4616
rect 268476 4632 268528 4684
rect 266176 4607 266228 4616
rect 266176 4573 266185 4607
rect 266185 4573 266219 4607
rect 266219 4573 266228 4607
rect 266176 4564 266228 4573
rect 267648 4564 267700 4616
rect 269212 4564 269264 4616
rect 269856 4607 269908 4616
rect 269856 4573 269865 4607
rect 269865 4573 269899 4607
rect 269899 4573 269908 4607
rect 269856 4564 269908 4573
rect 271052 4564 271104 4616
rect 271144 4564 271196 4616
rect 271972 4564 272024 4616
rect 259184 4496 259236 4548
rect 260840 4496 260892 4548
rect 263600 4496 263652 4548
rect 267188 4496 267240 4548
rect 267280 4539 267332 4548
rect 267280 4505 267289 4539
rect 267289 4505 267323 4539
rect 267323 4505 267332 4539
rect 267280 4496 267332 4505
rect 267556 4496 267608 4548
rect 269028 4496 269080 4548
rect 271696 4496 271748 4548
rect 259828 4428 259880 4480
rect 261576 4471 261628 4480
rect 261576 4437 261585 4471
rect 261585 4437 261619 4471
rect 261619 4437 261628 4471
rect 261576 4428 261628 4437
rect 269764 4428 269816 4480
rect 270408 4428 270460 4480
rect 271052 4428 271104 4480
rect 68546 4326 68598 4378
rect 68610 4326 68662 4378
rect 68674 4326 68726 4378
rect 68738 4326 68790 4378
rect 68802 4326 68854 4378
rect 136143 4326 136195 4378
rect 136207 4326 136259 4378
rect 136271 4326 136323 4378
rect 136335 4326 136387 4378
rect 136399 4326 136451 4378
rect 203740 4326 203792 4378
rect 203804 4326 203856 4378
rect 203868 4326 203920 4378
rect 203932 4326 203984 4378
rect 203996 4326 204048 4378
rect 271337 4326 271389 4378
rect 271401 4326 271453 4378
rect 271465 4326 271517 4378
rect 271529 4326 271581 4378
rect 271593 4326 271645 4378
rect 4436 4156 4488 4208
rect 38384 4224 38436 4276
rect 41880 4224 41932 4276
rect 18052 4088 18104 4140
rect 36728 4088 36780 4140
rect 37832 4156 37884 4208
rect 38660 4156 38712 4208
rect 38752 4199 38804 4208
rect 38752 4165 38761 4199
rect 38761 4165 38795 4199
rect 38795 4165 38804 4199
rect 38752 4156 38804 4165
rect 44364 4156 44416 4208
rect 44456 4199 44508 4208
rect 44456 4165 44465 4199
rect 44465 4165 44499 4199
rect 44499 4165 44508 4199
rect 44456 4156 44508 4165
rect 45744 4224 45796 4276
rect 48412 4224 48464 4276
rect 49792 4267 49844 4276
rect 49792 4233 49801 4267
rect 49801 4233 49835 4267
rect 49835 4233 49844 4267
rect 49792 4224 49844 4233
rect 51080 4224 51132 4276
rect 55864 4224 55916 4276
rect 100668 4224 100720 4276
rect 105820 4224 105872 4276
rect 38016 4131 38068 4140
rect 38016 4097 38025 4131
rect 38025 4097 38059 4131
rect 38059 4097 38068 4131
rect 38016 4088 38068 4097
rect 38384 4131 38436 4140
rect 38384 4097 38393 4131
rect 38393 4097 38427 4131
rect 38427 4097 38436 4131
rect 38384 4088 38436 4097
rect 42616 4131 42668 4140
rect 42616 4097 42625 4131
rect 42625 4097 42659 4131
rect 42659 4097 42668 4131
rect 42616 4088 42668 4097
rect 43352 4088 43404 4140
rect 45560 4199 45612 4208
rect 45560 4165 45569 4199
rect 45569 4165 45603 4199
rect 45603 4165 45612 4199
rect 45560 4156 45612 4165
rect 49148 4156 49200 4208
rect 49516 4156 49568 4208
rect 44732 4131 44784 4140
rect 44732 4097 44741 4131
rect 44741 4097 44775 4131
rect 44775 4097 44784 4131
rect 44732 4088 44784 4097
rect 45100 4088 45152 4140
rect 48596 4088 48648 4140
rect 49056 4088 49108 4140
rect 50896 4131 50948 4140
rect 50896 4097 50905 4131
rect 50905 4097 50939 4131
rect 50939 4097 50948 4131
rect 50896 4088 50948 4097
rect 51172 4156 51224 4208
rect 51724 4156 51776 4208
rect 94504 4156 94556 4208
rect 51816 4088 51868 4140
rect 12808 4020 12860 4072
rect 36912 4020 36964 4072
rect 38476 4020 38528 4072
rect 42524 4020 42576 4072
rect 45468 4020 45520 4072
rect 47124 4020 47176 4072
rect 47952 4020 48004 4072
rect 51632 4020 51684 4072
rect 52092 4020 52144 4072
rect 92572 4088 92624 4140
rect 92940 4131 92992 4140
rect 92940 4097 92949 4131
rect 92949 4097 92983 4131
rect 92983 4097 92992 4131
rect 92940 4088 92992 4097
rect 93584 4131 93636 4140
rect 93584 4097 93593 4131
rect 93593 4097 93627 4131
rect 93627 4097 93636 4131
rect 93584 4088 93636 4097
rect 94596 4131 94648 4140
rect 94596 4097 94605 4131
rect 94605 4097 94639 4131
rect 94639 4097 94648 4131
rect 94596 4088 94648 4097
rect 8024 3952 8076 4004
rect 36544 3952 36596 4004
rect 36820 3952 36872 4004
rect 37372 3952 37424 4004
rect 38936 3995 38988 4004
rect 38936 3961 38945 3995
rect 38945 3961 38979 3995
rect 38979 3961 38988 3995
rect 38936 3952 38988 3961
rect 39028 3952 39080 4004
rect 44088 3952 44140 4004
rect 94412 4020 94464 4072
rect 94780 4063 94832 4072
rect 94780 4029 94789 4063
rect 94789 4029 94823 4063
rect 94823 4029 94832 4063
rect 94780 4020 94832 4029
rect 95148 4020 95200 4072
rect 96344 4088 96396 4140
rect 98644 4156 98696 4208
rect 99196 4156 99248 4208
rect 101496 4156 101548 4208
rect 102048 4131 102100 4140
rect 102048 4097 102057 4131
rect 102057 4097 102091 4131
rect 102091 4097 102100 4131
rect 102048 4088 102100 4097
rect 105544 4156 105596 4208
rect 106004 4156 106056 4208
rect 106280 4156 106332 4208
rect 106924 4156 106976 4208
rect 108120 4156 108172 4208
rect 111616 4224 111668 4276
rect 118240 4224 118292 4276
rect 116676 4156 116728 4208
rect 96160 4063 96212 4072
rect 96160 4029 96169 4063
rect 96169 4029 96203 4063
rect 96203 4029 96212 4063
rect 96160 4020 96212 4029
rect 96896 4063 96948 4072
rect 96896 4029 96905 4063
rect 96905 4029 96939 4063
rect 96939 4029 96948 4063
rect 96896 4020 96948 4029
rect 89720 3952 89772 4004
rect 93216 3952 93268 4004
rect 96712 3952 96764 4004
rect 98276 4020 98328 4072
rect 97816 3952 97868 4004
rect 101220 4020 101272 4072
rect 102968 4020 103020 4072
rect 108764 4131 108816 4140
rect 108764 4097 108773 4131
rect 108773 4097 108807 4131
rect 108807 4097 108816 4131
rect 108764 4088 108816 4097
rect 105176 4020 105228 4072
rect 105360 4020 105412 4072
rect 105912 4063 105964 4072
rect 105912 4029 105921 4063
rect 105921 4029 105955 4063
rect 105955 4029 105964 4063
rect 105912 4020 105964 4029
rect 106004 4020 106056 4072
rect 108120 4020 108172 4072
rect 108856 4020 108908 4072
rect 109960 4088 110012 4140
rect 110236 4131 110288 4140
rect 110236 4097 110245 4131
rect 110245 4097 110279 4131
rect 110279 4097 110288 4131
rect 110236 4088 110288 4097
rect 114192 4131 114244 4140
rect 114192 4097 114201 4131
rect 114201 4097 114235 4131
rect 114235 4097 114244 4131
rect 114192 4088 114244 4097
rect 117044 4131 117096 4140
rect 117044 4097 117053 4131
rect 117053 4097 117087 4131
rect 117087 4097 117096 4131
rect 117044 4088 117096 4097
rect 120080 4156 120132 4208
rect 122104 4156 122156 4208
rect 110512 4063 110564 4072
rect 29000 3884 29052 3936
rect 36728 3884 36780 3936
rect 41144 3884 41196 3936
rect 41880 3884 41932 3936
rect 42432 3884 42484 3936
rect 44456 3884 44508 3936
rect 45744 3927 45796 3936
rect 45744 3893 45753 3927
rect 45753 3893 45787 3927
rect 45787 3893 45796 3927
rect 45744 3884 45796 3893
rect 47676 3884 47728 3936
rect 48412 3884 48464 3936
rect 66720 3927 66772 3936
rect 66720 3893 66729 3927
rect 66729 3893 66763 3927
rect 66763 3893 66772 3927
rect 66720 3884 66772 3893
rect 93308 3884 93360 3936
rect 95240 3884 95292 3936
rect 102876 3952 102928 4004
rect 100208 3884 100260 3936
rect 104164 3884 104216 3936
rect 104348 3884 104400 3936
rect 105268 3995 105320 4004
rect 105268 3961 105277 3995
rect 105277 3961 105311 3995
rect 105311 3961 105320 3995
rect 105268 3952 105320 3961
rect 108764 3952 108816 4004
rect 105452 3884 105504 3936
rect 107844 3884 107896 3936
rect 108856 3927 108908 3936
rect 108856 3893 108865 3927
rect 108865 3893 108899 3927
rect 108899 3893 108908 3927
rect 108856 3884 108908 3893
rect 109316 3884 109368 3936
rect 110512 4029 110521 4063
rect 110521 4029 110555 4063
rect 110555 4029 110564 4063
rect 110512 4020 110564 4029
rect 110788 4020 110840 4072
rect 111156 4020 111208 4072
rect 111616 4063 111668 4072
rect 111616 4029 111625 4063
rect 111625 4029 111659 4063
rect 111659 4029 111668 4063
rect 111616 4020 111668 4029
rect 111800 4063 111852 4072
rect 111800 4029 111809 4063
rect 111809 4029 111843 4063
rect 111843 4029 111852 4063
rect 111800 4020 111852 4029
rect 111984 4020 112036 4072
rect 114560 4020 114612 4072
rect 114744 4063 114796 4072
rect 114744 4029 114753 4063
rect 114753 4029 114787 4063
rect 114787 4029 114796 4063
rect 114744 4020 114796 4029
rect 112168 3952 112220 4004
rect 109776 3884 109828 3936
rect 110328 3884 110380 3936
rect 111708 3884 111760 3936
rect 117228 4063 117280 4072
rect 117228 4029 117237 4063
rect 117237 4029 117271 4063
rect 117271 4029 117280 4063
rect 117228 4020 117280 4029
rect 118240 4131 118292 4140
rect 118240 4097 118249 4131
rect 118249 4097 118283 4131
rect 118283 4097 118292 4131
rect 118240 4088 118292 4097
rect 120448 4131 120500 4140
rect 120448 4097 120457 4131
rect 120457 4097 120491 4131
rect 120491 4097 120500 4131
rect 120448 4088 120500 4097
rect 121000 4088 121052 4140
rect 117964 4063 118016 4072
rect 117964 4029 117973 4063
rect 117973 4029 118007 4063
rect 118007 4029 118016 4063
rect 117964 4020 118016 4029
rect 118056 4063 118108 4072
rect 118056 4029 118090 4063
rect 118090 4029 118108 4063
rect 118056 4020 118108 4029
rect 121460 4063 121512 4072
rect 121460 4029 121469 4063
rect 121469 4029 121503 4063
rect 121503 4029 121512 4063
rect 121460 4020 121512 4029
rect 122472 4020 122524 4072
rect 120264 3952 120316 4004
rect 121920 3952 121972 4004
rect 122012 3952 122064 4004
rect 138848 4156 138900 4208
rect 141148 4156 141200 4208
rect 142712 4156 142764 4208
rect 139400 4131 139452 4140
rect 139400 4097 139409 4131
rect 139409 4097 139443 4131
rect 139443 4097 139452 4131
rect 139400 4088 139452 4097
rect 141884 4088 141936 4140
rect 142988 4088 143040 4140
rect 145104 4156 145156 4208
rect 148416 4224 148468 4276
rect 150992 4224 151044 4276
rect 153844 4224 153896 4276
rect 155684 4224 155736 4276
rect 165988 4224 166040 4276
rect 167276 4224 167328 4276
rect 167368 4224 167420 4276
rect 170864 4224 170916 4276
rect 176660 4224 176712 4276
rect 209320 4224 209372 4276
rect 210148 4224 210200 4276
rect 150348 4156 150400 4208
rect 139032 4020 139084 4072
rect 139768 4020 139820 4072
rect 120080 3884 120132 3936
rect 120908 3884 120960 3936
rect 139492 3952 139544 4004
rect 140688 4063 140740 4072
rect 140688 4029 140697 4063
rect 140697 4029 140731 4063
rect 140731 4029 140740 4063
rect 140688 4020 140740 4029
rect 140964 4063 141016 4072
rect 140964 4029 140973 4063
rect 140973 4029 141007 4063
rect 141007 4029 141016 4063
rect 140964 4020 141016 4029
rect 142528 4020 142580 4072
rect 144736 4020 144788 4072
rect 145840 4063 145892 4072
rect 145840 4029 145849 4063
rect 145849 4029 145883 4063
rect 145883 4029 145892 4063
rect 145840 4020 145892 4029
rect 146852 4131 146904 4140
rect 146852 4097 146861 4131
rect 146861 4097 146895 4131
rect 146895 4097 146904 4131
rect 146852 4088 146904 4097
rect 147496 4131 147548 4140
rect 147496 4097 147505 4131
rect 147505 4097 147539 4131
rect 147539 4097 147548 4131
rect 147496 4088 147548 4097
rect 147956 4131 148008 4140
rect 147956 4097 147965 4131
rect 147965 4097 147999 4131
rect 147999 4097 148008 4131
rect 147956 4088 148008 4097
rect 149152 4088 149204 4140
rect 152832 4156 152884 4208
rect 154948 4156 155000 4208
rect 156236 4156 156288 4208
rect 160284 4156 160336 4208
rect 161296 4156 161348 4208
rect 163596 4156 163648 4208
rect 167184 4156 167236 4208
rect 168012 4156 168064 4208
rect 205640 4156 205692 4208
rect 215576 4156 215628 4208
rect 215944 4224 215996 4276
rect 216772 4224 216824 4276
rect 220912 4224 220964 4276
rect 221004 4224 221056 4276
rect 216312 4156 216364 4208
rect 150808 4131 150860 4140
rect 150808 4097 150817 4131
rect 150817 4097 150851 4131
rect 150851 4097 150860 4131
rect 150808 4088 150860 4097
rect 153200 4131 153252 4140
rect 153200 4097 153209 4131
rect 153209 4097 153243 4131
rect 153243 4097 153252 4131
rect 153200 4088 153252 4097
rect 146208 4020 146260 4072
rect 138940 3927 138992 3936
rect 138940 3893 138949 3927
rect 138949 3893 138983 3927
rect 138983 3893 138992 3927
rect 138940 3884 138992 3893
rect 142160 3952 142212 4004
rect 139676 3884 139728 3936
rect 140780 3884 140832 3936
rect 142344 3884 142396 3936
rect 143264 3952 143316 4004
rect 143448 3884 143500 3936
rect 145564 3884 145616 3936
rect 147864 3952 147916 4004
rect 149060 4020 149112 4072
rect 149428 4020 149480 4072
rect 149980 3952 150032 4004
rect 152004 4063 152056 4072
rect 152004 4029 152013 4063
rect 152013 4029 152047 4063
rect 152047 4029 152056 4063
rect 152004 4020 152056 4029
rect 153476 4020 153528 4072
rect 153936 4020 153988 4072
rect 154120 4063 154172 4072
rect 154120 4029 154129 4063
rect 154129 4029 154163 4063
rect 154163 4029 154172 4063
rect 154120 4020 154172 4029
rect 154212 4063 154264 4072
rect 154212 4029 154246 4063
rect 154246 4029 154264 4063
rect 154212 4020 154264 4029
rect 155224 4020 155276 4072
rect 156236 4020 156288 4072
rect 157064 4063 157116 4072
rect 157064 4029 157073 4063
rect 157073 4029 157107 4063
rect 157107 4029 157116 4063
rect 157064 4020 157116 4029
rect 152188 3952 152240 4004
rect 147312 3884 147364 3936
rect 149244 3884 149296 3936
rect 152740 3884 152792 3936
rect 154948 3952 155000 4004
rect 158168 3952 158220 4004
rect 158444 4063 158496 4072
rect 158444 4029 158453 4063
rect 158453 4029 158487 4063
rect 158487 4029 158496 4063
rect 158444 4020 158496 4029
rect 158536 4020 158588 4072
rect 164332 4088 164384 4140
rect 167736 4088 167788 4140
rect 190460 4131 190512 4140
rect 190460 4097 190469 4131
rect 190469 4097 190503 4131
rect 190503 4097 190512 4131
rect 190460 4088 190512 4097
rect 206560 4131 206612 4140
rect 206560 4097 206569 4131
rect 206569 4097 206603 4131
rect 206603 4097 206612 4131
rect 206560 4088 206612 4097
rect 206652 4131 206704 4140
rect 206652 4097 206661 4131
rect 206661 4097 206695 4131
rect 206695 4097 206704 4131
rect 206652 4088 206704 4097
rect 206744 4131 206796 4140
rect 206744 4097 206753 4131
rect 206753 4097 206787 4131
rect 206787 4097 206796 4131
rect 206744 4088 206796 4097
rect 213184 4131 213236 4140
rect 213184 4097 213193 4131
rect 213193 4097 213227 4131
rect 213227 4097 213236 4131
rect 213184 4088 213236 4097
rect 160008 4063 160060 4072
rect 160008 4029 160017 4063
rect 160017 4029 160051 4063
rect 160051 4029 160060 4063
rect 160008 4020 160060 4029
rect 168196 4020 168248 4072
rect 160376 3952 160428 4004
rect 161388 3952 161440 4004
rect 154580 3884 154632 3936
rect 158536 3884 158588 3936
rect 164240 3884 164292 3936
rect 164332 3884 164384 3936
rect 167368 3884 167420 3936
rect 167460 3884 167512 3936
rect 168288 3927 168340 3936
rect 168288 3893 168297 3927
rect 168297 3893 168331 3927
rect 168331 3893 168340 3927
rect 168288 3884 168340 3893
rect 191196 3884 191248 3936
rect 207480 4063 207532 4072
rect 207480 4029 207489 4063
rect 207489 4029 207523 4063
rect 207523 4029 207532 4063
rect 207480 4020 207532 4029
rect 209320 4063 209372 4072
rect 209320 4029 209329 4063
rect 209329 4029 209363 4063
rect 209363 4029 209372 4063
rect 209320 4020 209372 4029
rect 209780 4063 209832 4072
rect 209780 4029 209789 4063
rect 209789 4029 209823 4063
rect 209823 4029 209832 4063
rect 209780 4020 209832 4029
rect 209964 4063 210016 4072
rect 209964 4029 209973 4063
rect 209973 4029 210007 4063
rect 210007 4029 210016 4063
rect 209964 4020 210016 4029
rect 208308 3952 208360 4004
rect 209228 3952 209280 4004
rect 212080 4020 212132 4072
rect 213920 4063 213972 4072
rect 213920 4029 213929 4063
rect 213929 4029 213963 4063
rect 213963 4029 213972 4063
rect 213920 4020 213972 4029
rect 216588 4020 216640 4072
rect 216680 4020 216732 4072
rect 217876 4156 217928 4208
rect 216956 4088 217008 4140
rect 220268 4131 220320 4140
rect 220268 4097 220277 4131
rect 220277 4097 220311 4131
rect 220311 4097 220320 4131
rect 220268 4088 220320 4097
rect 223304 4224 223356 4276
rect 225144 4224 225196 4276
rect 242992 4224 243044 4276
rect 226984 4156 227036 4208
rect 217692 4020 217744 4072
rect 218152 4020 218204 4072
rect 218428 4063 218480 4072
rect 218428 4029 218437 4063
rect 218437 4029 218471 4063
rect 218471 4029 218480 4063
rect 218428 4020 218480 4029
rect 218704 4063 218756 4072
rect 218704 4029 218713 4063
rect 218713 4029 218747 4063
rect 218747 4029 218756 4063
rect 218704 4020 218756 4029
rect 218796 4063 218848 4072
rect 218796 4029 218830 4063
rect 218830 4029 218848 4063
rect 218796 4020 218848 4029
rect 218980 4063 219032 4072
rect 218980 4029 218989 4063
rect 218989 4029 219023 4063
rect 219023 4029 219032 4063
rect 218980 4020 219032 4029
rect 219164 4020 219216 4072
rect 219348 4020 219400 4072
rect 221004 4063 221056 4072
rect 221004 4029 221013 4063
rect 221013 4029 221047 4063
rect 221047 4029 221056 4063
rect 221004 4020 221056 4029
rect 221188 4020 221240 4072
rect 221924 4020 221976 4072
rect 222292 4020 222344 4072
rect 223304 4020 223356 4072
rect 223580 4063 223632 4072
rect 223580 4029 223589 4063
rect 223589 4029 223623 4063
rect 223623 4029 223632 4063
rect 223580 4020 223632 4029
rect 223856 4097 223865 4106
rect 223865 4097 223899 4106
rect 223899 4097 223908 4106
rect 223856 4054 223908 4097
rect 224132 4131 224184 4140
rect 224132 4097 224141 4131
rect 224141 4097 224175 4131
rect 224175 4097 224184 4131
rect 224132 4088 224184 4097
rect 224776 4131 224828 4140
rect 224776 4097 224785 4131
rect 224785 4097 224819 4131
rect 224819 4097 224828 4131
rect 224776 4088 224828 4097
rect 227260 4088 227312 4140
rect 211804 3952 211856 4004
rect 213184 3952 213236 4004
rect 215300 3952 215352 4004
rect 209688 3884 209740 3936
rect 217968 3952 218020 4004
rect 219808 3952 219860 4004
rect 220360 3952 220412 4004
rect 220728 3995 220780 4004
rect 220728 3961 220737 3995
rect 220737 3961 220771 3995
rect 220771 3961 220780 3995
rect 220728 3952 220780 3961
rect 216036 3927 216088 3936
rect 216036 3893 216045 3927
rect 216045 3893 216079 3927
rect 216079 3893 216088 3927
rect 216036 3884 216088 3893
rect 217416 3884 217468 3936
rect 221096 3884 221148 3936
rect 222108 3884 222160 3936
rect 224776 3884 224828 3936
rect 225420 4063 225472 4072
rect 225420 4029 225429 4063
rect 225429 4029 225463 4063
rect 225463 4029 225472 4063
rect 225420 4020 225472 4029
rect 226708 4063 226760 4072
rect 226708 4029 226717 4063
rect 226717 4029 226751 4063
rect 226751 4029 226760 4063
rect 226708 4020 226760 4029
rect 227628 4020 227680 4072
rect 229836 4020 229888 4072
rect 242900 4020 242952 4072
rect 247040 4224 247092 4276
rect 245016 4131 245068 4140
rect 245016 4097 245030 4131
rect 245030 4097 245064 4131
rect 245064 4097 245068 4131
rect 245016 4088 245068 4097
rect 246856 4156 246908 4208
rect 251272 4156 251324 4208
rect 247132 4088 247184 4140
rect 247224 4088 247276 4140
rect 247592 4131 247644 4140
rect 247592 4097 247601 4131
rect 247601 4097 247635 4131
rect 247635 4097 247644 4131
rect 247592 4088 247644 4097
rect 250996 4131 251048 4140
rect 250996 4097 251005 4131
rect 251005 4097 251039 4131
rect 251039 4097 251048 4131
rect 250996 4088 251048 4097
rect 252560 4156 252612 4208
rect 252652 4088 252704 4140
rect 252928 4088 252980 4140
rect 253664 4088 253716 4140
rect 253848 4156 253900 4208
rect 254124 4131 254176 4140
rect 254124 4097 254133 4131
rect 254133 4097 254167 4131
rect 254167 4097 254176 4131
rect 254124 4088 254176 4097
rect 257896 4156 257948 4208
rect 258264 4224 258316 4276
rect 266268 4224 266320 4276
rect 266452 4224 266504 4276
rect 268568 4267 268620 4276
rect 268568 4233 268577 4267
rect 268577 4233 268611 4267
rect 268611 4233 268620 4267
rect 268568 4224 268620 4233
rect 270776 4267 270828 4276
rect 270776 4233 270785 4267
rect 270785 4233 270819 4267
rect 270819 4233 270828 4267
rect 270776 4224 270828 4233
rect 258540 4156 258592 4208
rect 259828 4199 259880 4208
rect 259828 4165 259837 4199
rect 259837 4165 259871 4199
rect 259871 4165 259880 4199
rect 259828 4156 259880 4165
rect 257344 4131 257396 4140
rect 257344 4097 257353 4131
rect 257353 4097 257387 4131
rect 257387 4097 257396 4131
rect 257344 4088 257396 4097
rect 257436 4088 257488 4140
rect 257620 4131 257672 4140
rect 257620 4097 257629 4131
rect 257629 4097 257663 4131
rect 257663 4097 257672 4131
rect 257620 4088 257672 4097
rect 248420 4020 248472 4072
rect 248696 4063 248748 4072
rect 248696 4029 248705 4063
rect 248705 4029 248739 4063
rect 248739 4029 248748 4063
rect 248696 4020 248748 4029
rect 249432 4020 249484 4072
rect 250812 4020 250864 4072
rect 251364 4020 251416 4072
rect 253020 4063 253072 4072
rect 253020 4029 253029 4063
rect 253029 4029 253063 4063
rect 253063 4029 253072 4063
rect 253020 4020 253072 4029
rect 254584 4020 254636 4072
rect 227352 3952 227404 4004
rect 227444 3952 227496 4004
rect 244188 3952 244240 4004
rect 244464 3952 244516 4004
rect 257068 4020 257120 4072
rect 261760 4088 261812 4140
rect 228180 3884 228232 3936
rect 229744 3884 229796 3936
rect 244280 3884 244332 3936
rect 252836 3927 252888 3936
rect 252836 3893 252845 3927
rect 252845 3893 252879 3927
rect 252879 3893 252888 3927
rect 252836 3884 252888 3893
rect 254032 3884 254084 3936
rect 254124 3927 254176 3936
rect 254124 3893 254133 3927
rect 254133 3893 254167 3927
rect 254167 3893 254176 3927
rect 254124 3884 254176 3893
rect 259276 4020 259328 4072
rect 260748 4063 260800 4072
rect 260748 4029 260757 4063
rect 260757 4029 260791 4063
rect 260791 4029 260800 4063
rect 260748 4020 260800 4029
rect 257896 3952 257948 4004
rect 265532 4088 265584 4140
rect 267740 4156 267792 4208
rect 266912 4088 266964 4140
rect 267004 4131 267056 4140
rect 267004 4097 267013 4131
rect 267013 4097 267047 4131
rect 267047 4097 267056 4131
rect 267004 4088 267056 4097
rect 267096 4131 267148 4140
rect 267096 4097 267105 4131
rect 267105 4097 267139 4131
rect 267139 4097 267148 4131
rect 267096 4088 267148 4097
rect 269304 4131 269356 4140
rect 269304 4097 269313 4131
rect 269313 4097 269347 4131
rect 269347 4097 269356 4131
rect 269304 4088 269356 4097
rect 270868 4088 270920 4140
rect 272064 4088 272116 4140
rect 267280 4020 267332 4072
rect 257344 3927 257396 3936
rect 257344 3893 257353 3927
rect 257353 3893 257387 3927
rect 257387 3893 257396 3927
rect 257344 3884 257396 3893
rect 257436 3884 257488 3936
rect 258816 3927 258868 3936
rect 258816 3893 258825 3927
rect 258825 3893 258859 3927
rect 258859 3893 258868 3927
rect 258816 3884 258868 3893
rect 259276 3927 259328 3936
rect 259276 3893 259285 3927
rect 259285 3893 259319 3927
rect 259319 3893 259328 3927
rect 259276 3884 259328 3893
rect 261760 3884 261812 3936
rect 262036 3884 262088 3936
rect 269488 3995 269540 4004
rect 269488 3961 269497 3995
rect 269497 3961 269531 3995
rect 269531 3961 269540 3995
rect 269488 3952 269540 3961
rect 270500 3952 270552 4004
rect 264796 3884 264848 3936
rect 265808 3884 265860 3936
rect 267740 3884 267792 3936
rect 34748 3782 34800 3834
rect 34812 3782 34864 3834
rect 34876 3782 34928 3834
rect 34940 3782 34992 3834
rect 35004 3782 35056 3834
rect 102345 3782 102397 3834
rect 102409 3782 102461 3834
rect 102473 3782 102525 3834
rect 102537 3782 102589 3834
rect 102601 3782 102653 3834
rect 169942 3782 169994 3834
rect 170006 3782 170058 3834
rect 170070 3782 170122 3834
rect 170134 3782 170186 3834
rect 170198 3782 170250 3834
rect 237539 3782 237591 3834
rect 237603 3782 237655 3834
rect 237667 3782 237719 3834
rect 237731 3782 237783 3834
rect 237795 3782 237847 3834
rect 44456 3680 44508 3732
rect 48136 3680 48188 3732
rect 67640 3612 67692 3664
rect 37372 3544 37424 3596
rect 38476 3544 38528 3596
rect 23204 3476 23256 3528
rect 36636 3519 36688 3528
rect 36636 3485 36645 3519
rect 36645 3485 36679 3519
rect 36679 3485 36688 3519
rect 36636 3476 36688 3485
rect 36820 3476 36872 3528
rect 7380 3408 7432 3460
rect 23572 3383 23624 3392
rect 23572 3349 23581 3383
rect 23581 3349 23615 3383
rect 23615 3349 23624 3383
rect 23572 3340 23624 3349
rect 36360 3383 36412 3392
rect 36360 3349 36369 3383
rect 36369 3349 36403 3383
rect 36403 3349 36412 3383
rect 36360 3340 36412 3349
rect 37280 3476 37332 3528
rect 41052 3519 41104 3528
rect 41052 3485 41061 3519
rect 41061 3485 41095 3519
rect 41095 3485 41104 3519
rect 41052 3476 41104 3485
rect 41144 3519 41196 3528
rect 41144 3485 41153 3519
rect 41153 3485 41187 3519
rect 41187 3485 41196 3519
rect 41144 3476 41196 3485
rect 41512 3451 41564 3460
rect 41512 3417 41521 3451
rect 41521 3417 41555 3451
rect 41555 3417 41564 3451
rect 41512 3408 41564 3417
rect 37372 3340 37424 3392
rect 39488 3340 39540 3392
rect 41236 3340 41288 3392
rect 41328 3340 41380 3392
rect 42524 3544 42576 3596
rect 43904 3476 43956 3528
rect 43996 3519 44048 3528
rect 43996 3485 44005 3519
rect 44005 3485 44039 3519
rect 44039 3485 44048 3519
rect 43996 3476 44048 3485
rect 43352 3408 43404 3460
rect 43812 3408 43864 3460
rect 45468 3544 45520 3596
rect 47768 3544 47820 3596
rect 47952 3544 48004 3596
rect 51632 3544 51684 3596
rect 92480 3680 92532 3732
rect 92572 3723 92624 3732
rect 92572 3689 92581 3723
rect 92581 3689 92615 3723
rect 92615 3689 92624 3723
rect 92572 3680 92624 3689
rect 92204 3612 92256 3664
rect 94136 3612 94188 3664
rect 94688 3612 94740 3664
rect 48780 3476 48832 3528
rect 48964 3519 49016 3528
rect 48964 3485 48973 3519
rect 48973 3485 49007 3519
rect 49007 3485 49016 3519
rect 48964 3476 49016 3485
rect 50436 3476 50488 3528
rect 50896 3519 50948 3528
rect 50896 3485 50905 3519
rect 50905 3485 50939 3519
rect 50939 3485 50948 3519
rect 50896 3476 50948 3485
rect 48228 3451 48280 3460
rect 48228 3417 48237 3451
rect 48237 3417 48271 3451
rect 48271 3417 48280 3451
rect 48228 3408 48280 3417
rect 48412 3408 48464 3460
rect 48596 3451 48648 3460
rect 48596 3417 48605 3451
rect 48605 3417 48639 3451
rect 48639 3417 48648 3451
rect 48596 3408 48648 3417
rect 42064 3383 42116 3392
rect 42064 3349 42073 3383
rect 42073 3349 42107 3383
rect 42107 3349 42116 3383
rect 42064 3340 42116 3349
rect 43444 3340 43496 3392
rect 44364 3383 44416 3392
rect 44364 3349 44373 3383
rect 44373 3349 44407 3383
rect 44407 3349 44416 3383
rect 44364 3340 44416 3349
rect 51540 3408 51592 3460
rect 94504 3544 94556 3596
rect 94872 3587 94924 3596
rect 94872 3553 94881 3587
rect 94881 3553 94915 3587
rect 94915 3553 94924 3587
rect 94872 3544 94924 3553
rect 95056 3544 95108 3596
rect 95516 3544 95568 3596
rect 91928 3519 91980 3528
rect 91928 3485 91937 3519
rect 91937 3485 91971 3519
rect 91971 3485 91980 3519
rect 91928 3476 91980 3485
rect 49332 3383 49384 3392
rect 49332 3349 49341 3383
rect 49341 3349 49375 3383
rect 49375 3349 49384 3383
rect 49332 3340 49384 3349
rect 49516 3383 49568 3392
rect 49516 3349 49525 3383
rect 49525 3349 49559 3383
rect 49559 3349 49568 3383
rect 49516 3340 49568 3349
rect 50436 3340 50488 3392
rect 51632 3383 51684 3392
rect 51632 3349 51641 3383
rect 51641 3349 51675 3383
rect 51675 3349 51684 3383
rect 51632 3340 51684 3349
rect 51816 3383 51868 3392
rect 51816 3349 51825 3383
rect 51825 3349 51859 3383
rect 51859 3349 51868 3383
rect 51816 3340 51868 3349
rect 52092 3340 52144 3392
rect 92664 3408 92716 3460
rect 93216 3519 93268 3528
rect 93216 3485 93225 3519
rect 93225 3485 93259 3519
rect 93259 3485 93268 3519
rect 93216 3476 93268 3485
rect 93952 3519 94004 3528
rect 93952 3485 93961 3519
rect 93961 3485 93995 3519
rect 93995 3485 94004 3519
rect 93952 3476 94004 3485
rect 94044 3476 94096 3528
rect 96896 3680 96948 3732
rect 96988 3723 97040 3732
rect 96988 3689 96997 3723
rect 96997 3689 97031 3723
rect 97031 3689 97040 3723
rect 96988 3680 97040 3689
rect 101772 3680 101824 3732
rect 101956 3680 102008 3732
rect 105360 3723 105412 3732
rect 105360 3689 105369 3723
rect 105369 3689 105403 3723
rect 105403 3689 105412 3723
rect 105360 3680 105412 3689
rect 106188 3723 106240 3732
rect 106188 3689 106197 3723
rect 106197 3689 106231 3723
rect 106231 3689 106240 3723
rect 106188 3680 106240 3689
rect 106372 3680 106424 3732
rect 108764 3680 108816 3732
rect 95976 3612 96028 3664
rect 97724 3612 97776 3664
rect 100760 3612 100812 3664
rect 104164 3655 104216 3664
rect 104164 3621 104173 3655
rect 104173 3621 104207 3655
rect 104207 3621 104216 3655
rect 104164 3612 104216 3621
rect 105176 3612 105228 3664
rect 99288 3587 99340 3596
rect 99288 3553 99297 3587
rect 99297 3553 99331 3587
rect 99331 3553 99340 3587
rect 99288 3544 99340 3553
rect 101404 3544 101456 3596
rect 103704 3587 103756 3596
rect 103704 3553 103713 3587
rect 103713 3553 103747 3587
rect 103747 3553 103756 3587
rect 103704 3544 103756 3553
rect 104440 3587 104492 3596
rect 104440 3553 104449 3587
rect 104449 3553 104483 3587
rect 104483 3553 104492 3587
rect 104440 3544 104492 3553
rect 104557 3587 104609 3596
rect 104557 3553 104566 3587
rect 104566 3553 104600 3587
rect 104600 3553 104609 3587
rect 104557 3544 104609 3553
rect 105636 3544 105688 3596
rect 96804 3476 96856 3528
rect 96896 3476 96948 3528
rect 97356 3476 97408 3528
rect 101864 3519 101916 3528
rect 101864 3485 101873 3519
rect 101873 3485 101907 3519
rect 101907 3485 101916 3519
rect 101864 3476 101916 3485
rect 102232 3476 102284 3528
rect 93952 3340 94004 3392
rect 99380 3408 99432 3460
rect 100944 3451 100996 3460
rect 100944 3417 100953 3451
rect 100953 3417 100987 3451
rect 100987 3417 100996 3451
rect 100944 3408 100996 3417
rect 103152 3451 103204 3460
rect 103152 3417 103161 3451
rect 103161 3417 103195 3451
rect 103195 3417 103204 3451
rect 105544 3476 105596 3528
rect 106556 3612 106608 3664
rect 111616 3723 111668 3732
rect 111616 3689 111625 3723
rect 111625 3689 111659 3723
rect 111659 3689 111668 3723
rect 111616 3680 111668 3689
rect 111708 3680 111760 3732
rect 117412 3612 117464 3664
rect 118148 3612 118200 3664
rect 118424 3655 118476 3664
rect 118424 3621 118433 3655
rect 118433 3621 118467 3655
rect 118467 3621 118476 3655
rect 118424 3612 118476 3621
rect 121460 3680 121512 3732
rect 122472 3723 122524 3732
rect 122472 3689 122481 3723
rect 122481 3689 122515 3723
rect 122515 3689 122524 3723
rect 122472 3680 122524 3689
rect 140688 3680 140740 3732
rect 120908 3612 120960 3664
rect 106096 3544 106148 3596
rect 108856 3587 108908 3596
rect 108856 3553 108865 3587
rect 108865 3553 108899 3587
rect 108899 3553 108908 3587
rect 108856 3544 108908 3553
rect 109408 3544 109460 3596
rect 110420 3587 110472 3596
rect 110420 3553 110429 3587
rect 110429 3553 110463 3587
rect 110463 3553 110472 3587
rect 110420 3544 110472 3553
rect 110696 3587 110748 3596
rect 110696 3553 110705 3587
rect 110705 3553 110739 3587
rect 110739 3553 110748 3587
rect 110696 3544 110748 3553
rect 111524 3544 111576 3596
rect 111800 3544 111852 3596
rect 112536 3544 112588 3596
rect 113732 3587 113784 3596
rect 113732 3553 113741 3587
rect 113741 3553 113775 3587
rect 113775 3553 113784 3587
rect 113732 3544 113784 3553
rect 114836 3544 114888 3596
rect 117688 3544 117740 3596
rect 118516 3544 118568 3596
rect 119160 3544 119212 3596
rect 120080 3587 120132 3596
rect 120080 3553 120089 3587
rect 120089 3553 120123 3587
rect 120123 3553 120132 3587
rect 120080 3544 120132 3553
rect 122288 3544 122340 3596
rect 106188 3519 106240 3528
rect 106188 3485 106197 3519
rect 106197 3485 106231 3519
rect 106231 3485 106240 3519
rect 106188 3476 106240 3485
rect 106280 3476 106332 3528
rect 103152 3408 103204 3417
rect 105728 3408 105780 3460
rect 110880 3476 110932 3528
rect 114928 3519 114980 3528
rect 114928 3485 114937 3519
rect 114937 3485 114971 3519
rect 114971 3485 114980 3519
rect 114928 3476 114980 3485
rect 117320 3476 117372 3528
rect 117872 3476 117924 3528
rect 118884 3476 118936 3528
rect 118976 3519 119028 3528
rect 118976 3485 118985 3519
rect 118985 3485 119019 3519
rect 119019 3485 119028 3519
rect 118976 3476 119028 3485
rect 122104 3476 122156 3528
rect 123024 3476 123076 3528
rect 112168 3408 112220 3460
rect 98460 3340 98512 3392
rect 103060 3340 103112 3392
rect 103704 3340 103756 3392
rect 107660 3340 107712 3392
rect 110420 3340 110472 3392
rect 111248 3340 111300 3392
rect 119252 3340 119304 3392
rect 139492 3612 139544 3664
rect 142252 3680 142304 3732
rect 145840 3680 145892 3732
rect 149244 3723 149296 3732
rect 149244 3689 149253 3723
rect 149253 3689 149287 3723
rect 149287 3689 149296 3723
rect 149244 3680 149296 3689
rect 144736 3612 144788 3664
rect 145932 3612 145984 3664
rect 148508 3612 148560 3664
rect 151452 3680 151504 3732
rect 150808 3612 150860 3664
rect 152832 3612 152884 3664
rect 153660 3612 153712 3664
rect 154304 3680 154356 3732
rect 155224 3723 155276 3732
rect 155224 3689 155233 3723
rect 155233 3689 155267 3723
rect 155267 3689 155276 3723
rect 155224 3680 155276 3689
rect 156328 3655 156380 3664
rect 156328 3621 156337 3655
rect 156337 3621 156371 3655
rect 156371 3621 156380 3655
rect 156328 3612 156380 3621
rect 149520 3544 149572 3596
rect 152648 3544 152700 3596
rect 153384 3587 153436 3596
rect 153384 3553 153393 3587
rect 153393 3553 153427 3587
rect 153427 3553 153436 3587
rect 153384 3544 153436 3553
rect 153936 3544 153988 3596
rect 154948 3544 155000 3596
rect 155224 3544 155276 3596
rect 156604 3587 156656 3596
rect 156604 3553 156613 3587
rect 156613 3553 156647 3587
rect 156647 3553 156656 3587
rect 156604 3544 156656 3553
rect 138940 3476 138992 3528
rect 139124 3519 139176 3528
rect 139124 3485 139133 3519
rect 139133 3485 139167 3519
rect 139167 3485 139176 3519
rect 139124 3476 139176 3485
rect 139584 3519 139636 3528
rect 139584 3485 139593 3519
rect 139593 3485 139627 3519
rect 139627 3485 139636 3519
rect 139584 3476 139636 3485
rect 141516 3476 141568 3528
rect 141608 3476 141660 3528
rect 141884 3519 141936 3528
rect 141884 3485 141893 3519
rect 141893 3485 141927 3519
rect 141927 3485 141936 3519
rect 141884 3476 141936 3485
rect 139492 3408 139544 3460
rect 141976 3408 142028 3460
rect 142344 3476 142396 3528
rect 142528 3408 142580 3460
rect 143264 3451 143316 3460
rect 143264 3417 143273 3451
rect 143273 3417 143307 3451
rect 143307 3417 143316 3451
rect 143264 3408 143316 3417
rect 143632 3408 143684 3460
rect 144828 3408 144880 3460
rect 138296 3383 138348 3392
rect 138296 3349 138305 3383
rect 138305 3349 138339 3383
rect 138339 3349 138348 3383
rect 138296 3340 138348 3349
rect 139032 3340 139084 3392
rect 145564 3451 145616 3460
rect 145564 3417 145573 3451
rect 145573 3417 145607 3451
rect 145607 3417 145616 3451
rect 145564 3408 145616 3417
rect 145932 3408 145984 3460
rect 149152 3519 149204 3528
rect 149152 3485 149161 3519
rect 149161 3485 149195 3519
rect 149195 3485 149204 3519
rect 149152 3476 149204 3485
rect 149428 3519 149480 3528
rect 149428 3485 149437 3519
rect 149437 3485 149471 3519
rect 149471 3485 149480 3519
rect 149428 3476 149480 3485
rect 152740 3519 152792 3528
rect 152740 3485 152749 3519
rect 152749 3485 152783 3519
rect 152783 3485 152792 3519
rect 152740 3476 152792 3485
rect 153292 3476 153344 3528
rect 154488 3476 154540 3528
rect 154580 3519 154632 3528
rect 154580 3485 154589 3519
rect 154589 3485 154623 3519
rect 154623 3485 154632 3519
rect 154580 3476 154632 3485
rect 155592 3476 155644 3528
rect 156880 3519 156932 3528
rect 156880 3485 156889 3519
rect 156889 3485 156923 3519
rect 156923 3485 156932 3519
rect 156880 3476 156932 3485
rect 147220 3451 147272 3460
rect 147220 3417 147229 3451
rect 147229 3417 147263 3451
rect 147263 3417 147272 3451
rect 147220 3408 147272 3417
rect 149244 3408 149296 3460
rect 149612 3408 149664 3460
rect 150440 3451 150492 3460
rect 150440 3417 150449 3451
rect 150449 3417 150483 3451
rect 150483 3417 150492 3451
rect 150440 3408 150492 3417
rect 151728 3408 151780 3460
rect 160100 3680 160152 3732
rect 172704 3680 172756 3732
rect 207480 3680 207532 3732
rect 211344 3680 211396 3732
rect 159640 3612 159692 3664
rect 182088 3612 182140 3664
rect 208676 3612 208728 3664
rect 159364 3519 159416 3528
rect 159364 3485 159373 3519
rect 159373 3485 159407 3519
rect 159407 3485 159416 3519
rect 159364 3476 159416 3485
rect 168380 3544 168432 3596
rect 171784 3544 171836 3596
rect 189724 3544 189776 3596
rect 207020 3587 207072 3596
rect 207020 3553 207029 3587
rect 207029 3553 207063 3587
rect 207063 3553 207072 3587
rect 207020 3544 207072 3553
rect 207572 3544 207624 3596
rect 207664 3587 207716 3596
rect 207664 3553 207673 3587
rect 207673 3553 207707 3587
rect 207707 3553 207716 3587
rect 207664 3544 207716 3553
rect 209872 3544 209924 3596
rect 212080 3655 212132 3664
rect 212080 3621 212089 3655
rect 212089 3621 212123 3655
rect 212123 3621 212132 3655
rect 212080 3612 212132 3621
rect 168288 3476 168340 3528
rect 207940 3519 207992 3528
rect 207940 3485 207949 3519
rect 207949 3485 207983 3519
rect 207983 3485 207992 3519
rect 207940 3476 207992 3485
rect 208216 3519 208268 3528
rect 208216 3485 208225 3519
rect 208225 3485 208259 3519
rect 208259 3485 208268 3519
rect 208216 3476 208268 3485
rect 210332 3519 210384 3528
rect 210332 3485 210341 3519
rect 210341 3485 210375 3519
rect 210375 3485 210384 3519
rect 210332 3476 210384 3485
rect 210516 3519 210568 3528
rect 210516 3485 210525 3519
rect 210525 3485 210559 3519
rect 210559 3485 210568 3519
rect 210516 3476 210568 3485
rect 210976 3476 211028 3528
rect 211344 3476 211396 3528
rect 211528 3519 211580 3528
rect 211528 3485 211537 3519
rect 211537 3485 211571 3519
rect 211571 3485 211580 3519
rect 211528 3476 211580 3485
rect 211712 3519 211764 3528
rect 211712 3485 211721 3519
rect 211721 3485 211755 3519
rect 211755 3485 211764 3519
rect 211712 3476 211764 3485
rect 213000 3680 213052 3732
rect 218704 3680 218756 3732
rect 224684 3680 224736 3732
rect 214196 3612 214248 3664
rect 215392 3612 215444 3664
rect 216036 3612 216088 3664
rect 217968 3612 218020 3664
rect 218520 3612 218572 3664
rect 219532 3612 219584 3664
rect 219900 3612 219952 3664
rect 221188 3612 221240 3664
rect 227352 3655 227404 3664
rect 227352 3621 227361 3655
rect 227361 3621 227395 3655
rect 227395 3621 227404 3655
rect 227352 3612 227404 3621
rect 227628 3612 227680 3664
rect 228180 3680 228232 3732
rect 243636 3680 243688 3732
rect 245660 3680 245712 3732
rect 246488 3723 246540 3732
rect 246488 3689 246497 3723
rect 246497 3689 246531 3723
rect 246531 3689 246540 3723
rect 246488 3680 246540 3689
rect 246672 3723 246724 3732
rect 246672 3689 246681 3723
rect 246681 3689 246715 3723
rect 246715 3689 246724 3723
rect 246672 3680 246724 3689
rect 247592 3680 247644 3732
rect 251640 3680 251692 3732
rect 252560 3723 252612 3732
rect 252560 3689 252569 3723
rect 252569 3689 252603 3723
rect 252603 3689 252612 3723
rect 252560 3680 252612 3689
rect 252836 3680 252888 3732
rect 254124 3680 254176 3732
rect 257344 3680 257396 3732
rect 258632 3680 258684 3732
rect 259000 3680 259052 3732
rect 264796 3680 264848 3732
rect 267740 3680 267792 3732
rect 268200 3680 268252 3732
rect 268844 3680 268896 3732
rect 269120 3680 269172 3732
rect 270684 3680 270736 3732
rect 161204 3408 161256 3460
rect 187148 3408 187200 3460
rect 209228 3408 209280 3460
rect 210148 3408 210200 3460
rect 146300 3340 146352 3392
rect 152464 3340 152516 3392
rect 153292 3340 153344 3392
rect 155868 3340 155920 3392
rect 156144 3340 156196 3392
rect 158536 3383 158588 3392
rect 158536 3349 158545 3383
rect 158545 3349 158579 3383
rect 158579 3349 158588 3383
rect 158536 3340 158588 3349
rect 158628 3340 158680 3392
rect 167736 3383 167788 3392
rect 167736 3349 167745 3383
rect 167745 3349 167779 3383
rect 167779 3349 167788 3383
rect 167736 3340 167788 3349
rect 206744 3340 206796 3392
rect 207940 3340 207992 3392
rect 209044 3340 209096 3392
rect 212356 3408 212408 3460
rect 213000 3519 213052 3528
rect 213000 3485 213009 3519
rect 213009 3485 213043 3519
rect 213043 3485 213052 3519
rect 213000 3476 213052 3485
rect 214012 3476 214064 3528
rect 215576 3519 215628 3528
rect 215576 3485 215585 3519
rect 215585 3485 215619 3519
rect 215619 3485 215628 3519
rect 215576 3476 215628 3485
rect 216496 3519 216548 3528
rect 216496 3485 216505 3519
rect 216505 3485 216539 3519
rect 216539 3485 216548 3519
rect 216496 3476 216548 3485
rect 217416 3587 217468 3596
rect 217416 3553 217425 3587
rect 217425 3553 217459 3587
rect 217459 3553 217468 3587
rect 217416 3544 217468 3553
rect 221096 3587 221148 3596
rect 221096 3553 221105 3587
rect 221105 3553 221139 3587
rect 221139 3553 221148 3587
rect 221096 3544 221148 3553
rect 221372 3544 221424 3596
rect 216680 3519 216732 3528
rect 216680 3485 216689 3519
rect 216689 3485 216723 3519
rect 216723 3485 216732 3519
rect 216680 3476 216732 3485
rect 211436 3340 211488 3392
rect 211528 3340 211580 3392
rect 215116 3408 215168 3460
rect 217692 3408 217744 3460
rect 222568 3587 222620 3596
rect 222568 3553 222577 3587
rect 222577 3553 222611 3587
rect 222611 3553 222620 3587
rect 222568 3544 222620 3553
rect 222752 3544 222804 3596
rect 223948 3544 224000 3596
rect 224224 3544 224276 3596
rect 225880 3544 225932 3596
rect 226248 3544 226300 3596
rect 229744 3612 229796 3664
rect 229836 3612 229888 3664
rect 241796 3612 241848 3664
rect 244372 3612 244424 3664
rect 223764 3519 223816 3528
rect 223764 3485 223773 3519
rect 223773 3485 223807 3519
rect 223807 3485 223816 3519
rect 223764 3476 223816 3485
rect 224040 3476 224092 3528
rect 225512 3519 225564 3528
rect 225512 3485 225521 3519
rect 225521 3485 225555 3519
rect 225555 3485 225564 3519
rect 225512 3476 225564 3485
rect 225696 3519 225748 3528
rect 225696 3485 225705 3519
rect 225705 3485 225739 3519
rect 225739 3485 225748 3519
rect 225696 3476 225748 3485
rect 226708 3519 226760 3528
rect 226708 3485 226717 3519
rect 226717 3485 226751 3519
rect 226751 3485 226760 3519
rect 226708 3476 226760 3485
rect 219164 3408 219216 3460
rect 219624 3408 219676 3460
rect 220820 3408 220872 3460
rect 220912 3408 220964 3460
rect 221464 3408 221516 3460
rect 231860 3544 231912 3596
rect 227720 3476 227772 3528
rect 238760 3544 238812 3596
rect 236276 3476 236328 3528
rect 244004 3544 244056 3596
rect 244556 3544 244608 3596
rect 246856 3544 246908 3596
rect 247316 3587 247368 3596
rect 247316 3553 247325 3587
rect 247325 3553 247359 3587
rect 247359 3553 247368 3587
rect 247316 3544 247368 3553
rect 249248 3544 249300 3596
rect 253296 3612 253348 3664
rect 251640 3544 251692 3596
rect 254032 3587 254084 3596
rect 254032 3553 254041 3587
rect 254041 3553 254075 3587
rect 254075 3553 254084 3587
rect 254032 3544 254084 3553
rect 255136 3544 255188 3596
rect 268016 3612 268068 3664
rect 213736 3383 213788 3392
rect 213736 3349 213745 3383
rect 213745 3349 213779 3383
rect 213779 3349 213788 3383
rect 213736 3340 213788 3349
rect 216588 3340 216640 3392
rect 222108 3340 222160 3392
rect 223948 3340 224000 3392
rect 244004 3408 244056 3460
rect 244280 3408 244332 3460
rect 246948 3476 247000 3528
rect 247040 3519 247092 3528
rect 247040 3485 247049 3519
rect 247049 3485 247083 3519
rect 247083 3485 247092 3519
rect 247040 3476 247092 3485
rect 250996 3476 251048 3528
rect 251364 3476 251416 3528
rect 258724 3544 258776 3596
rect 259368 3476 259420 3528
rect 260656 3476 260708 3528
rect 265900 3544 265952 3596
rect 266544 3544 266596 3596
rect 225880 3340 225932 3392
rect 227720 3383 227772 3392
rect 227720 3349 227729 3383
rect 227729 3349 227763 3383
rect 227763 3349 227772 3383
rect 227720 3340 227772 3349
rect 229744 3340 229796 3392
rect 245016 3408 245068 3460
rect 244648 3383 244700 3392
rect 244648 3349 244657 3383
rect 244657 3349 244691 3383
rect 244691 3349 244700 3383
rect 244648 3340 244700 3349
rect 244832 3340 244884 3392
rect 246580 3408 246632 3460
rect 247224 3408 247276 3460
rect 248144 3451 248196 3460
rect 248144 3417 248153 3451
rect 248153 3417 248187 3451
rect 248187 3417 248196 3451
rect 248144 3408 248196 3417
rect 245568 3383 245620 3392
rect 245568 3349 245577 3383
rect 245577 3349 245611 3383
rect 245611 3349 245620 3383
rect 245568 3340 245620 3349
rect 248420 3340 248472 3392
rect 249616 3340 249668 3392
rect 252652 3408 252704 3460
rect 253940 3408 253992 3460
rect 254308 3408 254360 3460
rect 259276 3408 259328 3460
rect 259736 3451 259788 3460
rect 259736 3417 259745 3451
rect 259745 3417 259779 3451
rect 259779 3417 259788 3451
rect 259736 3408 259788 3417
rect 267464 3519 267516 3528
rect 267464 3485 267473 3519
rect 267473 3485 267507 3519
rect 267507 3485 267516 3519
rect 267464 3476 267516 3485
rect 268108 3519 268160 3528
rect 268108 3485 268117 3519
rect 268117 3485 268151 3519
rect 268151 3485 268160 3519
rect 268108 3476 268160 3485
rect 268752 3519 268804 3528
rect 268752 3485 268761 3519
rect 268761 3485 268795 3519
rect 268795 3485 268804 3519
rect 268752 3476 268804 3485
rect 270776 3612 270828 3664
rect 271788 3612 271840 3664
rect 270592 3476 270644 3528
rect 271880 3476 271932 3528
rect 254124 3340 254176 3392
rect 258908 3340 258960 3392
rect 260472 3340 260524 3392
rect 262128 3340 262180 3392
rect 267924 3408 267976 3460
rect 267740 3340 267792 3392
rect 268936 3340 268988 3392
rect 271236 3408 271288 3460
rect 271144 3340 271196 3392
rect 272156 3340 272208 3392
rect 68546 3238 68598 3290
rect 68610 3238 68662 3290
rect 68674 3238 68726 3290
rect 68738 3238 68790 3290
rect 68802 3238 68854 3290
rect 136143 3238 136195 3290
rect 136207 3238 136259 3290
rect 136271 3238 136323 3290
rect 136335 3238 136387 3290
rect 136399 3238 136451 3290
rect 203740 3238 203792 3290
rect 203804 3238 203856 3290
rect 203868 3238 203920 3290
rect 203932 3238 203984 3290
rect 203996 3238 204048 3290
rect 271337 3238 271389 3290
rect 271401 3238 271453 3290
rect 271465 3238 271517 3290
rect 271529 3238 271581 3290
rect 271593 3238 271645 3290
rect 23480 3136 23532 3188
rect 39120 3136 39172 3188
rect 39488 3136 39540 3188
rect 42432 3136 42484 3188
rect 24952 3068 25004 3120
rect 22100 3000 22152 3052
rect 23296 3000 23348 3052
rect 23664 3043 23716 3052
rect 23664 3009 23673 3043
rect 23673 3009 23707 3043
rect 23707 3009 23716 3043
rect 23664 3000 23716 3009
rect 24492 3043 24544 3052
rect 24492 3009 24501 3043
rect 24501 3009 24535 3043
rect 24535 3009 24544 3043
rect 24492 3000 24544 3009
rect 24584 3043 24636 3052
rect 24584 3009 24593 3043
rect 24593 3009 24627 3043
rect 24627 3009 24636 3043
rect 24584 3000 24636 3009
rect 25412 3000 25464 3052
rect 26240 3000 26292 3052
rect 37648 3111 37700 3120
rect 37648 3077 37657 3111
rect 37657 3077 37691 3111
rect 37691 3077 37700 3111
rect 37648 3068 37700 3077
rect 37924 3111 37976 3120
rect 37924 3077 37933 3111
rect 37933 3077 37967 3111
rect 37967 3077 37976 3111
rect 37924 3068 37976 3077
rect 38016 3111 38068 3120
rect 38016 3077 38025 3111
rect 38025 3077 38059 3111
rect 38059 3077 38068 3111
rect 38016 3068 38068 3077
rect 39212 3068 39264 3120
rect 38568 3000 38620 3052
rect 43168 3068 43220 3120
rect 43260 3111 43312 3120
rect 43260 3077 43269 3111
rect 43269 3077 43303 3111
rect 43303 3077 43312 3111
rect 43260 3068 43312 3077
rect 43352 3111 43404 3120
rect 43352 3077 43361 3111
rect 43361 3077 43395 3111
rect 43395 3077 43404 3111
rect 43352 3068 43404 3077
rect 44088 3179 44140 3188
rect 44088 3145 44097 3179
rect 44097 3145 44131 3179
rect 44131 3145 44140 3179
rect 44088 3136 44140 3145
rect 47492 3136 47544 3188
rect 49516 3136 49568 3188
rect 93032 3136 93084 3188
rect 93308 3136 93360 3188
rect 47952 3111 48004 3120
rect 47952 3077 47961 3111
rect 47961 3077 47995 3111
rect 47995 3077 48004 3111
rect 47952 3068 48004 3077
rect 49056 3111 49108 3120
rect 49056 3077 49065 3111
rect 49065 3077 49099 3111
rect 49099 3077 49108 3111
rect 49056 3068 49108 3077
rect 51816 3068 51868 3120
rect 91192 3068 91244 3120
rect 31944 2932 31996 2984
rect 38476 2932 38528 2984
rect 40592 2932 40644 2984
rect 41144 2932 41196 2984
rect 43812 2932 43864 2984
rect 48044 3000 48096 3052
rect 48504 3000 48556 3052
rect 48688 3043 48740 3052
rect 48688 3009 48697 3043
rect 48697 3009 48731 3043
rect 48731 3009 48740 3043
rect 48688 3000 48740 3009
rect 49148 3000 49200 3052
rect 54668 3000 54720 3052
rect 89352 3043 89404 3052
rect 89352 3009 89361 3043
rect 89361 3009 89395 3043
rect 89395 3009 89404 3043
rect 89352 3000 89404 3009
rect 90916 3000 90968 3052
rect 91836 3043 91888 3052
rect 91836 3009 91845 3043
rect 91845 3009 91879 3043
rect 91879 3009 91888 3043
rect 91836 3000 91888 3009
rect 96436 3179 96488 3188
rect 96436 3145 96445 3179
rect 96445 3145 96479 3179
rect 96479 3145 96488 3179
rect 96436 3136 96488 3145
rect 96528 3136 96580 3188
rect 97264 3136 97316 3188
rect 97632 3136 97684 3188
rect 97908 3136 97960 3188
rect 47676 2932 47728 2984
rect 47768 2932 47820 2984
rect 66352 2975 66404 2984
rect 66352 2941 66361 2975
rect 66361 2941 66395 2975
rect 66395 2941 66404 2975
rect 66352 2932 66404 2941
rect 94136 3043 94188 3052
rect 94136 3009 94145 3043
rect 94145 3009 94179 3043
rect 94179 3009 94188 3043
rect 94136 3000 94188 3009
rect 94320 3000 94372 3052
rect 94504 3000 94556 3052
rect 94964 3043 95016 3052
rect 94964 3009 94973 3043
rect 94973 3009 95007 3043
rect 95007 3009 95016 3043
rect 94964 3000 95016 3009
rect 96344 3000 96396 3052
rect 93400 2932 93452 2984
rect 96160 2932 96212 2984
rect 19248 2864 19300 2916
rect 25964 2864 26016 2916
rect 44180 2864 44232 2916
rect 49240 2907 49292 2916
rect 49240 2873 49249 2907
rect 49249 2873 49283 2907
rect 49283 2873 49292 2907
rect 49240 2864 49292 2873
rect 95424 2864 95476 2916
rect 95700 2864 95752 2916
rect 96436 2864 96488 2916
rect 96620 3000 96672 3052
rect 99748 3111 99800 3120
rect 99748 3077 99757 3111
rect 99757 3077 99791 3111
rect 99791 3077 99800 3111
rect 99748 3068 99800 3077
rect 101588 3068 101640 3120
rect 103704 3111 103756 3120
rect 103704 3077 103713 3111
rect 103713 3077 103747 3111
rect 103747 3077 103756 3111
rect 103704 3068 103756 3077
rect 103612 3000 103664 3052
rect 104992 3136 105044 3188
rect 106188 3136 106240 3188
rect 106280 3179 106332 3188
rect 106280 3145 106289 3179
rect 106289 3145 106323 3179
rect 106323 3145 106332 3179
rect 106280 3136 106332 3145
rect 105360 3043 105412 3052
rect 105360 3009 105369 3043
rect 105369 3009 105403 3043
rect 105403 3009 105412 3043
rect 105360 3000 105412 3009
rect 105636 3043 105688 3052
rect 105636 3009 105645 3043
rect 105645 3009 105679 3043
rect 105679 3009 105688 3043
rect 105636 3000 105688 3009
rect 99012 2932 99064 2984
rect 99380 2864 99432 2916
rect 101496 2932 101548 2984
rect 105452 2975 105504 2984
rect 105452 2941 105486 2975
rect 105486 2941 105504 2975
rect 113364 3136 113416 3188
rect 147220 3136 147272 3188
rect 105452 2932 105504 2941
rect 104992 2864 105044 2916
rect 105176 2864 105228 2916
rect 22100 2796 22152 2848
rect 23848 2839 23900 2848
rect 23848 2805 23857 2839
rect 23857 2805 23891 2839
rect 23891 2805 23900 2839
rect 23848 2796 23900 2805
rect 24400 2796 24452 2848
rect 25780 2839 25832 2848
rect 25780 2805 25789 2839
rect 25789 2805 25823 2839
rect 25823 2805 25832 2839
rect 25780 2796 25832 2805
rect 26516 2839 26568 2848
rect 26516 2805 26525 2839
rect 26525 2805 26559 2839
rect 26559 2805 26568 2839
rect 26516 2796 26568 2805
rect 54484 2839 54536 2848
rect 54484 2805 54493 2839
rect 54493 2805 54527 2839
rect 54527 2805 54536 2839
rect 54484 2796 54536 2805
rect 89536 2839 89588 2848
rect 89536 2805 89545 2839
rect 89545 2805 89579 2839
rect 89579 2805 89588 2839
rect 89536 2796 89588 2805
rect 90824 2839 90876 2848
rect 90824 2805 90833 2839
rect 90833 2805 90867 2839
rect 90867 2805 90876 2839
rect 90824 2796 90876 2805
rect 92020 2839 92072 2848
rect 92020 2805 92029 2839
rect 92029 2805 92063 2839
rect 92063 2805 92072 2839
rect 92020 2796 92072 2805
rect 92756 2839 92808 2848
rect 92756 2805 92765 2839
rect 92765 2805 92799 2839
rect 92799 2805 92808 2839
rect 92756 2796 92808 2805
rect 96988 2796 97040 2848
rect 97356 2796 97408 2848
rect 104348 2796 104400 2848
rect 104716 2796 104768 2848
rect 106464 2932 106516 2984
rect 108948 2975 109000 2984
rect 108948 2941 108957 2975
rect 108957 2941 108991 2975
rect 108991 2941 109000 2975
rect 108948 2932 109000 2941
rect 106372 2864 106424 2916
rect 106188 2796 106240 2848
rect 110236 3043 110288 3052
rect 110236 3009 110245 3043
rect 110245 3009 110279 3043
rect 110279 3009 110288 3043
rect 110236 3000 110288 3009
rect 110512 2975 110564 2984
rect 110512 2941 110521 2975
rect 110521 2941 110555 2975
rect 110555 2941 110564 2975
rect 110512 2932 110564 2941
rect 110420 2864 110472 2916
rect 115020 3043 115072 3052
rect 115020 3009 115029 3043
rect 115029 3009 115063 3043
rect 115063 3009 115072 3043
rect 115020 3000 115072 3009
rect 119252 3000 119304 3052
rect 119988 3043 120040 3052
rect 119988 3009 119997 3043
rect 119997 3009 120031 3043
rect 120031 3009 120040 3043
rect 119988 3000 120040 3009
rect 111616 2932 111668 2984
rect 109592 2839 109644 2848
rect 109592 2805 109601 2839
rect 109601 2805 109635 2839
rect 109635 2805 109644 2839
rect 109592 2796 109644 2805
rect 111708 2864 111760 2916
rect 113456 2975 113508 2984
rect 113456 2941 113465 2975
rect 113465 2941 113499 2975
rect 113499 2941 113508 2975
rect 113456 2932 113508 2941
rect 115204 2975 115256 2984
rect 115204 2941 115213 2975
rect 115213 2941 115247 2975
rect 115247 2941 115256 2975
rect 115204 2932 115256 2941
rect 117504 2975 117556 2984
rect 117504 2941 117513 2975
rect 117513 2941 117547 2975
rect 117547 2941 117556 2975
rect 117504 2932 117556 2941
rect 118608 2932 118660 2984
rect 118976 2932 119028 2984
rect 120724 2975 120776 2984
rect 120724 2941 120733 2975
rect 120733 2941 120767 2975
rect 120767 2941 120776 2975
rect 120724 2932 120776 2941
rect 121644 2932 121696 2984
rect 121736 2864 121788 2916
rect 135352 2975 135404 2984
rect 135352 2941 135361 2975
rect 135361 2941 135395 2975
rect 135395 2941 135404 2975
rect 135352 2932 135404 2941
rect 138296 3068 138348 3120
rect 140872 3068 140924 3120
rect 145656 3068 145708 3120
rect 138940 3000 138992 3052
rect 139032 3043 139084 3052
rect 139032 3009 139041 3043
rect 139041 3009 139075 3043
rect 139075 3009 139084 3043
rect 139032 3000 139084 3009
rect 139676 3043 139728 3052
rect 139676 3009 139685 3043
rect 139685 3009 139719 3043
rect 139719 3009 139728 3043
rect 139676 3000 139728 3009
rect 148232 3000 148284 3052
rect 149336 3043 149388 3052
rect 149336 3009 149345 3043
rect 149345 3009 149379 3043
rect 149379 3009 149388 3043
rect 149336 3000 149388 3009
rect 149612 3043 149664 3052
rect 149612 3009 149621 3043
rect 149621 3009 149655 3043
rect 149655 3009 149664 3043
rect 149612 3000 149664 3009
rect 139952 2932 140004 2984
rect 141148 2932 141200 2984
rect 142068 2975 142120 2984
rect 142068 2941 142077 2975
rect 142077 2941 142111 2975
rect 142111 2941 142120 2975
rect 142068 2932 142120 2941
rect 139492 2907 139544 2916
rect 139492 2873 139501 2907
rect 139501 2873 139535 2907
rect 139535 2873 139544 2907
rect 139492 2864 139544 2873
rect 143540 2975 143592 2984
rect 143540 2941 143549 2975
rect 143549 2941 143583 2975
rect 143583 2941 143592 2975
rect 143540 2932 143592 2941
rect 144552 2932 144604 2984
rect 144644 2864 144696 2916
rect 146484 2975 146536 2984
rect 146484 2941 146493 2975
rect 146493 2941 146527 2975
rect 146527 2941 146536 2975
rect 146484 2932 146536 2941
rect 149152 2932 149204 2984
rect 150440 3136 150492 3188
rect 156236 3136 156288 3188
rect 160284 3136 160336 3188
rect 171784 3136 171836 3188
rect 152464 3068 152516 3120
rect 152556 3000 152608 3052
rect 155040 3068 155092 3120
rect 159364 3068 159416 3120
rect 209688 3136 209740 3188
rect 209780 3136 209832 3188
rect 210976 3136 211028 3188
rect 211620 3136 211672 3188
rect 213000 3136 213052 3188
rect 213460 3136 213512 3188
rect 213828 3136 213880 3188
rect 218796 3136 218848 3188
rect 154672 3000 154724 3052
rect 147404 2864 147456 2916
rect 148508 2864 148560 2916
rect 151268 2932 151320 2984
rect 152832 2932 152884 2984
rect 153660 2932 153712 2984
rect 156144 3043 156196 3052
rect 156144 3009 156153 3043
rect 156153 3009 156187 3043
rect 156187 3009 156196 3043
rect 156144 3000 156196 3009
rect 159088 3000 159140 3052
rect 160284 3000 160336 3052
rect 155776 2932 155828 2984
rect 156420 2932 156472 2984
rect 206652 3068 206704 3120
rect 165712 3000 165764 3052
rect 170312 3000 170364 3052
rect 191288 3000 191340 3052
rect 206560 3000 206612 3052
rect 208860 3068 208912 3120
rect 211988 3068 212040 3120
rect 215116 3111 215168 3120
rect 215116 3077 215125 3111
rect 215125 3077 215159 3111
rect 215159 3077 215168 3111
rect 215116 3068 215168 3077
rect 216772 3068 216824 3120
rect 218428 3068 218480 3120
rect 220912 3179 220964 3188
rect 220912 3145 220921 3179
rect 220921 3145 220955 3179
rect 220955 3145 220964 3179
rect 220912 3136 220964 3145
rect 167920 2975 167972 2984
rect 167920 2941 167929 2975
rect 167929 2941 167963 2975
rect 167963 2941 167972 2975
rect 167920 2932 167972 2941
rect 203156 2975 203208 2984
rect 203156 2941 203165 2975
rect 203165 2941 203199 2975
rect 203199 2941 203208 2975
rect 203156 2932 203208 2941
rect 207940 3043 207992 3052
rect 207940 3009 207949 3043
rect 207949 3009 207983 3043
rect 207983 3009 207992 3043
rect 207940 3000 207992 3009
rect 208768 3000 208820 3052
rect 209964 3043 210016 3052
rect 209964 3009 209998 3043
rect 209998 3009 210016 3043
rect 209964 3000 210016 3009
rect 210148 3043 210200 3052
rect 210148 3009 210157 3043
rect 210157 3009 210191 3043
rect 210191 3009 210200 3043
rect 210148 3000 210200 3009
rect 211344 3043 211396 3052
rect 211344 3009 211353 3043
rect 211353 3009 211387 3043
rect 211387 3009 211396 3043
rect 211344 3000 211396 3009
rect 211436 3043 211488 3052
rect 211436 3009 211445 3043
rect 211445 3009 211479 3043
rect 211479 3009 211488 3043
rect 211436 3000 211488 3009
rect 211620 3043 211672 3052
rect 211620 3009 211629 3043
rect 211629 3009 211663 3043
rect 211663 3009 211672 3043
rect 211620 3000 211672 3009
rect 212356 3000 212408 3052
rect 212540 3000 212592 3052
rect 208676 2932 208728 2984
rect 209136 2975 209188 2984
rect 209136 2941 209145 2975
rect 209145 2941 209179 2975
rect 209179 2941 209188 2975
rect 209136 2932 209188 2941
rect 116124 2796 116176 2848
rect 120080 2796 120132 2848
rect 138204 2839 138256 2848
rect 138204 2805 138213 2839
rect 138213 2805 138247 2839
rect 138247 2805 138256 2839
rect 138204 2796 138256 2805
rect 143264 2796 143316 2848
rect 145472 2796 145524 2848
rect 150348 2796 150400 2848
rect 152924 2796 152976 2848
rect 153016 2796 153068 2848
rect 206192 2864 206244 2916
rect 208308 2907 208360 2916
rect 208308 2873 208317 2907
rect 208317 2873 208351 2907
rect 208351 2873 208360 2907
rect 208308 2864 208360 2873
rect 209596 2907 209648 2916
rect 155132 2796 155184 2848
rect 156236 2796 156288 2848
rect 158444 2796 158496 2848
rect 158628 2839 158680 2848
rect 158628 2805 158637 2839
rect 158637 2805 158671 2839
rect 158671 2805 158680 2839
rect 158628 2796 158680 2805
rect 159364 2839 159416 2848
rect 159364 2805 159373 2839
rect 159373 2805 159407 2839
rect 159407 2805 159416 2839
rect 159364 2796 159416 2805
rect 191104 2839 191156 2848
rect 191104 2805 191113 2839
rect 191113 2805 191147 2839
rect 191147 2805 191156 2839
rect 191104 2796 191156 2805
rect 207664 2796 207716 2848
rect 209596 2873 209605 2907
rect 209605 2873 209639 2907
rect 209639 2873 209648 2907
rect 209596 2864 209648 2873
rect 211160 2864 211212 2916
rect 213000 2932 213052 2984
rect 213828 2932 213880 2984
rect 214288 2975 214340 2984
rect 214288 2941 214297 2975
rect 214297 2941 214331 2975
rect 214331 2941 214340 2975
rect 214288 2932 214340 2941
rect 214932 2975 214984 2984
rect 214932 2941 214941 2975
rect 214941 2941 214975 2975
rect 214975 2941 214984 2975
rect 214932 2932 214984 2941
rect 215392 2975 215444 2984
rect 215392 2941 215401 2975
rect 215401 2941 215435 2975
rect 215435 2941 215444 2975
rect 215392 2932 215444 2941
rect 209964 2796 210016 2848
rect 216680 2864 216732 2916
rect 218336 2975 218388 2984
rect 218336 2941 218345 2975
rect 218345 2941 218379 2975
rect 218379 2941 218388 2975
rect 218336 2932 218388 2941
rect 218428 2932 218480 2984
rect 219348 2932 219400 2984
rect 219624 2975 219676 2984
rect 219624 2941 219633 2975
rect 219633 2941 219667 2975
rect 219667 2941 219676 2975
rect 219624 2932 219676 2941
rect 220636 3043 220688 3052
rect 220636 3009 220645 3043
rect 220645 3009 220679 3043
rect 220679 3009 220688 3043
rect 220636 3000 220688 3009
rect 221372 3000 221424 3052
rect 221648 3043 221700 3052
rect 221648 3009 221657 3043
rect 221657 3009 221691 3043
rect 221691 3009 221700 3043
rect 221648 3000 221700 3009
rect 221832 3043 221884 3052
rect 221832 3009 221841 3043
rect 221841 3009 221875 3043
rect 221875 3009 221884 3043
rect 221832 3000 221884 3009
rect 223396 3043 223448 3052
rect 223396 3009 223405 3043
rect 223405 3009 223439 3043
rect 223439 3009 223448 3043
rect 223396 3000 223448 3009
rect 225236 3111 225288 3120
rect 225236 3077 225245 3111
rect 225245 3077 225279 3111
rect 225279 3077 225288 3111
rect 225236 3068 225288 3077
rect 225696 3179 225748 3188
rect 225696 3145 225705 3179
rect 225705 3145 225739 3179
rect 225739 3145 225748 3179
rect 225696 3136 225748 3145
rect 225788 3136 225840 3188
rect 227444 3136 227496 3188
rect 227996 3136 228048 3188
rect 228364 3136 228416 3188
rect 244372 3136 244424 3188
rect 244924 3136 244976 3188
rect 245016 3136 245068 3188
rect 244004 3111 244056 3120
rect 244004 3077 244013 3111
rect 244013 3077 244047 3111
rect 244047 3077 244056 3111
rect 244004 3068 244056 3077
rect 244832 3068 244884 3120
rect 245108 3111 245160 3120
rect 245108 3077 245117 3111
rect 245117 3077 245151 3111
rect 245151 3077 245160 3111
rect 245108 3068 245160 3077
rect 248604 3068 248656 3120
rect 264244 3136 264296 3188
rect 267280 3179 267332 3188
rect 267280 3145 267289 3179
rect 267289 3145 267323 3179
rect 267323 3145 267332 3179
rect 267280 3136 267332 3145
rect 267832 3136 267884 3188
rect 269580 3136 269632 3188
rect 223764 3000 223816 3052
rect 224316 3043 224368 3052
rect 224316 3009 224325 3043
rect 224325 3009 224359 3043
rect 224359 3009 224368 3043
rect 224316 3000 224368 3009
rect 224592 3043 224644 3052
rect 224592 3009 224601 3043
rect 224601 3009 224635 3043
rect 224635 3009 224644 3043
rect 224592 3000 224644 3009
rect 225880 3043 225932 3052
rect 225880 3009 225889 3043
rect 225889 3009 225923 3043
rect 225923 3009 225932 3043
rect 225880 3000 225932 3009
rect 225972 3000 226024 3052
rect 227720 3000 227772 3052
rect 243360 3000 243412 3052
rect 244280 3043 244332 3052
rect 244280 3009 244289 3043
rect 244289 3009 244323 3043
rect 244323 3009 244332 3043
rect 244280 3000 244332 3009
rect 248420 3000 248472 3052
rect 248696 3043 248748 3052
rect 248696 3009 248705 3043
rect 248705 3009 248739 3043
rect 248739 3009 248748 3043
rect 248696 3000 248748 3009
rect 250076 3000 250128 3052
rect 220820 2932 220872 2984
rect 219256 2864 219308 2916
rect 220544 2864 220596 2916
rect 221372 2864 221424 2916
rect 213000 2796 213052 2848
rect 216496 2796 216548 2848
rect 217876 2796 217928 2848
rect 220636 2796 220688 2848
rect 221556 2839 221608 2848
rect 221556 2805 221565 2839
rect 221565 2805 221599 2839
rect 221599 2805 221608 2839
rect 221556 2796 221608 2805
rect 221648 2796 221700 2848
rect 222752 2796 222804 2848
rect 223672 2932 223724 2984
rect 224132 2932 224184 2984
rect 235816 2932 235868 2984
rect 229744 2864 229796 2916
rect 244372 2932 244424 2984
rect 246856 2932 246908 2984
rect 247408 2932 247460 2984
rect 250536 2975 250588 2984
rect 250536 2941 250545 2975
rect 250545 2941 250579 2975
rect 250579 2941 250588 2975
rect 250536 2932 250588 2941
rect 251180 2975 251232 2984
rect 251180 2941 251189 2975
rect 251189 2941 251223 2975
rect 251223 2941 251232 2975
rect 251180 2932 251232 2941
rect 244556 2864 244608 2916
rect 244648 2864 244700 2916
rect 256516 3000 256568 3052
rect 268016 3068 268068 3120
rect 253848 2975 253900 2984
rect 253848 2941 253857 2975
rect 253857 2941 253891 2975
rect 253891 2941 253900 2975
rect 253848 2932 253900 2941
rect 245660 2796 245712 2848
rect 246304 2796 246356 2848
rect 258172 2932 258224 2984
rect 260012 3000 260064 3052
rect 260472 3043 260524 3052
rect 260472 3009 260481 3043
rect 260481 3009 260515 3043
rect 260515 3009 260524 3043
rect 260472 3000 260524 3009
rect 261024 3000 261076 3052
rect 261116 3043 261168 3052
rect 261116 3009 261125 3043
rect 261125 3009 261159 3043
rect 261159 3009 261168 3043
rect 261116 3000 261168 3009
rect 260288 2975 260340 2984
rect 260288 2941 260297 2975
rect 260297 2941 260331 2975
rect 260331 2941 260340 2975
rect 260288 2932 260340 2941
rect 260564 2932 260616 2984
rect 267740 3000 267792 3052
rect 268660 3068 268712 3120
rect 269028 3000 269080 3052
rect 269856 3043 269908 3052
rect 269856 3009 269865 3043
rect 269865 3009 269899 3043
rect 269899 3009 269908 3043
rect 269856 3000 269908 3009
rect 270960 3043 271012 3052
rect 270960 3009 270969 3043
rect 270969 3009 271003 3043
rect 271003 3009 271012 3043
rect 270960 3000 271012 3009
rect 268660 2932 268712 2984
rect 258816 2864 258868 2916
rect 260472 2864 260524 2916
rect 266820 2864 266872 2916
rect 267556 2864 267608 2916
rect 258264 2796 258316 2848
rect 259092 2796 259144 2848
rect 259828 2796 259880 2848
rect 267648 2796 267700 2848
rect 267924 2839 267976 2848
rect 267924 2805 267933 2839
rect 267933 2805 267967 2839
rect 267967 2805 267976 2839
rect 267924 2796 267976 2805
rect 270684 2796 270736 2848
rect 34748 2694 34800 2746
rect 34812 2694 34864 2746
rect 34876 2694 34928 2746
rect 34940 2694 34992 2746
rect 35004 2694 35056 2746
rect 102345 2694 102397 2746
rect 102409 2694 102461 2746
rect 102473 2694 102525 2746
rect 102537 2694 102589 2746
rect 102601 2694 102653 2746
rect 169942 2694 169994 2746
rect 170006 2694 170058 2746
rect 170070 2694 170122 2746
rect 170134 2694 170186 2746
rect 170198 2694 170250 2746
rect 237539 2694 237591 2746
rect 237603 2694 237655 2746
rect 237667 2694 237719 2746
rect 237731 2694 237783 2746
rect 237795 2694 237847 2746
rect 848 2592 900 2644
rect 22836 2592 22888 2644
rect 23664 2592 23716 2644
rect 25044 2592 25096 2644
rect 27620 2635 27672 2644
rect 27620 2601 27629 2635
rect 27629 2601 27663 2635
rect 27663 2601 27672 2635
rect 27620 2592 27672 2601
rect 43536 2635 43588 2644
rect 43536 2601 43545 2635
rect 43545 2601 43579 2635
rect 43579 2601 43588 2635
rect 43536 2592 43588 2601
rect 47492 2592 47544 2644
rect 51816 2592 51868 2644
rect 55220 2592 55272 2644
rect 1860 2524 1912 2576
rect 21272 2524 21324 2576
rect 4804 2499 4856 2508
rect 4804 2465 4813 2499
rect 4813 2465 4847 2499
rect 4847 2465 4856 2499
rect 4804 2456 4856 2465
rect 5540 2456 5592 2508
rect 23480 2524 23532 2576
rect 24308 2524 24360 2576
rect 24768 2524 24820 2576
rect 22468 2456 22520 2508
rect 23388 2499 23440 2508
rect 23388 2465 23397 2499
rect 23397 2465 23431 2499
rect 23431 2465 23440 2499
rect 23388 2456 23440 2465
rect 4528 2431 4580 2440
rect 4528 2397 4537 2431
rect 4537 2397 4571 2431
rect 4571 2397 4580 2431
rect 4528 2388 4580 2397
rect 6736 2431 6788 2440
rect 6736 2397 6745 2431
rect 6745 2397 6779 2431
rect 6779 2397 6788 2431
rect 6736 2388 6788 2397
rect 7012 2431 7064 2440
rect 7012 2397 7021 2431
rect 7021 2397 7055 2431
rect 7055 2397 7064 2431
rect 7012 2388 7064 2397
rect 14832 2431 14884 2440
rect 14832 2397 14841 2431
rect 14841 2397 14875 2431
rect 14875 2397 14884 2431
rect 14832 2388 14884 2397
rect 15108 2431 15160 2440
rect 15108 2397 15117 2431
rect 15117 2397 15151 2431
rect 15151 2397 15160 2431
rect 15108 2388 15160 2397
rect 22100 2388 22152 2440
rect 22284 2388 22336 2440
rect 23296 2388 23348 2440
rect 24400 2431 24452 2440
rect 24400 2397 24409 2431
rect 24409 2397 24443 2431
rect 24443 2397 24452 2431
rect 24400 2388 24452 2397
rect 24584 2388 24636 2440
rect 26056 2456 26108 2508
rect 38476 2456 38528 2508
rect 26332 2388 26384 2440
rect 27436 2431 27488 2440
rect 27436 2397 27445 2431
rect 27445 2397 27479 2431
rect 27479 2397 27488 2431
rect 27436 2388 27488 2397
rect 29736 2431 29788 2440
rect 29736 2397 29745 2431
rect 29745 2397 29779 2431
rect 29779 2397 29788 2431
rect 29736 2388 29788 2397
rect 31944 2431 31996 2440
rect 31944 2397 31953 2431
rect 31953 2397 31987 2431
rect 31987 2397 31996 2431
rect 31944 2388 31996 2397
rect 32772 2431 32824 2440
rect 32772 2397 32781 2431
rect 32781 2397 32815 2431
rect 32815 2397 32824 2431
rect 32772 2388 32824 2397
rect 38200 2388 38252 2440
rect 32496 2320 32548 2372
rect 38016 2320 38068 2372
rect 38476 2363 38528 2372
rect 38476 2329 38485 2363
rect 38485 2329 38519 2363
rect 38519 2329 38528 2363
rect 38476 2320 38528 2329
rect 38936 2388 38988 2440
rect 40132 2388 40184 2440
rect 40500 2431 40552 2440
rect 40500 2397 40509 2431
rect 40509 2397 40543 2431
rect 40543 2397 40552 2431
rect 40500 2388 40552 2397
rect 40960 2431 41012 2440
rect 40960 2397 40969 2431
rect 40969 2397 41003 2431
rect 41003 2397 41012 2431
rect 40960 2388 41012 2397
rect 41052 2388 41104 2440
rect 41328 2456 41380 2508
rect 43996 2456 44048 2508
rect 42892 2388 42944 2440
rect 42984 2431 43036 2440
rect 42984 2397 42993 2431
rect 42993 2397 43027 2431
rect 43027 2397 43036 2431
rect 42984 2388 43036 2397
rect 40592 2363 40644 2372
rect 40592 2329 40601 2363
rect 40601 2329 40635 2363
rect 40635 2329 40644 2363
rect 40592 2320 40644 2329
rect 43352 2388 43404 2440
rect 53840 2388 53892 2440
rect 54300 2524 54352 2576
rect 84936 2592 84988 2644
rect 104256 2592 104308 2644
rect 104348 2592 104400 2644
rect 107568 2592 107620 2644
rect 107660 2592 107712 2644
rect 108672 2592 108724 2644
rect 108764 2592 108816 2644
rect 114744 2592 114796 2644
rect 66168 2456 66220 2508
rect 54208 2431 54260 2440
rect 54208 2397 54217 2431
rect 54217 2397 54251 2431
rect 54251 2397 54260 2431
rect 54208 2388 54260 2397
rect 55496 2431 55548 2440
rect 55496 2397 55505 2431
rect 55505 2397 55539 2431
rect 55539 2397 55548 2431
rect 55496 2388 55548 2397
rect 57520 2388 57572 2440
rect 59176 2388 59228 2440
rect 61660 2388 61712 2440
rect 62212 2431 62264 2440
rect 62212 2397 62221 2431
rect 62221 2397 62255 2431
rect 62255 2397 62264 2431
rect 62212 2388 62264 2397
rect 62672 2388 62724 2440
rect 65432 2388 65484 2440
rect 66720 2388 66772 2440
rect 76472 2431 76524 2440
rect 76472 2397 76481 2431
rect 76481 2397 76515 2431
rect 76515 2397 76524 2431
rect 76472 2388 76524 2397
rect 78680 2431 78732 2440
rect 78680 2397 78689 2431
rect 78689 2397 78723 2431
rect 78723 2397 78732 2431
rect 78680 2388 78732 2397
rect 78956 2431 79008 2440
rect 78956 2397 78965 2431
rect 78965 2397 78999 2431
rect 78999 2397 79008 2431
rect 78956 2388 79008 2397
rect 22192 2252 22244 2304
rect 25872 2252 25924 2304
rect 29920 2295 29972 2304
rect 29920 2261 29929 2295
rect 29929 2261 29963 2295
rect 29963 2261 29972 2295
rect 29920 2252 29972 2261
rect 32680 2252 32732 2304
rect 38292 2252 38344 2304
rect 38384 2252 38436 2304
rect 39856 2252 39908 2304
rect 40224 2295 40276 2304
rect 40224 2261 40233 2295
rect 40233 2261 40267 2295
rect 40267 2261 40276 2295
rect 40224 2252 40276 2261
rect 41328 2295 41380 2304
rect 41328 2261 41337 2295
rect 41337 2261 41371 2295
rect 41371 2261 41380 2295
rect 41328 2252 41380 2261
rect 41512 2295 41564 2304
rect 41512 2261 41521 2295
rect 41521 2261 41555 2295
rect 41555 2261 41564 2295
rect 41512 2252 41564 2261
rect 42248 2295 42300 2304
rect 42248 2261 42257 2295
rect 42257 2261 42291 2295
rect 42291 2261 42300 2295
rect 42248 2252 42300 2261
rect 43352 2295 43404 2304
rect 43352 2261 43361 2295
rect 43361 2261 43395 2295
rect 43395 2261 43404 2295
rect 43352 2252 43404 2261
rect 53748 2252 53800 2304
rect 57980 2295 58032 2304
rect 57980 2261 57989 2295
rect 57989 2261 58023 2295
rect 58023 2261 58032 2295
rect 57980 2252 58032 2261
rect 59360 2252 59412 2304
rect 59820 2252 59872 2304
rect 61476 2252 61528 2304
rect 62396 2295 62448 2304
rect 62396 2261 62405 2295
rect 62405 2261 62439 2295
rect 62439 2261 62448 2295
rect 62396 2252 62448 2261
rect 63132 2295 63184 2304
rect 63132 2261 63141 2295
rect 63141 2261 63175 2295
rect 63175 2261 63184 2295
rect 63132 2252 63184 2261
rect 65984 2295 66036 2304
rect 65984 2261 65993 2295
rect 65993 2261 66027 2295
rect 66027 2261 66036 2295
rect 65984 2252 66036 2261
rect 81624 2431 81676 2440
rect 81624 2397 81633 2431
rect 81633 2397 81667 2431
rect 81667 2397 81676 2431
rect 81624 2388 81676 2397
rect 83832 2431 83884 2440
rect 83832 2397 83841 2431
rect 83841 2397 83875 2431
rect 83875 2397 83884 2431
rect 83832 2388 83884 2397
rect 84108 2499 84160 2508
rect 84108 2465 84117 2499
rect 84117 2465 84151 2499
rect 84151 2465 84160 2499
rect 84108 2456 84160 2465
rect 94688 2524 94740 2576
rect 94780 2524 94832 2576
rect 93860 2456 93912 2508
rect 94596 2456 94648 2508
rect 95240 2499 95292 2508
rect 95240 2465 95249 2499
rect 95249 2465 95283 2499
rect 95283 2465 95292 2499
rect 95240 2456 95292 2465
rect 97632 2524 97684 2576
rect 97724 2524 97776 2576
rect 96712 2456 96764 2508
rect 99656 2499 99708 2508
rect 99656 2465 99665 2499
rect 99665 2465 99699 2499
rect 99699 2465 99708 2499
rect 99656 2456 99708 2465
rect 100024 2456 100076 2508
rect 102140 2499 102192 2508
rect 102140 2465 102149 2499
rect 102149 2465 102183 2499
rect 102183 2465 102192 2499
rect 102140 2456 102192 2465
rect 104808 2499 104860 2508
rect 104808 2465 104817 2499
rect 104817 2465 104851 2499
rect 104851 2465 104860 2499
rect 104808 2456 104860 2465
rect 106188 2499 106240 2508
rect 106188 2465 106197 2499
rect 106197 2465 106231 2499
rect 106231 2465 106240 2499
rect 106188 2456 106240 2465
rect 107200 2499 107252 2508
rect 107200 2465 107209 2499
rect 107209 2465 107243 2499
rect 107243 2465 107252 2499
rect 107200 2456 107252 2465
rect 107660 2499 107712 2508
rect 107660 2465 107669 2499
rect 107669 2465 107703 2499
rect 107703 2465 107712 2499
rect 107660 2456 107712 2465
rect 84936 2388 84988 2440
rect 88524 2388 88576 2440
rect 88984 2388 89036 2440
rect 89076 2431 89128 2440
rect 89076 2397 89085 2431
rect 89085 2397 89119 2431
rect 89119 2397 89128 2431
rect 89076 2388 89128 2397
rect 90272 2388 90324 2440
rect 91100 2388 91152 2440
rect 92204 2431 92256 2440
rect 92204 2397 92213 2431
rect 92213 2397 92247 2431
rect 92247 2397 92256 2431
rect 92204 2388 92256 2397
rect 92848 2431 92900 2440
rect 92848 2397 92857 2431
rect 92857 2397 92891 2431
rect 92891 2397 92900 2431
rect 92848 2388 92900 2397
rect 94412 2388 94464 2440
rect 95516 2431 95568 2440
rect 95516 2397 95525 2431
rect 95525 2397 95559 2431
rect 95559 2397 95568 2431
rect 95516 2388 95568 2397
rect 98736 2388 98788 2440
rect 100944 2388 100996 2440
rect 101312 2431 101364 2440
rect 101312 2397 101321 2431
rect 101321 2397 101355 2431
rect 101355 2397 101364 2431
rect 101312 2388 101364 2397
rect 81164 2320 81216 2372
rect 92296 2320 92348 2372
rect 92572 2320 92624 2372
rect 88524 2295 88576 2304
rect 88524 2261 88533 2295
rect 88533 2261 88567 2295
rect 88567 2261 88576 2295
rect 88524 2252 88576 2261
rect 88800 2252 88852 2304
rect 90180 2295 90232 2304
rect 90180 2261 90189 2295
rect 90189 2261 90223 2295
rect 90223 2261 90232 2295
rect 90180 2252 90232 2261
rect 91192 2252 91244 2304
rect 93768 2295 93820 2304
rect 93768 2261 93777 2295
rect 93777 2261 93811 2295
rect 93811 2261 93820 2295
rect 93768 2252 93820 2261
rect 96068 2320 96120 2372
rect 97908 2320 97960 2372
rect 99012 2363 99064 2372
rect 99012 2329 99021 2363
rect 99021 2329 99055 2363
rect 99055 2329 99064 2363
rect 99012 2320 99064 2329
rect 100484 2320 100536 2372
rect 101496 2320 101548 2372
rect 106372 2320 106424 2372
rect 109040 2456 109092 2508
rect 109500 2499 109552 2508
rect 109500 2465 109509 2499
rect 109509 2465 109543 2499
rect 109543 2465 109552 2499
rect 109500 2456 109552 2465
rect 113364 2456 113416 2508
rect 108488 2388 108540 2440
rect 110696 2388 110748 2440
rect 112076 2388 112128 2440
rect 112168 2431 112220 2440
rect 112168 2397 112177 2431
rect 112177 2397 112211 2431
rect 112211 2397 112220 2431
rect 112168 2388 112220 2397
rect 114560 2524 114612 2576
rect 117320 2524 117372 2576
rect 113824 2456 113876 2508
rect 96252 2252 96304 2304
rect 96436 2252 96488 2304
rect 98828 2252 98880 2304
rect 99104 2252 99156 2304
rect 104900 2252 104952 2304
rect 107844 2252 107896 2304
rect 108580 2252 108632 2304
rect 110236 2252 110288 2304
rect 112352 2363 112404 2372
rect 112352 2329 112361 2363
rect 112361 2329 112395 2363
rect 112395 2329 112404 2363
rect 112352 2320 112404 2329
rect 117228 2388 117280 2440
rect 117320 2388 117372 2440
rect 124220 2635 124272 2644
rect 124220 2601 124229 2635
rect 124229 2601 124263 2635
rect 124263 2601 124272 2635
rect 124220 2592 124272 2601
rect 133880 2592 133932 2644
rect 139952 2592 140004 2644
rect 138940 2524 138992 2576
rect 140964 2592 141016 2644
rect 141148 2635 141200 2644
rect 141148 2601 141157 2635
rect 141157 2601 141191 2635
rect 141191 2601 141200 2635
rect 141148 2592 141200 2601
rect 142252 2592 142304 2644
rect 142436 2592 142488 2644
rect 146668 2592 146720 2644
rect 141792 2524 141844 2576
rect 153016 2592 153068 2644
rect 153752 2592 153804 2644
rect 155224 2592 155276 2644
rect 156420 2592 156472 2644
rect 149060 2524 149112 2576
rect 152740 2524 152792 2576
rect 152924 2524 152976 2576
rect 118700 2456 118752 2508
rect 120264 2499 120316 2508
rect 120264 2465 120273 2499
rect 120273 2465 120307 2499
rect 120307 2465 120316 2499
rect 120264 2456 120316 2465
rect 118976 2388 119028 2440
rect 121920 2456 121972 2508
rect 124772 2499 124824 2508
rect 124772 2465 124781 2499
rect 124781 2465 124815 2499
rect 124815 2465 124824 2499
rect 124772 2456 124824 2465
rect 130200 2456 130252 2508
rect 135352 2456 135404 2508
rect 139308 2499 139360 2508
rect 139308 2465 139317 2499
rect 139317 2465 139351 2499
rect 139351 2465 139360 2499
rect 139308 2456 139360 2465
rect 139952 2499 140004 2508
rect 139952 2465 139961 2499
rect 139961 2465 139995 2499
rect 139995 2465 140004 2499
rect 139952 2456 140004 2465
rect 121184 2388 121236 2440
rect 124312 2388 124364 2440
rect 124956 2431 125008 2440
rect 124956 2397 124965 2431
rect 124965 2397 124999 2431
rect 124999 2397 125008 2431
rect 124956 2388 125008 2397
rect 126060 2431 126112 2440
rect 126060 2397 126069 2431
rect 126069 2397 126103 2431
rect 126103 2397 126112 2431
rect 126060 2388 126112 2397
rect 126704 2388 126756 2440
rect 128360 2388 128412 2440
rect 129004 2431 129056 2440
rect 129004 2397 129013 2431
rect 129013 2397 129047 2431
rect 129047 2397 129056 2431
rect 129004 2388 129056 2397
rect 129648 2388 129700 2440
rect 131764 2388 131816 2440
rect 133512 2388 133564 2440
rect 133696 2388 133748 2440
rect 134340 2388 134392 2440
rect 128820 2320 128872 2372
rect 115020 2252 115072 2304
rect 116032 2252 116084 2304
rect 117596 2252 117648 2304
rect 118056 2252 118108 2304
rect 122656 2295 122708 2304
rect 122656 2261 122665 2295
rect 122665 2261 122699 2295
rect 122699 2261 122708 2295
rect 122656 2252 122708 2261
rect 125140 2295 125192 2304
rect 125140 2261 125149 2295
rect 125149 2261 125183 2295
rect 125183 2261 125192 2295
rect 125140 2252 125192 2261
rect 126244 2295 126296 2304
rect 126244 2261 126253 2295
rect 126253 2261 126287 2295
rect 126287 2261 126296 2295
rect 126244 2252 126296 2261
rect 126980 2295 127032 2304
rect 126980 2261 126989 2295
rect 126989 2261 127023 2295
rect 127023 2261 127032 2295
rect 126980 2252 127032 2261
rect 128452 2295 128504 2304
rect 128452 2261 128461 2295
rect 128461 2261 128495 2295
rect 128495 2261 128504 2295
rect 128452 2252 128504 2261
rect 129188 2295 129240 2304
rect 129188 2261 129197 2295
rect 129197 2261 129231 2295
rect 129231 2261 129240 2295
rect 129188 2252 129240 2261
rect 130752 2295 130804 2304
rect 130752 2261 130761 2295
rect 130761 2261 130795 2295
rect 130795 2261 130804 2295
rect 130752 2252 130804 2261
rect 131672 2295 131724 2304
rect 131672 2261 131681 2295
rect 131681 2261 131715 2295
rect 131715 2261 131724 2295
rect 131672 2252 131724 2261
rect 133236 2295 133288 2304
rect 133236 2261 133245 2295
rect 133245 2261 133279 2295
rect 133279 2261 133288 2295
rect 133236 2252 133288 2261
rect 135352 2252 135404 2304
rect 139492 2431 139544 2440
rect 139492 2397 139501 2431
rect 139501 2397 139535 2431
rect 139535 2397 139544 2431
rect 139492 2388 139544 2397
rect 140228 2431 140280 2440
rect 140228 2397 140237 2431
rect 140237 2397 140271 2431
rect 140271 2397 140280 2431
rect 140228 2388 140280 2397
rect 140320 2431 140372 2440
rect 140688 2456 140740 2508
rect 143356 2456 143408 2508
rect 146300 2499 146352 2508
rect 146300 2465 146309 2499
rect 146309 2465 146343 2499
rect 146343 2465 146352 2499
rect 146300 2456 146352 2465
rect 148600 2499 148652 2508
rect 148600 2465 148609 2499
rect 148609 2465 148643 2499
rect 148643 2465 148652 2499
rect 148600 2456 148652 2465
rect 148784 2499 148836 2508
rect 148784 2465 148793 2499
rect 148793 2465 148827 2499
rect 148827 2465 148836 2499
rect 148784 2456 148836 2465
rect 150256 2499 150308 2508
rect 150256 2465 150265 2499
rect 150265 2465 150299 2499
rect 150299 2465 150308 2499
rect 150256 2456 150308 2465
rect 150808 2456 150860 2508
rect 151360 2499 151412 2508
rect 151360 2465 151369 2499
rect 151369 2465 151403 2499
rect 151403 2465 151412 2499
rect 151360 2456 151412 2465
rect 151820 2456 151872 2508
rect 154488 2524 154540 2576
rect 158444 2524 158496 2576
rect 166540 2524 166592 2576
rect 168380 2524 168432 2576
rect 140320 2397 140354 2431
rect 140354 2397 140372 2431
rect 140320 2388 140372 2397
rect 141608 2431 141660 2440
rect 141608 2397 141617 2431
rect 141617 2397 141651 2431
rect 141651 2397 141660 2431
rect 141608 2388 141660 2397
rect 141976 2431 142028 2440
rect 141976 2397 141985 2431
rect 141985 2397 142019 2431
rect 142019 2397 142028 2431
rect 141976 2388 142028 2397
rect 142160 2388 142212 2440
rect 145380 2431 145432 2440
rect 145380 2397 145389 2431
rect 145389 2397 145423 2431
rect 145423 2397 145432 2431
rect 145380 2388 145432 2397
rect 141240 2320 141292 2372
rect 144736 2320 144788 2372
rect 146392 2320 146444 2372
rect 150900 2431 150952 2440
rect 150900 2397 150909 2431
rect 150909 2397 150943 2431
rect 150943 2397 150952 2431
rect 150900 2388 150952 2397
rect 148508 2320 148560 2372
rect 150440 2320 150492 2372
rect 153384 2388 153436 2440
rect 154120 2388 154172 2440
rect 154488 2388 154540 2440
rect 155592 2431 155644 2440
rect 155592 2397 155601 2431
rect 155601 2397 155635 2431
rect 155635 2397 155644 2431
rect 155592 2388 155644 2397
rect 156604 2431 156656 2440
rect 156604 2397 156613 2431
rect 156613 2397 156647 2431
rect 156647 2397 156656 2431
rect 156604 2388 156656 2397
rect 156972 2388 157024 2440
rect 156420 2320 156472 2372
rect 156696 2320 156748 2372
rect 157708 2431 157760 2440
rect 157708 2397 157717 2431
rect 157717 2397 157751 2431
rect 157751 2397 157760 2431
rect 157708 2388 157760 2397
rect 158444 2388 158496 2440
rect 159916 2431 159968 2440
rect 159916 2397 159925 2431
rect 159925 2397 159959 2431
rect 159959 2397 159968 2431
rect 159916 2388 159968 2397
rect 160008 2431 160060 2440
rect 160008 2397 160017 2431
rect 160017 2397 160051 2431
rect 160051 2397 160060 2431
rect 160008 2388 160060 2397
rect 161480 2431 161532 2440
rect 161480 2397 161489 2431
rect 161489 2397 161523 2431
rect 161523 2397 161532 2431
rect 161480 2388 161532 2397
rect 163964 2388 164016 2440
rect 165620 2388 165672 2440
rect 165804 2431 165856 2440
rect 165804 2397 165813 2431
rect 165813 2397 165847 2431
rect 165847 2397 165856 2431
rect 165804 2388 165856 2397
rect 167460 2388 167512 2440
rect 167920 2431 167972 2440
rect 167920 2397 167929 2431
rect 167929 2397 167963 2431
rect 167963 2397 167972 2431
rect 167920 2388 167972 2397
rect 168012 2431 168064 2440
rect 168012 2397 168021 2431
rect 168021 2397 168055 2431
rect 168055 2397 168064 2431
rect 168012 2388 168064 2397
rect 168288 2388 168340 2440
rect 158996 2363 159048 2372
rect 158996 2329 159005 2363
rect 159005 2329 159039 2363
rect 159039 2329 159048 2363
rect 158996 2320 159048 2329
rect 167736 2320 167788 2372
rect 140780 2252 140832 2304
rect 140964 2252 141016 2304
rect 144276 2252 144328 2304
rect 146852 2252 146904 2304
rect 148324 2252 148376 2304
rect 151084 2252 151136 2304
rect 151452 2252 151504 2304
rect 153476 2252 153528 2304
rect 157248 2252 157300 2304
rect 160836 2295 160888 2304
rect 160836 2261 160845 2295
rect 160845 2261 160879 2295
rect 160879 2261 160888 2295
rect 160836 2252 160888 2261
rect 161664 2295 161716 2304
rect 161664 2261 161673 2295
rect 161673 2261 161707 2295
rect 161707 2261 161716 2295
rect 161664 2252 161716 2261
rect 162400 2295 162452 2304
rect 162400 2261 162409 2295
rect 162409 2261 162443 2295
rect 162443 2261 162452 2295
rect 162400 2252 162452 2261
rect 163872 2295 163924 2304
rect 163872 2261 163881 2295
rect 163881 2261 163915 2295
rect 163915 2261 163924 2295
rect 163872 2252 163924 2261
rect 165252 2295 165304 2304
rect 165252 2261 165261 2295
rect 165261 2261 165295 2295
rect 165295 2261 165304 2295
rect 165252 2252 165304 2261
rect 165988 2295 166040 2304
rect 165988 2261 165997 2295
rect 165997 2261 166031 2295
rect 166031 2261 166040 2295
rect 165988 2252 166040 2261
rect 166816 2295 166868 2304
rect 166816 2261 166825 2295
rect 166825 2261 166859 2295
rect 166859 2261 166868 2295
rect 166816 2252 166868 2261
rect 168196 2295 168248 2304
rect 168196 2261 168205 2295
rect 168205 2261 168239 2295
rect 168239 2261 168248 2295
rect 168196 2252 168248 2261
rect 168288 2252 168340 2304
rect 176660 2431 176712 2440
rect 176660 2397 176669 2431
rect 176669 2397 176703 2431
rect 176703 2397 176712 2431
rect 176660 2388 176712 2397
rect 176936 2431 176988 2440
rect 176936 2397 176945 2431
rect 176945 2397 176979 2431
rect 176979 2397 176988 2431
rect 176936 2388 176988 2397
rect 179604 2431 179656 2440
rect 179604 2397 179613 2431
rect 179613 2397 179647 2431
rect 179647 2397 179656 2431
rect 179604 2388 179656 2397
rect 172428 2320 172480 2372
rect 181812 2431 181864 2440
rect 181812 2397 181821 2431
rect 181821 2397 181855 2431
rect 181855 2397 181864 2431
rect 181812 2388 181864 2397
rect 184756 2431 184808 2440
rect 184756 2397 184765 2431
rect 184765 2397 184799 2431
rect 184799 2397 184808 2431
rect 184756 2388 184808 2397
rect 190460 2592 190512 2644
rect 191840 2592 191892 2644
rect 198740 2635 198792 2644
rect 198740 2601 198749 2635
rect 198749 2601 198783 2635
rect 198783 2601 198792 2635
rect 198740 2592 198792 2601
rect 192392 2524 192444 2576
rect 192852 2524 192904 2576
rect 217600 2592 217652 2644
rect 200212 2524 200264 2576
rect 201500 2524 201552 2576
rect 202788 2456 202840 2508
rect 186964 2431 187016 2440
rect 186964 2397 186973 2431
rect 186973 2397 187007 2431
rect 187007 2397 187016 2431
rect 186964 2388 187016 2397
rect 190920 2388 190972 2440
rect 191012 2388 191064 2440
rect 192208 2388 192260 2440
rect 195704 2388 195756 2440
rect 196164 2431 196216 2440
rect 196164 2397 196173 2431
rect 196173 2397 196207 2431
rect 196207 2397 196216 2431
rect 196164 2388 196216 2397
rect 197544 2388 197596 2440
rect 198280 2388 198332 2440
rect 199752 2388 199804 2440
rect 200212 2431 200264 2440
rect 200212 2397 200221 2431
rect 200221 2397 200255 2431
rect 200255 2397 200264 2431
rect 200212 2388 200264 2397
rect 201040 2431 201092 2440
rect 201040 2397 201049 2431
rect 201049 2397 201083 2431
rect 201083 2397 201092 2431
rect 201040 2388 201092 2397
rect 202696 2388 202748 2440
rect 203156 2431 203208 2440
rect 203156 2397 203165 2431
rect 203165 2397 203199 2431
rect 203199 2397 203208 2431
rect 203156 2388 203208 2397
rect 191196 2363 191248 2372
rect 191196 2329 191205 2363
rect 191205 2329 191239 2363
rect 191239 2329 191248 2363
rect 191196 2320 191248 2329
rect 191380 2320 191432 2372
rect 218152 2567 218204 2576
rect 218152 2533 218161 2567
rect 218161 2533 218195 2567
rect 218195 2533 218204 2567
rect 218152 2524 218204 2533
rect 219256 2592 219308 2644
rect 224500 2592 224552 2644
rect 222016 2524 222068 2576
rect 225788 2524 225840 2576
rect 226984 2635 227036 2644
rect 226984 2601 226993 2635
rect 226993 2601 227027 2635
rect 227027 2601 227036 2635
rect 226984 2592 227036 2601
rect 227076 2592 227128 2644
rect 228272 2592 228324 2644
rect 243912 2592 243964 2644
rect 245476 2592 245528 2644
rect 248880 2592 248932 2644
rect 228456 2524 228508 2576
rect 230572 2524 230624 2576
rect 230756 2524 230808 2576
rect 233056 2524 233108 2576
rect 246856 2524 246908 2576
rect 248512 2524 248564 2576
rect 209688 2456 209740 2508
rect 208676 2388 208728 2440
rect 208952 2431 209004 2440
rect 208952 2397 208961 2431
rect 208961 2397 208995 2431
rect 208995 2397 209004 2431
rect 208952 2388 209004 2397
rect 209044 2388 209096 2440
rect 211896 2363 211948 2372
rect 211896 2329 211905 2363
rect 211905 2329 211939 2363
rect 211939 2329 211948 2363
rect 211896 2320 211948 2329
rect 191012 2252 191064 2304
rect 194600 2252 194652 2304
rect 196072 2252 196124 2304
rect 196624 2252 196676 2304
rect 197360 2252 197412 2304
rect 201224 2295 201276 2304
rect 201224 2261 201233 2295
rect 201233 2261 201267 2295
rect 201267 2261 201276 2295
rect 201224 2252 201276 2261
rect 204076 2295 204128 2304
rect 204076 2261 204085 2295
rect 204085 2261 204119 2295
rect 204119 2261 204128 2295
rect 204076 2252 204128 2261
rect 208124 2295 208176 2304
rect 208124 2261 208133 2295
rect 208133 2261 208167 2295
rect 208167 2261 208176 2295
rect 208124 2252 208176 2261
rect 212540 2499 212592 2508
rect 212540 2465 212549 2499
rect 212549 2465 212583 2499
rect 212583 2465 212592 2499
rect 212540 2456 212592 2465
rect 213828 2456 213880 2508
rect 216772 2499 216824 2508
rect 216772 2465 216781 2499
rect 216781 2465 216815 2499
rect 216815 2465 216824 2499
rect 216772 2456 216824 2465
rect 217508 2499 217560 2508
rect 217508 2465 217517 2499
rect 217517 2465 217551 2499
rect 217551 2465 217560 2499
rect 217508 2456 217560 2465
rect 217600 2456 217652 2508
rect 221832 2456 221884 2508
rect 223120 2499 223172 2508
rect 223120 2465 223129 2499
rect 223129 2465 223163 2499
rect 223163 2465 223172 2499
rect 223120 2456 223172 2465
rect 212356 2431 212408 2440
rect 212356 2397 212365 2431
rect 212365 2397 212399 2431
rect 212399 2397 212408 2431
rect 212356 2388 212408 2397
rect 214380 2388 214432 2440
rect 214472 2252 214524 2304
rect 217692 2431 217744 2440
rect 217692 2397 217701 2431
rect 217701 2397 217735 2431
rect 217735 2397 217744 2431
rect 217692 2388 217744 2397
rect 218428 2431 218480 2440
rect 218428 2397 218437 2431
rect 218437 2397 218471 2431
rect 218471 2397 218480 2431
rect 218428 2388 218480 2397
rect 218612 2388 218664 2440
rect 218704 2431 218756 2440
rect 218704 2397 218713 2431
rect 218713 2397 218747 2431
rect 218747 2397 218756 2431
rect 218704 2388 218756 2397
rect 220544 2431 220596 2440
rect 220544 2397 220553 2431
rect 220553 2397 220587 2431
rect 220587 2397 220596 2431
rect 220544 2388 220596 2397
rect 220636 2431 220688 2440
rect 220636 2397 220645 2431
rect 220645 2397 220679 2431
rect 220679 2397 220688 2431
rect 220636 2388 220688 2397
rect 220820 2388 220872 2440
rect 221372 2431 221424 2440
rect 221372 2397 221381 2431
rect 221381 2397 221415 2431
rect 221415 2397 221424 2431
rect 221372 2388 221424 2397
rect 222568 2320 222620 2372
rect 224132 2388 224184 2440
rect 225788 2388 225840 2440
rect 226800 2388 226852 2440
rect 228456 2388 228508 2440
rect 219624 2252 219676 2304
rect 219716 2252 219768 2304
rect 225420 2320 225472 2372
rect 240048 2456 240100 2508
rect 242900 2456 242952 2508
rect 248604 2456 248656 2508
rect 230940 2388 230992 2440
rect 231768 2388 231820 2440
rect 232596 2388 232648 2440
rect 232964 2431 233016 2440
rect 232964 2397 232973 2431
rect 232973 2397 233007 2431
rect 233007 2397 233016 2431
rect 232964 2388 233016 2397
rect 234988 2431 235040 2440
rect 234988 2397 234997 2431
rect 234997 2397 235031 2431
rect 235031 2397 235040 2431
rect 234988 2388 235040 2397
rect 235816 2431 235868 2440
rect 235816 2397 235825 2431
rect 235825 2397 235859 2431
rect 235859 2397 235868 2431
rect 235816 2388 235868 2397
rect 229928 2320 229980 2372
rect 236920 2388 236972 2440
rect 243452 2431 243504 2440
rect 243452 2397 243461 2431
rect 243461 2397 243495 2431
rect 243495 2397 243504 2431
rect 243452 2388 243504 2397
rect 243728 2431 243780 2440
rect 243728 2397 243737 2431
rect 243737 2397 243771 2431
rect 243771 2397 243780 2431
rect 243728 2388 243780 2397
rect 244188 2388 244240 2440
rect 245016 2431 245068 2440
rect 245016 2397 245025 2431
rect 245025 2397 245059 2431
rect 245059 2397 245068 2431
rect 245016 2388 245068 2397
rect 248788 2431 248840 2440
rect 248788 2397 248797 2431
rect 248797 2397 248831 2431
rect 248831 2397 248840 2431
rect 248788 2388 248840 2397
rect 256516 2524 256568 2576
rect 259736 2524 259788 2576
rect 251456 2499 251508 2508
rect 251456 2465 251465 2499
rect 251465 2465 251499 2499
rect 251499 2465 251508 2499
rect 251456 2456 251508 2465
rect 253480 2456 253532 2508
rect 252652 2388 252704 2440
rect 254860 2431 254912 2440
rect 254860 2397 254869 2431
rect 254869 2397 254903 2431
rect 254903 2397 254912 2431
rect 254860 2388 254912 2397
rect 246304 2363 246356 2372
rect 246304 2329 246313 2363
rect 246313 2329 246347 2363
rect 246347 2329 246356 2363
rect 246304 2320 246356 2329
rect 252376 2320 252428 2372
rect 253112 2363 253164 2372
rect 253112 2329 253121 2363
rect 253121 2329 253155 2363
rect 253155 2329 253164 2363
rect 253112 2320 253164 2329
rect 224224 2295 224276 2304
rect 224224 2261 224233 2295
rect 224233 2261 224267 2295
rect 224267 2261 224276 2295
rect 224224 2252 224276 2261
rect 224776 2295 224828 2304
rect 224776 2261 224785 2295
rect 224785 2261 224819 2295
rect 224819 2261 224828 2295
rect 224776 2252 224828 2261
rect 225696 2295 225748 2304
rect 225696 2261 225705 2295
rect 225705 2261 225739 2295
rect 225739 2261 225748 2295
rect 225696 2252 225748 2261
rect 226340 2252 226392 2304
rect 227996 2295 228048 2304
rect 227996 2261 228005 2295
rect 228005 2261 228039 2295
rect 228039 2261 228048 2295
rect 227996 2252 228048 2261
rect 230020 2295 230072 2304
rect 230020 2261 230029 2295
rect 230029 2261 230063 2295
rect 230063 2261 230072 2295
rect 230020 2252 230072 2261
rect 231584 2295 231636 2304
rect 231584 2261 231593 2295
rect 231593 2261 231627 2295
rect 231627 2261 231636 2295
rect 231584 2252 231636 2261
rect 232412 2295 232464 2304
rect 232412 2261 232421 2295
rect 232421 2261 232455 2295
rect 232455 2261 232464 2295
rect 232412 2252 232464 2261
rect 233148 2295 233200 2304
rect 233148 2261 233157 2295
rect 233157 2261 233191 2295
rect 233191 2261 233200 2295
rect 233148 2252 233200 2261
rect 235172 2295 235224 2304
rect 235172 2261 235181 2295
rect 235181 2261 235215 2295
rect 235215 2261 235224 2295
rect 235172 2252 235224 2261
rect 236184 2295 236236 2304
rect 236184 2261 236193 2295
rect 236193 2261 236227 2295
rect 236227 2261 236236 2295
rect 236184 2252 236236 2261
rect 236828 2295 236880 2304
rect 236828 2261 236837 2295
rect 236837 2261 236871 2295
rect 236871 2261 236880 2295
rect 236828 2252 236880 2261
rect 243636 2252 243688 2304
rect 256424 2431 256476 2440
rect 256424 2397 256433 2431
rect 256433 2397 256467 2431
rect 256467 2397 256476 2431
rect 256424 2388 256476 2397
rect 257528 2320 257580 2372
rect 258356 2320 258408 2372
rect 260104 2363 260156 2372
rect 260104 2329 260113 2363
rect 260113 2329 260147 2363
rect 260147 2329 260156 2363
rect 260104 2320 260156 2329
rect 261576 2499 261628 2508
rect 261576 2465 261585 2499
rect 261585 2465 261619 2499
rect 261619 2465 261628 2499
rect 261576 2456 261628 2465
rect 262220 2524 262272 2576
rect 267004 2592 267056 2644
rect 269856 2592 269908 2644
rect 267924 2524 267976 2576
rect 261024 2388 261076 2440
rect 261484 2388 261536 2440
rect 263140 2431 263192 2440
rect 263140 2397 263149 2431
rect 263149 2397 263183 2431
rect 263183 2397 263192 2431
rect 263140 2388 263192 2397
rect 263968 2499 264020 2508
rect 263968 2465 263977 2499
rect 263977 2465 264011 2499
rect 264011 2465 264020 2499
rect 263968 2456 264020 2465
rect 267556 2456 267608 2508
rect 264336 2388 264388 2440
rect 265164 2431 265216 2440
rect 265164 2397 265173 2431
rect 265173 2397 265207 2431
rect 265207 2397 265216 2431
rect 265164 2388 265216 2397
rect 267004 2388 267056 2440
rect 268292 2388 268344 2440
rect 268476 2431 268528 2440
rect 268476 2397 268485 2431
rect 268485 2397 268519 2431
rect 268519 2397 268528 2431
rect 268476 2388 268528 2397
rect 268660 2456 268712 2508
rect 269120 2431 269172 2440
rect 269120 2397 269129 2431
rect 269129 2397 269163 2431
rect 269163 2397 269172 2431
rect 269120 2388 269172 2397
rect 270040 2388 270092 2440
rect 263968 2320 264020 2372
rect 264244 2320 264296 2372
rect 268384 2320 268436 2372
rect 259920 2252 259972 2304
rect 260196 2295 260248 2304
rect 260196 2261 260205 2295
rect 260205 2261 260239 2295
rect 260239 2261 260248 2295
rect 260196 2252 260248 2261
rect 263324 2295 263376 2304
rect 263324 2261 263333 2295
rect 263333 2261 263367 2295
rect 263367 2261 263376 2295
rect 263324 2252 263376 2261
rect 264888 2252 264940 2304
rect 266912 2295 266964 2304
rect 266912 2261 266921 2295
rect 266921 2261 266955 2295
rect 266955 2261 266964 2295
rect 266912 2252 266964 2261
rect 269212 2252 269264 2304
rect 270132 2252 270184 2304
rect 270776 2295 270828 2304
rect 270776 2261 270785 2295
rect 270785 2261 270819 2295
rect 270819 2261 270828 2295
rect 270776 2252 270828 2261
rect 68546 2150 68598 2202
rect 68610 2150 68662 2202
rect 68674 2150 68726 2202
rect 68738 2150 68790 2202
rect 68802 2150 68854 2202
rect 136143 2150 136195 2202
rect 136207 2150 136259 2202
rect 136271 2150 136323 2202
rect 136335 2150 136387 2202
rect 136399 2150 136451 2202
rect 203740 2150 203792 2202
rect 203804 2150 203856 2202
rect 203868 2150 203920 2202
rect 203932 2150 203984 2202
rect 203996 2150 204048 2202
rect 271337 2150 271389 2202
rect 271401 2150 271453 2202
rect 271465 2150 271517 2202
rect 271529 2150 271581 2202
rect 271593 2150 271645 2202
rect 1860 2048 1912 2100
rect 12072 2091 12124 2100
rect 12072 2057 12081 2091
rect 12081 2057 12115 2091
rect 12115 2057 12124 2091
rect 12072 2048 12124 2057
rect 12808 2091 12860 2100
rect 12808 2057 12817 2091
rect 12817 2057 12851 2091
rect 12851 2057 12860 2091
rect 12808 2048 12860 2057
rect 1676 1955 1728 1964
rect 1676 1921 1685 1955
rect 1685 1921 1719 1955
rect 1719 1921 1728 1955
rect 1676 1912 1728 1921
rect 5540 1912 5592 1964
rect 3792 1887 3844 1896
rect 3792 1853 3801 1887
rect 3801 1853 3835 1887
rect 3835 1853 3844 1887
rect 3792 1844 3844 1853
rect 5172 1887 5224 1896
rect 5172 1853 5181 1887
rect 5181 1853 5215 1887
rect 5215 1853 5224 1887
rect 5172 1844 5224 1853
rect 7380 1955 7432 1964
rect 7380 1921 7389 1955
rect 7389 1921 7423 1955
rect 7423 1921 7432 1955
rect 7380 1912 7432 1921
rect 8668 1955 8720 1964
rect 8668 1921 8677 1955
rect 8677 1921 8711 1955
rect 8711 1921 8720 1955
rect 8668 1912 8720 1921
rect 11980 1955 12032 1964
rect 11980 1921 11989 1955
rect 11989 1921 12023 1955
rect 12023 1921 12032 1955
rect 11980 1912 12032 1921
rect 12716 1955 12768 1964
rect 12716 1921 12725 1955
rect 12725 1921 12759 1955
rect 12759 1921 12768 1955
rect 12716 1912 12768 1921
rect 14372 1955 14424 1964
rect 14372 1921 14381 1955
rect 14381 1921 14415 1955
rect 14415 1921 14424 1955
rect 14372 1912 14424 1921
rect 7104 1887 7156 1896
rect 7104 1853 7113 1887
rect 7113 1853 7147 1887
rect 7147 1853 7156 1887
rect 7104 1844 7156 1853
rect 8392 1887 8444 1896
rect 8392 1853 8401 1887
rect 8401 1853 8435 1887
rect 8435 1853 8444 1887
rect 8392 1844 8444 1853
rect 9680 1887 9732 1896
rect 9680 1853 9689 1887
rect 9689 1853 9723 1887
rect 9723 1853 9732 1887
rect 9680 1844 9732 1853
rect 14096 1887 14148 1896
rect 14096 1853 14105 1887
rect 14105 1853 14139 1887
rect 14139 1853 14148 1887
rect 14096 1844 14148 1853
rect 15476 1887 15528 1896
rect 15476 1853 15485 1887
rect 15485 1853 15519 1887
rect 15519 1853 15528 1887
rect 15476 1844 15528 1853
rect 15844 1980 15896 2032
rect 17868 1955 17920 1964
rect 17868 1921 17877 1955
rect 17877 1921 17911 1955
rect 17911 1921 17920 1955
rect 17868 1912 17920 1921
rect 18052 1955 18104 1964
rect 18052 1921 18061 1955
rect 18061 1921 18095 1955
rect 18095 1921 18104 1955
rect 18052 1912 18104 1921
rect 22192 1912 22244 1964
rect 22284 1955 22336 1964
rect 22284 1921 22293 1955
rect 22293 1921 22327 1955
rect 22327 1921 22336 1955
rect 22284 1912 22336 1921
rect 22376 1912 22428 1964
rect 15844 1776 15896 1828
rect 22468 1844 22520 1896
rect 23112 1887 23164 1896
rect 23112 1853 23121 1887
rect 23121 1853 23155 1887
rect 23155 1853 23164 1887
rect 23112 1844 23164 1853
rect 23296 1955 23348 1964
rect 23296 1921 23305 1955
rect 23305 1921 23339 1955
rect 23339 1921 23348 1955
rect 23296 1912 23348 1921
rect 24124 1912 24176 1964
rect 24952 1955 25004 1964
rect 24952 1921 24961 1955
rect 24961 1921 24995 1955
rect 24995 1921 25004 1955
rect 24952 1912 25004 1921
rect 25872 2023 25924 2032
rect 25872 1989 25881 2023
rect 25881 1989 25915 2023
rect 25915 1989 25924 2023
rect 25872 1980 25924 1989
rect 37648 2048 37700 2100
rect 38476 2048 38528 2100
rect 26332 1912 26384 1964
rect 27344 1912 27396 1964
rect 32496 1955 32548 1964
rect 32496 1921 32505 1955
rect 32505 1921 32539 1955
rect 32539 1921 32548 1955
rect 32496 1912 32548 1921
rect 32680 1912 32732 1964
rect 27620 1844 27672 1896
rect 27712 1887 27764 1896
rect 27712 1853 27721 1887
rect 27721 1853 27755 1887
rect 27755 1853 27764 1887
rect 27712 1844 27764 1853
rect 28540 1887 28592 1896
rect 28540 1853 28549 1887
rect 28549 1853 28583 1887
rect 28583 1853 28592 1887
rect 28540 1844 28592 1853
rect 29460 1844 29512 1896
rect 29736 1887 29788 1896
rect 29736 1853 29745 1887
rect 29745 1853 29779 1887
rect 29779 1853 29788 1887
rect 29736 1844 29788 1853
rect 30104 1844 30156 1896
rect 30748 1887 30800 1896
rect 30748 1853 30757 1887
rect 30757 1853 30791 1887
rect 30791 1853 30800 1887
rect 30748 1844 30800 1853
rect 31300 1844 31352 1896
rect 31852 1844 31904 1896
rect 38568 1980 38620 2032
rect 38108 1955 38160 1964
rect 38108 1921 38117 1955
rect 38117 1921 38151 1955
rect 38151 1921 38160 1955
rect 38108 1912 38160 1921
rect 39028 1980 39080 2032
rect 39304 1980 39356 2032
rect 39396 2023 39448 2032
rect 39396 1989 39405 2023
rect 39405 1989 39439 2023
rect 39439 1989 39448 2023
rect 39396 1980 39448 1989
rect 40592 2048 40644 2100
rect 41512 2048 41564 2100
rect 73436 2048 73488 2100
rect 73620 2048 73672 2100
rect 80060 2048 80112 2100
rect 89352 2048 89404 2100
rect 90272 2091 90324 2100
rect 90272 2057 90281 2091
rect 90281 2057 90315 2091
rect 90315 2057 90324 2091
rect 90272 2048 90324 2057
rect 91100 2091 91152 2100
rect 91100 2057 91109 2091
rect 91109 2057 91143 2091
rect 91143 2057 91152 2091
rect 91100 2048 91152 2057
rect 91836 2048 91888 2100
rect 93216 2048 93268 2100
rect 94136 2048 94188 2100
rect 94688 2048 94740 2100
rect 96068 2048 96120 2100
rect 96436 2091 96488 2100
rect 96436 2057 96445 2091
rect 96445 2057 96479 2091
rect 96479 2057 96488 2091
rect 96436 2048 96488 2057
rect 39580 1980 39632 2032
rect 40040 1980 40092 2032
rect 53288 2023 53340 2032
rect 53288 1989 53297 2023
rect 53297 1989 53331 2023
rect 53331 1989 53340 2023
rect 53288 1980 53340 1989
rect 55496 1980 55548 2032
rect 45468 1955 45520 1964
rect 45468 1921 45477 1955
rect 45477 1921 45511 1955
rect 45511 1921 45520 1955
rect 45468 1912 45520 1921
rect 53748 1912 53800 1964
rect 54208 1912 54260 1964
rect 54576 1912 54628 1964
rect 56232 1980 56284 2032
rect 57520 2023 57572 2032
rect 57520 1989 57529 2023
rect 57529 1989 57563 2023
rect 57563 1989 57572 2023
rect 57520 1980 57572 1989
rect 59176 2023 59228 2032
rect 59176 1989 59185 2023
rect 59185 1989 59219 2023
rect 59219 1989 59228 2023
rect 59176 1980 59228 1989
rect 61660 2023 61712 2032
rect 61660 1989 61669 2023
rect 61669 1989 61703 2023
rect 61703 1989 61712 2023
rect 61660 1980 61712 1989
rect 62672 2023 62724 2032
rect 62672 1989 62681 2023
rect 62681 1989 62715 2023
rect 62715 1989 62724 2023
rect 62672 1980 62724 1989
rect 40132 1844 40184 1896
rect 41052 1844 41104 1896
rect 53288 1844 53340 1896
rect 54116 1844 54168 1896
rect 38384 1776 38436 1828
rect 45284 1819 45336 1828
rect 45284 1785 45293 1819
rect 45293 1785 45327 1819
rect 45327 1785 45336 1819
rect 45284 1776 45336 1785
rect 56416 1955 56468 1964
rect 56416 1921 56425 1955
rect 56425 1921 56459 1955
rect 56459 1921 56468 1955
rect 56416 1912 56468 1921
rect 56876 1912 56928 1964
rect 58072 1955 58124 1964
rect 58072 1921 58081 1955
rect 58081 1921 58115 1955
rect 58115 1921 58124 1955
rect 58072 1912 58124 1921
rect 58624 1912 58676 1964
rect 58532 1844 58584 1896
rect 59728 1955 59780 1964
rect 59728 1921 59737 1955
rect 59737 1921 59771 1955
rect 59771 1921 59780 1955
rect 59728 1912 59780 1921
rect 59820 1955 59872 1964
rect 59820 1921 59829 1955
rect 59829 1921 59863 1955
rect 59863 1921 59872 1955
rect 59820 1912 59872 1921
rect 60556 1955 60608 1964
rect 60556 1921 60565 1955
rect 60565 1921 60599 1955
rect 60599 1921 60608 1955
rect 60556 1912 60608 1921
rect 61292 1955 61344 1964
rect 61292 1921 61301 1955
rect 61301 1921 61335 1955
rect 61335 1921 61344 1955
rect 61292 1912 61344 1921
rect 62304 1955 62356 1964
rect 62304 1921 62313 1955
rect 62313 1921 62347 1955
rect 62347 1921 62356 1955
rect 62304 1912 62356 1921
rect 62488 1955 62540 1964
rect 62488 1921 62497 1955
rect 62497 1921 62531 1955
rect 62531 1921 62540 1955
rect 62488 1912 62540 1921
rect 63224 1912 63276 1964
rect 64052 1955 64104 1964
rect 64052 1921 64061 1955
rect 64061 1921 64095 1955
rect 64095 1921 64104 1955
rect 64052 1912 64104 1921
rect 65432 2023 65484 2032
rect 65432 1989 65441 2023
rect 65441 1989 65475 2023
rect 65475 1989 65484 2023
rect 65432 1980 65484 1989
rect 66168 1980 66220 2032
rect 66352 1955 66404 1964
rect 66352 1921 66361 1955
rect 66361 1921 66395 1955
rect 66395 1921 66404 1955
rect 66352 1912 66404 1921
rect 89904 1980 89956 2032
rect 71504 1955 71556 1964
rect 71504 1921 71513 1955
rect 71513 1921 71547 1955
rect 71547 1921 71556 1955
rect 71504 1912 71556 1921
rect 72240 1955 72292 1964
rect 72240 1921 72249 1955
rect 72249 1921 72283 1955
rect 72283 1921 72292 1955
rect 72240 1912 72292 1921
rect 73620 1912 73672 1964
rect 73712 1955 73764 1964
rect 73712 1921 73721 1955
rect 73721 1921 73755 1955
rect 73755 1921 73764 1955
rect 73712 1912 73764 1921
rect 65064 1887 65116 1896
rect 65064 1853 65073 1887
rect 65073 1853 65107 1887
rect 65107 1853 65116 1887
rect 65064 1844 65116 1853
rect 55588 1776 55640 1828
rect 22008 1708 22060 1760
rect 22100 1708 22152 1760
rect 22560 1708 22612 1760
rect 24124 1708 24176 1760
rect 25044 1751 25096 1760
rect 25044 1717 25053 1751
rect 25053 1717 25087 1751
rect 25087 1717 25096 1751
rect 25044 1708 25096 1717
rect 25964 1751 26016 1760
rect 25964 1717 25973 1751
rect 25973 1717 26007 1751
rect 26007 1717 26016 1751
rect 25964 1708 26016 1717
rect 27988 1708 28040 1760
rect 28816 1708 28868 1760
rect 30380 1751 30432 1760
rect 30380 1717 30389 1751
rect 30389 1717 30423 1751
rect 30423 1717 30432 1751
rect 30380 1708 30432 1717
rect 31024 1708 31076 1760
rect 32312 1708 32364 1760
rect 33140 1708 33192 1760
rect 35164 1751 35216 1760
rect 35164 1717 35173 1751
rect 35173 1717 35207 1751
rect 35207 1717 35216 1751
rect 35164 1708 35216 1717
rect 40408 1751 40460 1760
rect 40408 1717 40417 1751
rect 40417 1717 40451 1751
rect 40451 1717 40460 1751
rect 40408 1708 40460 1717
rect 52920 1751 52972 1760
rect 52920 1717 52929 1751
rect 52929 1717 52963 1751
rect 52963 1717 52972 1751
rect 52920 1708 52972 1717
rect 54300 1751 54352 1760
rect 54300 1717 54309 1751
rect 54309 1717 54343 1751
rect 54343 1717 54352 1751
rect 54300 1708 54352 1717
rect 55036 1751 55088 1760
rect 55036 1717 55045 1751
rect 55045 1717 55079 1751
rect 55079 1717 55088 1751
rect 55036 1708 55088 1717
rect 56232 1708 56284 1760
rect 56968 1708 57020 1760
rect 58256 1751 58308 1760
rect 58256 1717 58265 1751
rect 58265 1717 58299 1751
rect 58299 1717 58308 1751
rect 58256 1708 58308 1717
rect 59820 1708 59872 1760
rect 60740 1708 60792 1760
rect 63684 1708 63736 1760
rect 64420 1751 64472 1760
rect 64420 1717 64429 1751
rect 64429 1717 64463 1751
rect 64463 1717 64472 1751
rect 64420 1708 64472 1717
rect 67272 1751 67324 1760
rect 67272 1717 67281 1751
rect 67281 1717 67315 1751
rect 67315 1717 67324 1751
rect 67272 1708 67324 1717
rect 72056 1819 72108 1828
rect 72056 1785 72065 1819
rect 72065 1785 72099 1819
rect 72099 1785 72108 1819
rect 72056 1776 72108 1785
rect 73436 1776 73488 1828
rect 73344 1708 73396 1760
rect 75736 1887 75788 1896
rect 75736 1853 75745 1887
rect 75745 1853 75779 1887
rect 75779 1853 75788 1887
rect 75736 1844 75788 1853
rect 78588 1912 78640 1964
rect 77208 1887 77260 1896
rect 77208 1853 77217 1887
rect 77217 1853 77251 1887
rect 77251 1853 77260 1887
rect 77208 1844 77260 1853
rect 77484 1887 77536 1896
rect 77484 1853 77493 1887
rect 77493 1853 77527 1887
rect 77527 1853 77536 1887
rect 77484 1844 77536 1853
rect 79416 1887 79468 1896
rect 79416 1853 79425 1887
rect 79425 1853 79459 1887
rect 79459 1853 79468 1887
rect 79416 1844 79468 1853
rect 80888 1887 80940 1896
rect 80888 1853 80897 1887
rect 80897 1853 80931 1887
rect 80931 1853 80940 1887
rect 80888 1844 80940 1853
rect 81164 1955 81216 1964
rect 81164 1921 81173 1955
rect 81173 1921 81207 1955
rect 81207 1921 81216 1955
rect 81164 1912 81216 1921
rect 82360 1887 82412 1896
rect 82360 1853 82369 1887
rect 82369 1853 82403 1887
rect 82403 1853 82412 1887
rect 82360 1844 82412 1853
rect 82636 1887 82688 1896
rect 82636 1853 82645 1887
rect 82645 1853 82679 1887
rect 82679 1853 82688 1887
rect 82636 1844 82688 1853
rect 84568 1887 84620 1896
rect 84568 1853 84577 1887
rect 84577 1853 84611 1887
rect 84611 1853 84620 1887
rect 84568 1844 84620 1853
rect 84844 1955 84896 1964
rect 84844 1921 84853 1955
rect 84853 1921 84887 1955
rect 84887 1921 84896 1955
rect 84844 1912 84896 1921
rect 86040 1887 86092 1896
rect 86040 1853 86049 1887
rect 86049 1853 86083 1887
rect 86083 1853 86092 1887
rect 86040 1844 86092 1853
rect 86868 1912 86920 1964
rect 88248 1912 88300 1964
rect 89076 1955 89128 1964
rect 89076 1921 89085 1955
rect 89085 1921 89119 1955
rect 89119 1921 89128 1955
rect 91008 1980 91060 2032
rect 93768 1980 93820 2032
rect 97908 2048 97960 2100
rect 98736 2091 98788 2100
rect 98736 2057 98745 2091
rect 98745 2057 98779 2091
rect 98779 2057 98788 2091
rect 98736 2048 98788 2057
rect 98828 2048 98880 2100
rect 99932 1980 99984 2032
rect 101036 1980 101088 2032
rect 89076 1912 89128 1921
rect 88524 1844 88576 1896
rect 89628 1844 89680 1896
rect 89904 1887 89956 1896
rect 89904 1853 89913 1887
rect 89913 1853 89947 1887
rect 89947 1853 89956 1887
rect 89904 1844 89956 1853
rect 90732 1844 90784 1896
rect 91652 1955 91704 1964
rect 91652 1921 91661 1955
rect 91661 1921 91695 1955
rect 91695 1921 91704 1955
rect 91652 1912 91704 1921
rect 92572 1955 92624 1964
rect 92572 1921 92581 1955
rect 92581 1921 92615 1955
rect 92615 1921 92624 1955
rect 92572 1912 92624 1921
rect 93124 1912 93176 1964
rect 92388 1887 92440 1896
rect 92388 1853 92397 1887
rect 92397 1853 92431 1887
rect 92431 1853 92440 1887
rect 92388 1844 92440 1853
rect 93492 1844 93544 1896
rect 94228 1955 94280 1964
rect 94228 1921 94237 1955
rect 94237 1921 94271 1955
rect 94271 1921 94280 1955
rect 94228 1912 94280 1921
rect 95056 1844 95108 1896
rect 95884 1912 95936 1964
rect 95608 1844 95660 1896
rect 96344 1912 96396 1964
rect 96896 1955 96948 1964
rect 96896 1921 96905 1955
rect 96905 1921 96939 1955
rect 96939 1921 96948 1955
rect 96896 1912 96948 1921
rect 97834 1955 97886 1964
rect 97834 1921 97843 1955
rect 97843 1921 97877 1955
rect 97877 1921 97886 1955
rect 97834 1912 97886 1921
rect 97080 1887 97132 1896
rect 97080 1853 97089 1887
rect 97089 1853 97123 1887
rect 97123 1853 97132 1887
rect 97080 1844 97132 1853
rect 98092 1955 98144 1964
rect 98092 1921 98101 1955
rect 98101 1921 98135 1955
rect 98135 1921 98144 1955
rect 98092 1912 98144 1921
rect 107660 2048 107712 2100
rect 107752 2048 107804 2100
rect 108764 2048 108816 2100
rect 110880 2048 110932 2100
rect 107936 1980 107988 2032
rect 108304 1980 108356 2032
rect 110328 1980 110380 2032
rect 112536 2091 112588 2100
rect 112536 2057 112545 2091
rect 112545 2057 112579 2091
rect 112579 2057 112588 2091
rect 112536 2048 112588 2057
rect 114560 2048 114612 2100
rect 118976 2048 119028 2100
rect 120724 2048 120776 2100
rect 121092 2091 121144 2100
rect 121092 2057 121101 2091
rect 121101 2057 121135 2091
rect 121135 2057 121144 2091
rect 121092 2048 121144 2057
rect 124312 2091 124364 2100
rect 124312 2057 124321 2091
rect 124321 2057 124355 2091
rect 124355 2057 124364 2091
rect 124312 2048 124364 2057
rect 126704 2091 126756 2100
rect 126704 2057 126713 2091
rect 126713 2057 126747 2091
rect 126747 2057 126756 2091
rect 126704 2048 126756 2057
rect 128360 2091 128412 2100
rect 128360 2057 128369 2091
rect 128369 2057 128403 2091
rect 128403 2057 128412 2091
rect 128360 2048 128412 2057
rect 117136 1980 117188 2032
rect 117228 2023 117280 2032
rect 117228 1989 117237 2023
rect 117237 1989 117271 2023
rect 117271 1989 117280 2023
rect 117228 1980 117280 1989
rect 104900 1955 104952 1964
rect 104900 1921 104909 1955
rect 104909 1921 104943 1955
rect 104943 1921 104952 1955
rect 104900 1912 104952 1921
rect 105820 1955 105872 1964
rect 105820 1921 105829 1955
rect 105829 1921 105863 1955
rect 105863 1921 105872 1955
rect 105820 1912 105872 1921
rect 106004 1912 106056 1964
rect 106096 1955 106148 1964
rect 106096 1921 106105 1955
rect 106105 1921 106139 1955
rect 106139 1921 106148 1955
rect 106096 1912 106148 1921
rect 110236 1912 110288 1964
rect 110512 1912 110564 1964
rect 111892 1955 111944 1964
rect 111892 1921 111901 1955
rect 111901 1921 111935 1955
rect 111935 1921 111944 1955
rect 111892 1912 111944 1921
rect 74632 1776 74684 1828
rect 94044 1776 94096 1828
rect 94780 1776 94832 1828
rect 97448 1776 97500 1828
rect 99288 1887 99340 1896
rect 99288 1853 99297 1887
rect 99297 1853 99331 1887
rect 99331 1853 99340 1887
rect 99288 1844 99340 1853
rect 101128 1844 101180 1896
rect 105084 1887 105136 1896
rect 105084 1853 105093 1887
rect 105093 1853 105127 1887
rect 105127 1853 105136 1887
rect 105084 1844 105136 1853
rect 81440 1708 81492 1760
rect 88340 1751 88392 1760
rect 88340 1717 88349 1751
rect 88349 1717 88383 1751
rect 88383 1717 88392 1751
rect 88340 1708 88392 1717
rect 89904 1708 89956 1760
rect 91376 1708 91428 1760
rect 91652 1708 91704 1760
rect 92940 1708 92992 1760
rect 94596 1708 94648 1760
rect 103244 1776 103296 1828
rect 104164 1776 104216 1828
rect 107660 1887 107712 1896
rect 107660 1853 107669 1887
rect 107669 1853 107703 1887
rect 107703 1853 107712 1887
rect 107660 1844 107712 1853
rect 109132 1844 109184 1896
rect 101680 1708 101732 1760
rect 108580 1776 108632 1828
rect 107844 1708 107896 1760
rect 107936 1708 107988 1760
rect 110880 1887 110932 1896
rect 110880 1853 110889 1887
rect 110889 1853 110923 1887
rect 110923 1853 110932 1887
rect 110880 1844 110932 1853
rect 111340 1819 111392 1828
rect 111340 1785 111349 1819
rect 111349 1785 111383 1819
rect 111383 1785 111392 1819
rect 111340 1776 111392 1785
rect 114836 1844 114888 1896
rect 115020 1887 115072 1896
rect 115020 1853 115029 1887
rect 115029 1853 115063 1887
rect 115063 1853 115072 1887
rect 115020 1844 115072 1853
rect 115204 1887 115256 1896
rect 115204 1853 115213 1887
rect 115213 1853 115247 1887
rect 115247 1853 115256 1887
rect 115204 1844 115256 1853
rect 115940 1955 115992 1964
rect 115940 1921 115949 1955
rect 115949 1921 115983 1955
rect 115983 1921 115992 1955
rect 115940 1912 115992 1921
rect 116032 1955 116084 1964
rect 116032 1921 116066 1955
rect 116066 1921 116084 1955
rect 116032 1912 116084 1921
rect 116216 1955 116268 1964
rect 116216 1921 116225 1955
rect 116225 1921 116259 1955
rect 116259 1921 116268 1955
rect 116216 1912 116268 1921
rect 117412 1912 117464 1964
rect 117688 1955 117740 1964
rect 117688 1921 117697 1955
rect 117697 1921 117731 1955
rect 117731 1921 117740 1955
rect 117688 1912 117740 1921
rect 115572 1844 115624 1896
rect 118148 1887 118200 1896
rect 115664 1819 115716 1828
rect 115664 1785 115673 1819
rect 115673 1785 115707 1819
rect 115707 1785 115716 1819
rect 115664 1776 115716 1785
rect 111984 1708 112036 1760
rect 118148 1853 118157 1887
rect 118157 1853 118191 1887
rect 118191 1853 118200 1887
rect 118148 1844 118200 1853
rect 120172 1912 120224 1964
rect 120724 1955 120776 1964
rect 120724 1921 120733 1955
rect 120733 1921 120767 1955
rect 120767 1921 120776 1955
rect 120724 1912 120776 1921
rect 121736 1980 121788 2032
rect 131764 2023 131816 2032
rect 131764 1989 131773 2023
rect 131773 1989 131807 2023
rect 131807 1989 131816 2023
rect 131764 1980 131816 1989
rect 133696 2091 133748 2100
rect 133696 2057 133705 2091
rect 133705 2057 133739 2091
rect 133739 2057 133748 2091
rect 133696 2048 133748 2057
rect 139492 2048 139544 2100
rect 139952 2048 140004 2100
rect 121460 1955 121512 1964
rect 121460 1921 121469 1955
rect 121469 1921 121503 1955
rect 121503 1921 121512 1955
rect 121460 1912 121512 1921
rect 122656 1912 122708 1964
rect 124956 1912 125008 1964
rect 125048 1912 125100 1964
rect 118148 1708 118200 1760
rect 118516 1887 118568 1896
rect 118516 1853 118550 1887
rect 118550 1853 118568 1887
rect 118516 1844 118568 1853
rect 119068 1844 119120 1896
rect 122104 1887 122156 1896
rect 122104 1853 122113 1887
rect 122113 1853 122147 1887
rect 122147 1853 122156 1887
rect 122104 1844 122156 1853
rect 122840 1887 122892 1896
rect 122840 1853 122849 1887
rect 122849 1853 122883 1887
rect 122883 1853 122892 1887
rect 123116 1887 123168 1896
rect 122840 1844 122892 1853
rect 123116 1853 123125 1887
rect 123125 1853 123159 1887
rect 123159 1853 123168 1887
rect 123116 1844 123168 1853
rect 124036 1844 124088 1896
rect 126336 1955 126388 1964
rect 126336 1921 126345 1955
rect 126345 1921 126379 1955
rect 126379 1921 126388 1955
rect 126336 1912 126388 1921
rect 126428 1844 126480 1896
rect 127440 1844 127492 1896
rect 127992 1955 128044 1964
rect 127992 1921 128001 1955
rect 128001 1921 128035 1955
rect 128035 1921 128044 1955
rect 127992 1912 128044 1921
rect 128820 1955 128872 1964
rect 128820 1921 128829 1955
rect 128829 1921 128863 1955
rect 128863 1921 128872 1955
rect 128820 1912 128872 1921
rect 130108 1912 130160 1964
rect 129096 1887 129148 1896
rect 129096 1853 129105 1887
rect 129105 1853 129139 1887
rect 129139 1853 129148 1887
rect 129096 1844 129148 1853
rect 129648 1844 129700 1896
rect 131120 1912 131172 1964
rect 131856 1912 131908 1964
rect 138940 1980 138992 2032
rect 132592 1912 132644 1964
rect 133420 1912 133472 1964
rect 134340 1955 134392 1964
rect 134340 1921 134349 1955
rect 134349 1921 134383 1955
rect 134383 1921 134392 1955
rect 134340 1912 134392 1921
rect 135352 1955 135404 1964
rect 135352 1921 135361 1955
rect 135361 1921 135395 1955
rect 135395 1921 135404 1955
rect 135352 1912 135404 1921
rect 139032 1912 139084 1964
rect 140228 1980 140280 2032
rect 139768 1955 139820 1964
rect 139768 1921 139777 1955
rect 139777 1921 139811 1955
rect 139811 1921 139820 1955
rect 139768 1912 139820 1921
rect 140504 1955 140556 1964
rect 140504 1921 140513 1955
rect 140513 1921 140547 1955
rect 140547 1921 140556 1955
rect 140504 1912 140556 1921
rect 140872 2048 140924 2100
rect 141700 2048 141752 2100
rect 142344 2091 142396 2100
rect 142344 2057 142353 2091
rect 142353 2057 142387 2091
rect 142387 2057 142396 2091
rect 142344 2048 142396 2057
rect 144644 2091 144696 2100
rect 144644 2057 144653 2091
rect 144653 2057 144687 2091
rect 144687 2057 144696 2091
rect 144644 2048 144696 2057
rect 145748 2048 145800 2100
rect 147404 2048 147456 2100
rect 148600 2048 148652 2100
rect 152096 2048 152148 2100
rect 152556 2048 152608 2100
rect 152740 2048 152792 2100
rect 153844 2048 153896 2100
rect 153936 2048 153988 2100
rect 154948 2048 155000 2100
rect 159088 2048 159140 2100
rect 134156 1887 134208 1896
rect 134156 1853 134165 1887
rect 134165 1853 134199 1887
rect 134199 1853 134208 1887
rect 134156 1844 134208 1853
rect 141424 1955 141476 1964
rect 141424 1921 141433 1955
rect 141433 1921 141467 1955
rect 141467 1921 141476 1955
rect 141424 1912 141476 1921
rect 141700 1955 141752 1964
rect 141700 1921 141709 1955
rect 141709 1921 141743 1955
rect 141743 1921 141752 1955
rect 141700 1912 141752 1921
rect 142804 1955 142856 1964
rect 142804 1921 142813 1955
rect 142813 1921 142847 1955
rect 142847 1921 142856 1955
rect 142804 1912 142856 1921
rect 143724 1955 143776 1964
rect 143724 1921 143733 1955
rect 143733 1921 143767 1955
rect 143767 1921 143776 1955
rect 143724 1912 143776 1921
rect 143908 1912 143960 1964
rect 145196 1912 145248 1964
rect 146576 1955 146628 1964
rect 146576 1921 146585 1955
rect 146585 1921 146619 1955
rect 146619 1921 146628 1955
rect 146576 1912 146628 1921
rect 150624 1912 150676 1964
rect 151728 1955 151780 1964
rect 151728 1921 151737 1955
rect 151737 1921 151771 1955
rect 151771 1921 151780 1955
rect 151728 1912 151780 1921
rect 152004 1955 152056 1964
rect 152004 1921 152013 1955
rect 152013 1921 152047 1955
rect 152047 1921 152056 1955
rect 152004 1912 152056 1921
rect 153292 1955 153344 1964
rect 153292 1921 153301 1955
rect 153301 1921 153335 1955
rect 153335 1921 153344 1955
rect 153292 1912 153344 1921
rect 153384 1912 153436 1964
rect 154580 1955 154632 1964
rect 154580 1921 154589 1955
rect 154589 1921 154623 1955
rect 154623 1921 154632 1955
rect 154580 1912 154632 1921
rect 157340 1980 157392 2032
rect 158536 1980 158588 2032
rect 160192 2048 160244 2100
rect 160284 2091 160336 2100
rect 160284 2057 160293 2091
rect 160293 2057 160327 2091
rect 160327 2057 160336 2091
rect 160284 2048 160336 2057
rect 161480 2048 161532 2100
rect 163964 2091 164016 2100
rect 163964 2057 163973 2091
rect 163973 2057 164007 2091
rect 164007 2057 164016 2091
rect 163964 2048 164016 2057
rect 165620 2091 165672 2100
rect 165620 2057 165629 2091
rect 165629 2057 165663 2091
rect 165663 2057 165672 2091
rect 165620 2048 165672 2057
rect 165804 2048 165856 2100
rect 167460 2091 167512 2100
rect 167460 2057 167469 2091
rect 167469 2057 167503 2091
rect 167503 2057 167512 2091
rect 167460 2048 167512 2057
rect 190920 2091 190972 2100
rect 190920 2057 190929 2091
rect 190929 2057 190963 2091
rect 190963 2057 190972 2091
rect 190920 2048 190972 2057
rect 192208 2091 192260 2100
rect 192208 2057 192217 2091
rect 192217 2057 192251 2091
rect 192251 2057 192260 2091
rect 192208 2048 192260 2057
rect 156328 1912 156380 1964
rect 156788 1955 156840 1964
rect 156788 1921 156797 1955
rect 156797 1921 156831 1955
rect 156831 1921 156840 1955
rect 156788 1912 156840 1921
rect 158996 1912 159048 1964
rect 159272 1955 159324 1964
rect 159272 1921 159281 1955
rect 159281 1921 159315 1955
rect 159315 1921 159324 1955
rect 159272 1912 159324 1921
rect 160008 1912 160060 1964
rect 161112 1955 161164 1964
rect 161112 1921 161121 1955
rect 161121 1921 161155 1955
rect 161155 1921 161164 1955
rect 161112 1912 161164 1921
rect 161572 1912 161624 1964
rect 162400 1980 162452 2032
rect 162676 1912 162728 1964
rect 163596 1955 163648 1964
rect 163596 1921 163605 1955
rect 163605 1921 163639 1955
rect 163639 1921 163648 1955
rect 163596 1912 163648 1921
rect 141056 1844 141108 1896
rect 141608 1844 141660 1896
rect 139032 1776 139084 1828
rect 118608 1708 118660 1760
rect 120540 1751 120592 1760
rect 120540 1717 120549 1751
rect 120549 1717 120583 1751
rect 120583 1717 120592 1751
rect 120540 1708 120592 1717
rect 121644 1708 121696 1760
rect 122472 1751 122524 1760
rect 122472 1717 122481 1751
rect 122481 1717 122515 1751
rect 122515 1717 122524 1751
rect 122472 1708 122524 1717
rect 123208 1708 123260 1760
rect 125784 1751 125836 1760
rect 125784 1717 125793 1751
rect 125793 1717 125827 1751
rect 125827 1717 125836 1751
rect 125784 1708 125836 1717
rect 127624 1708 127676 1760
rect 130660 1708 130712 1760
rect 132684 1751 132736 1760
rect 132684 1717 132693 1751
rect 132693 1717 132727 1751
rect 132727 1717 132736 1751
rect 132684 1708 132736 1717
rect 134340 1708 134392 1760
rect 135260 1708 135312 1760
rect 140228 1708 140280 1760
rect 140688 1708 140740 1760
rect 140872 1708 140924 1760
rect 142436 1708 142488 1760
rect 144184 1844 144236 1896
rect 146392 1844 146444 1896
rect 146668 1844 146720 1896
rect 146852 1887 146904 1896
rect 146852 1853 146861 1887
rect 146861 1853 146895 1887
rect 146895 1853 146904 1887
rect 146852 1844 146904 1853
rect 143448 1819 143500 1828
rect 143448 1785 143457 1819
rect 143457 1785 143491 1819
rect 143491 1785 143500 1819
rect 143448 1776 143500 1785
rect 146300 1819 146352 1828
rect 146300 1785 146309 1819
rect 146309 1785 146343 1819
rect 146343 1785 146352 1819
rect 146300 1776 146352 1785
rect 144828 1708 144880 1760
rect 148508 1844 148560 1896
rect 148692 1844 148744 1896
rect 148968 1887 149020 1896
rect 148968 1853 149002 1887
rect 149002 1853 149020 1887
rect 148968 1844 149020 1853
rect 149336 1844 149388 1896
rect 149704 1844 149756 1896
rect 151544 1844 151596 1896
rect 150624 1776 150676 1828
rect 151268 1708 151320 1760
rect 151452 1819 151504 1828
rect 151452 1785 151461 1819
rect 151461 1785 151495 1819
rect 151495 1785 151504 1819
rect 151452 1776 151504 1785
rect 156604 1844 156656 1896
rect 157156 1844 157208 1896
rect 159180 1844 159232 1896
rect 162860 1844 162912 1896
rect 164516 1955 164568 1964
rect 164516 1921 164525 1955
rect 164525 1921 164559 1955
rect 164559 1921 164568 1955
rect 164516 1912 164568 1921
rect 165160 1912 165212 1964
rect 166264 1955 166316 1964
rect 166264 1921 166273 1955
rect 166273 1921 166307 1955
rect 166307 1921 166316 1955
rect 166264 1912 166316 1921
rect 167184 1980 167236 2032
rect 167092 1955 167144 1964
rect 167092 1921 167101 1955
rect 167101 1921 167135 1955
rect 167135 1921 167144 1955
rect 167092 1912 167144 1921
rect 173808 1980 173860 2032
rect 168012 1912 168064 1964
rect 169760 1912 169812 1964
rect 176844 1955 176896 1964
rect 176844 1921 176853 1955
rect 176853 1921 176887 1955
rect 176887 1921 176896 1955
rect 176844 1912 176896 1921
rect 179420 1955 179472 1964
rect 179420 1921 179429 1955
rect 179429 1921 179463 1955
rect 179463 1921 179472 1955
rect 179420 1912 179472 1921
rect 182088 1980 182140 2032
rect 184572 1955 184624 1964
rect 184572 1921 184581 1955
rect 184581 1921 184615 1955
rect 184615 1921 184624 1955
rect 184572 1912 184624 1921
rect 187148 1955 187200 1964
rect 187148 1921 187157 1955
rect 187157 1921 187191 1955
rect 187191 1921 187200 1955
rect 187148 1912 187200 1921
rect 190644 1980 190696 2032
rect 191012 1912 191064 1964
rect 166540 1844 166592 1896
rect 167828 1844 167880 1896
rect 172980 1887 173032 1896
rect 172980 1853 172989 1887
rect 172989 1853 173023 1887
rect 173023 1853 173032 1887
rect 172980 1844 173032 1853
rect 174452 1887 174504 1896
rect 174452 1853 174461 1887
rect 174461 1853 174495 1887
rect 174495 1853 174504 1887
rect 174452 1844 174504 1853
rect 174728 1887 174780 1896
rect 174728 1853 174737 1887
rect 174737 1853 174771 1887
rect 174771 1853 174780 1887
rect 174728 1844 174780 1853
rect 176568 1887 176620 1896
rect 176568 1853 176577 1887
rect 176577 1853 176611 1887
rect 176611 1853 176620 1887
rect 176568 1844 176620 1853
rect 177856 1887 177908 1896
rect 177856 1853 177865 1887
rect 177865 1853 177899 1887
rect 177899 1853 177908 1887
rect 177856 1844 177908 1853
rect 178132 1887 178184 1896
rect 178132 1853 178141 1887
rect 178141 1853 178175 1887
rect 178175 1853 178184 1887
rect 178132 1844 178184 1853
rect 179144 1887 179196 1896
rect 179144 1853 179153 1887
rect 179153 1853 179187 1887
rect 179187 1853 179196 1887
rect 179144 1844 179196 1853
rect 181720 1887 181772 1896
rect 181720 1853 181729 1887
rect 181729 1853 181763 1887
rect 181763 1853 181772 1887
rect 181720 1844 181772 1853
rect 183008 1887 183060 1896
rect 183008 1853 183017 1887
rect 183017 1853 183051 1887
rect 183051 1853 183060 1887
rect 183008 1844 183060 1853
rect 184296 1887 184348 1896
rect 184296 1853 184305 1887
rect 184305 1853 184339 1887
rect 184339 1853 184348 1887
rect 184296 1844 184348 1853
rect 186320 1844 186372 1896
rect 188160 1887 188212 1896
rect 188160 1853 188169 1887
rect 188169 1853 188203 1887
rect 188203 1853 188212 1887
rect 188160 1844 188212 1853
rect 191840 1887 191892 1896
rect 191840 1853 191849 1887
rect 191849 1853 191883 1887
rect 191883 1853 191892 1887
rect 191840 1844 191892 1853
rect 192852 1887 192904 1896
rect 192852 1853 192861 1887
rect 192861 1853 192895 1887
rect 192895 1853 192904 1887
rect 192852 1844 192904 1853
rect 193496 1912 193548 1964
rect 195336 1955 195388 1964
rect 195336 1921 195345 1955
rect 195345 1921 195379 1955
rect 195379 1921 195388 1955
rect 195336 1912 195388 1921
rect 195704 1955 195756 1964
rect 195704 1921 195713 1955
rect 195713 1921 195747 1955
rect 195747 1921 195756 1955
rect 195704 1912 195756 1921
rect 195980 1912 196032 1964
rect 196440 1980 196492 2032
rect 197544 2091 197596 2100
rect 197544 2057 197553 2091
rect 197553 2057 197587 2091
rect 197587 2057 197596 2091
rect 197544 2048 197596 2057
rect 199752 2091 199804 2100
rect 199752 2057 199761 2091
rect 199761 2057 199795 2091
rect 199795 2057 199804 2091
rect 199752 2048 199804 2057
rect 216588 2048 216640 2100
rect 216680 2048 216732 2100
rect 218428 2048 218480 2100
rect 197176 1955 197228 1964
rect 197176 1921 197185 1955
rect 197185 1921 197219 1955
rect 197219 1921 197228 1955
rect 197176 1912 197228 1921
rect 200212 1980 200264 2032
rect 202696 2023 202748 2032
rect 202696 1989 202705 2023
rect 202705 1989 202739 2023
rect 202739 1989 202748 2023
rect 202696 1980 202748 1989
rect 199384 1955 199436 1964
rect 199384 1921 199393 1955
rect 199393 1921 199427 1955
rect 199427 1921 199436 1955
rect 199384 1912 199436 1921
rect 194784 1844 194836 1896
rect 191196 1776 191248 1828
rect 198372 1887 198424 1896
rect 198372 1853 198381 1887
rect 198381 1853 198415 1887
rect 198415 1853 198424 1887
rect 200304 1955 200356 1964
rect 200304 1921 200313 1955
rect 200313 1921 200347 1955
rect 200347 1921 200356 1955
rect 200304 1912 200356 1921
rect 200672 1912 200724 1964
rect 202328 1955 202380 1964
rect 202328 1921 202337 1955
rect 202337 1921 202371 1955
rect 202371 1921 202380 1955
rect 202328 1912 202380 1921
rect 198372 1844 198424 1853
rect 201500 1844 201552 1896
rect 203248 1955 203300 1964
rect 203248 1921 203257 1955
rect 203257 1921 203291 1955
rect 203291 1921 203300 1955
rect 203248 1912 203300 1921
rect 209688 1980 209740 2032
rect 210700 1980 210752 2032
rect 202788 1844 202840 1896
rect 208492 1955 208544 1964
rect 208492 1921 208501 1955
rect 208501 1921 208535 1955
rect 208535 1921 208544 1955
rect 208492 1912 208544 1921
rect 208952 1955 209004 1964
rect 208952 1921 208961 1955
rect 208961 1921 208995 1955
rect 208995 1921 209004 1955
rect 208952 1912 209004 1921
rect 211344 1955 211396 1964
rect 211344 1921 211353 1955
rect 211353 1921 211387 1955
rect 211387 1921 211396 1955
rect 211344 1912 211396 1921
rect 211436 1955 211488 1964
rect 211436 1921 211445 1955
rect 211445 1921 211479 1955
rect 211479 1921 211488 1955
rect 211436 1912 211488 1921
rect 211620 1955 211672 1964
rect 211620 1921 211629 1955
rect 211629 1921 211663 1955
rect 211663 1921 211672 1955
rect 211620 1912 211672 1921
rect 211988 2023 212040 2032
rect 211988 1989 211997 2023
rect 211997 1989 212031 2023
rect 212031 1989 212040 2023
rect 211988 1980 212040 1989
rect 214472 2023 214524 2032
rect 214472 1989 214481 2023
rect 214481 1989 214515 2023
rect 214515 1989 214524 2023
rect 214472 1980 214524 1989
rect 219624 2091 219676 2100
rect 219624 2057 219633 2091
rect 219633 2057 219667 2091
rect 219667 2057 219676 2091
rect 219624 2048 219676 2057
rect 220728 2048 220780 2100
rect 221372 2048 221424 2100
rect 222660 2048 222712 2100
rect 224132 2091 224184 2100
rect 224132 2057 224141 2091
rect 224141 2057 224175 2091
rect 224175 2057 224184 2091
rect 224132 2048 224184 2057
rect 224500 2091 224552 2100
rect 224500 2057 224509 2091
rect 224509 2057 224543 2091
rect 224543 2057 224552 2091
rect 224500 2048 224552 2057
rect 225788 2091 225840 2100
rect 225788 2057 225797 2091
rect 225797 2057 225831 2091
rect 225831 2057 225840 2091
rect 225788 2048 225840 2057
rect 226800 2091 226852 2100
rect 226800 2057 226809 2091
rect 226809 2057 226843 2091
rect 226843 2057 226852 2091
rect 226800 2048 226852 2057
rect 228456 2091 228508 2100
rect 228456 2057 228465 2091
rect 228465 2057 228499 2091
rect 228499 2057 228508 2091
rect 228456 2048 228508 2057
rect 230940 2091 230992 2100
rect 230940 2057 230949 2091
rect 230949 2057 230983 2091
rect 230983 2057 230992 2091
rect 230940 2048 230992 2057
rect 231768 2091 231820 2100
rect 231768 2057 231777 2091
rect 231777 2057 231811 2091
rect 231811 2057 231820 2091
rect 231768 2048 231820 2057
rect 232596 2091 232648 2100
rect 232596 2057 232605 2091
rect 232605 2057 232639 2091
rect 232639 2057 232648 2091
rect 232596 2048 232648 2057
rect 232964 2048 233016 2100
rect 234988 2048 235040 2100
rect 236920 2091 236972 2100
rect 236920 2057 236929 2091
rect 236929 2057 236963 2091
rect 236963 2057 236972 2091
rect 236920 2048 236972 2057
rect 237012 2048 237064 2100
rect 213644 1955 213696 1964
rect 213644 1921 213678 1955
rect 213678 1921 213696 1955
rect 213644 1912 213696 1921
rect 213828 1955 213880 1964
rect 213828 1921 213837 1955
rect 213837 1921 213871 1955
rect 213871 1921 213880 1955
rect 213828 1912 213880 1921
rect 208308 1844 208360 1896
rect 209780 1887 209832 1896
rect 209780 1853 209789 1887
rect 209789 1853 209823 1887
rect 209823 1853 209832 1887
rect 209780 1844 209832 1853
rect 213092 1776 213144 1828
rect 213368 1844 213420 1896
rect 214656 1912 214708 1964
rect 221832 1980 221884 2032
rect 226432 1980 226484 2032
rect 154580 1708 154632 1760
rect 155960 1751 156012 1760
rect 155960 1717 155969 1751
rect 155969 1717 156003 1751
rect 156003 1717 156012 1751
rect 155960 1708 156012 1717
rect 161480 1751 161532 1760
rect 161480 1717 161489 1751
rect 161489 1717 161523 1751
rect 161523 1717 161532 1751
rect 161480 1708 161532 1717
rect 163136 1751 163188 1760
rect 163136 1717 163145 1751
rect 163145 1717 163179 1751
rect 163179 1717 163188 1751
rect 163136 1708 163188 1717
rect 164424 1708 164476 1760
rect 168380 1708 168432 1760
rect 193220 1751 193272 1760
rect 193220 1717 193229 1751
rect 193229 1717 193263 1751
rect 193263 1717 193272 1751
rect 193220 1708 193272 1717
rect 194048 1751 194100 1760
rect 194048 1717 194057 1751
rect 194057 1717 194091 1751
rect 194091 1717 194100 1751
rect 194048 1708 194100 1717
rect 194600 1708 194652 1760
rect 196072 1708 196124 1760
rect 200580 1751 200632 1760
rect 200580 1717 200589 1751
rect 200589 1717 200623 1751
rect 200623 1717 200632 1751
rect 200580 1708 200632 1717
rect 202880 1708 202932 1760
rect 210240 1708 210292 1760
rect 210700 1708 210752 1760
rect 213736 1708 213788 1760
rect 215852 1955 215904 1964
rect 215852 1921 215861 1955
rect 215861 1921 215895 1955
rect 215895 1921 215904 1955
rect 215852 1912 215904 1921
rect 216036 1912 216088 1964
rect 218704 1955 218756 1964
rect 218704 1921 218713 1955
rect 218713 1921 218747 1955
rect 218747 1921 218756 1955
rect 218704 1912 218756 1921
rect 218980 1955 219032 1964
rect 218980 1921 218989 1955
rect 218989 1921 219023 1955
rect 219023 1921 219032 1955
rect 218980 1912 219032 1921
rect 220176 1912 220228 1964
rect 221004 1955 221056 1962
rect 221004 1921 221031 1955
rect 221031 1921 221056 1955
rect 221004 1910 221056 1921
rect 221280 1955 221332 1964
rect 221280 1921 221289 1955
rect 221289 1921 221323 1955
rect 221323 1921 221332 1955
rect 221280 1912 221332 1921
rect 222016 1912 222068 1964
rect 224408 1912 224460 1964
rect 215484 1844 215536 1896
rect 216128 1887 216180 1896
rect 216128 1853 216137 1887
rect 216137 1853 216171 1887
rect 216171 1853 216180 1887
rect 216128 1844 216180 1853
rect 215576 1819 215628 1828
rect 215576 1785 215585 1819
rect 215585 1785 215619 1819
rect 215619 1785 215628 1819
rect 215576 1776 215628 1785
rect 214840 1708 214892 1760
rect 219348 1844 219400 1896
rect 219532 1844 219584 1896
rect 220360 1844 220412 1896
rect 218152 1776 218204 1828
rect 219440 1776 219492 1828
rect 220452 1776 220504 1828
rect 223396 1844 223448 1896
rect 224500 1844 224552 1896
rect 225420 1887 225472 1896
rect 225420 1853 225429 1887
rect 225429 1853 225463 1887
rect 225463 1853 225472 1887
rect 225420 1844 225472 1853
rect 226432 1887 226484 1896
rect 226432 1853 226441 1887
rect 226441 1853 226475 1887
rect 226475 1853 226484 1887
rect 226432 1844 226484 1853
rect 227260 1955 227312 1964
rect 227260 1921 227269 1955
rect 227269 1921 227303 1955
rect 227303 1921 227312 1955
rect 227260 1912 227312 1921
rect 228364 1980 228416 2032
rect 229836 1980 229888 2032
rect 227076 1844 227128 1896
rect 228916 1955 228968 1964
rect 228916 1921 228925 1955
rect 228925 1921 228959 1955
rect 228959 1921 228968 1955
rect 228916 1912 228968 1921
rect 229744 1955 229796 1964
rect 229744 1921 229753 1955
rect 229753 1921 229787 1955
rect 229787 1921 229796 1955
rect 229744 1912 229796 1921
rect 229928 1955 229980 1964
rect 229928 1921 229937 1955
rect 229937 1921 229971 1955
rect 229971 1921 229980 1955
rect 229928 1912 229980 1921
rect 231492 1980 231544 2032
rect 230664 1955 230716 1964
rect 230664 1921 230673 1955
rect 230673 1921 230707 1955
rect 230707 1921 230716 1955
rect 230664 1912 230716 1921
rect 230756 1955 230808 1964
rect 230756 1921 230765 1955
rect 230765 1921 230799 1955
rect 230799 1921 230808 1955
rect 230756 1912 230808 1921
rect 230848 1912 230900 1964
rect 232044 1912 232096 1964
rect 232780 1912 232832 1964
rect 233608 1912 233660 1964
rect 235632 1912 235684 1964
rect 236184 1980 236236 2032
rect 236000 1912 236052 1964
rect 236092 1912 236144 1964
rect 239496 2048 239548 2100
rect 243636 2048 243688 2100
rect 245384 1980 245436 2032
rect 231676 1844 231728 1896
rect 233516 1844 233568 1896
rect 241244 1887 241296 1896
rect 241244 1853 241253 1887
rect 241253 1853 241287 1887
rect 241287 1853 241296 1887
rect 241244 1844 241296 1853
rect 242808 1844 242860 1896
rect 244832 1887 244884 1896
rect 244832 1853 244841 1887
rect 244841 1853 244875 1887
rect 244875 1853 244884 1887
rect 244832 1844 244884 1853
rect 245936 1844 245988 1896
rect 246672 1887 246724 1896
rect 246672 1853 246681 1887
rect 246681 1853 246715 1887
rect 246715 1853 246724 1887
rect 246672 1844 246724 1853
rect 219532 1708 219584 1760
rect 221372 1708 221424 1760
rect 221924 1708 221976 1760
rect 223396 1751 223448 1760
rect 223396 1717 223405 1751
rect 223405 1717 223439 1751
rect 223439 1717 223448 1751
rect 223396 1708 223448 1717
rect 225512 1708 225564 1760
rect 227444 1751 227496 1760
rect 227444 1717 227453 1751
rect 227453 1717 227487 1751
rect 227487 1717 227496 1751
rect 227444 1708 227496 1717
rect 228548 1708 228600 1760
rect 230112 1751 230164 1760
rect 230112 1717 230121 1751
rect 230121 1717 230155 1751
rect 230155 1717 230164 1751
rect 230112 1708 230164 1717
rect 233700 1708 233752 1760
rect 235264 1751 235316 1760
rect 235264 1717 235273 1751
rect 235273 1717 235307 1751
rect 235307 1717 235316 1751
rect 235264 1708 235316 1717
rect 237380 1708 237432 1760
rect 245752 1776 245804 1828
rect 247408 1955 247460 1964
rect 247408 1921 247417 1955
rect 247417 1921 247451 1955
rect 247451 1921 247460 1955
rect 247408 1912 247460 1921
rect 248880 2048 248932 2100
rect 252376 1980 252428 2032
rect 255228 1980 255280 2032
rect 260288 2048 260340 2100
rect 261116 2048 261168 2100
rect 263140 2048 263192 2100
rect 255688 2023 255740 2032
rect 255688 1989 255697 2023
rect 255697 1989 255731 2023
rect 255731 1989 255740 2023
rect 255688 1980 255740 1989
rect 268844 2048 268896 2100
rect 263968 1980 264020 2032
rect 268568 1980 268620 2032
rect 247500 1844 247552 1896
rect 250536 1887 250588 1896
rect 250536 1853 250545 1887
rect 250545 1853 250579 1887
rect 250579 1853 250588 1887
rect 250536 1844 250588 1853
rect 249800 1776 249852 1828
rect 251272 1887 251324 1896
rect 251272 1853 251281 1887
rect 251281 1853 251315 1887
rect 251315 1853 251324 1887
rect 251272 1844 251324 1853
rect 251364 1844 251416 1896
rect 252560 1708 252612 1760
rect 255688 1708 255740 1760
rect 258448 1912 258500 1964
rect 258540 1912 258592 1964
rect 260472 1955 260524 1964
rect 260472 1921 260481 1955
rect 260481 1921 260515 1955
rect 260515 1921 260524 1955
rect 260472 1912 260524 1921
rect 261392 1912 261444 1964
rect 261484 1955 261536 1964
rect 261484 1921 261493 1955
rect 261493 1921 261527 1955
rect 261527 1921 261536 1955
rect 261484 1912 261536 1921
rect 261760 1912 261812 1964
rect 258172 1844 258224 1896
rect 260196 1844 260248 1896
rect 262864 1912 262916 1964
rect 264060 1912 264112 1964
rect 264336 1955 264388 1964
rect 264336 1921 264345 1955
rect 264345 1921 264379 1955
rect 264379 1921 264388 1955
rect 264336 1912 264388 1921
rect 264428 1912 264480 1964
rect 265164 1955 265216 1964
rect 265164 1921 265173 1955
rect 265173 1921 265207 1955
rect 265207 1921 265216 1955
rect 265164 1912 265216 1921
rect 265808 1955 265860 1964
rect 265808 1921 265817 1955
rect 265817 1921 265851 1955
rect 265851 1921 265860 1955
rect 265808 1912 265860 1921
rect 266544 1912 266596 1964
rect 267004 1955 267056 1964
rect 267004 1921 267013 1955
rect 267013 1921 267047 1955
rect 267047 1921 267056 1955
rect 267004 1912 267056 1921
rect 267372 1912 267424 1964
rect 267740 1912 267792 1964
rect 269120 1912 269172 1964
rect 269948 1980 270000 2032
rect 271144 1776 271196 1828
rect 272156 1776 272208 1828
rect 257712 1708 257764 1760
rect 257988 1708 258040 1760
rect 263140 1708 263192 1760
rect 264152 1708 264204 1760
rect 265624 1708 265676 1760
rect 266728 1708 266780 1760
rect 267832 1751 267884 1760
rect 267832 1717 267841 1751
rect 267841 1717 267875 1751
rect 267875 1717 267884 1751
rect 267832 1708 267884 1717
rect 268200 1708 268252 1760
rect 269764 1708 269816 1760
rect 34748 1606 34800 1658
rect 34812 1606 34864 1658
rect 34876 1606 34928 1658
rect 34940 1606 34992 1658
rect 35004 1606 35056 1658
rect 102345 1606 102397 1658
rect 102409 1606 102461 1658
rect 102473 1606 102525 1658
rect 102537 1606 102589 1658
rect 102601 1606 102653 1658
rect 169942 1606 169994 1658
rect 170006 1606 170058 1658
rect 170070 1606 170122 1658
rect 170134 1606 170186 1658
rect 170198 1606 170250 1658
rect 237539 1606 237591 1658
rect 237603 1606 237655 1658
rect 237667 1606 237719 1658
rect 237731 1606 237783 1658
rect 237795 1606 237847 1658
rect 20720 1504 20772 1556
rect 25044 1504 25096 1556
rect 27436 1504 27488 1556
rect 27620 1504 27672 1556
rect 54300 1504 54352 1556
rect 58072 1504 58124 1556
rect 62212 1504 62264 1556
rect 73436 1504 73488 1556
rect 24768 1436 24820 1488
rect 22652 1368 22704 1420
rect 23756 1368 23808 1420
rect 25136 1368 25188 1420
rect 25688 1368 25740 1420
rect 27068 1368 27120 1420
rect 31300 1436 31352 1488
rect 65064 1436 65116 1488
rect 82636 1436 82688 1488
rect 92388 1436 92440 1488
rect 92848 1504 92900 1556
rect 95516 1504 95568 1556
rect 96988 1504 97040 1556
rect 53840 1368 53892 1420
rect 54300 1411 54352 1420
rect 54300 1377 54309 1411
rect 54309 1377 54343 1411
rect 54343 1377 54352 1411
rect 54300 1368 54352 1377
rect 58164 1368 58216 1420
rect 59544 1368 59596 1420
rect 62028 1411 62080 1420
rect 62028 1377 62037 1411
rect 62037 1377 62071 1411
rect 62071 1377 62080 1411
rect 62028 1368 62080 1377
rect 66076 1368 66128 1420
rect 69112 1411 69164 1420
rect 69112 1377 69121 1411
rect 69121 1377 69155 1411
rect 69155 1377 69164 1411
rect 69112 1368 69164 1377
rect 1952 1275 2004 1284
rect 1952 1241 1961 1275
rect 1961 1241 1995 1275
rect 1995 1241 2004 1275
rect 1952 1232 2004 1241
rect 2872 1343 2924 1352
rect 2872 1309 2881 1343
rect 2881 1309 2915 1343
rect 2915 1309 2924 1343
rect 2872 1300 2924 1309
rect 5356 1300 5408 1352
rect 5448 1343 5500 1352
rect 5448 1309 5457 1343
rect 5457 1309 5491 1343
rect 5491 1309 5500 1343
rect 5448 1300 5500 1309
rect 7748 1343 7800 1352
rect 7748 1309 7757 1343
rect 7757 1309 7791 1343
rect 7791 1309 7800 1343
rect 7748 1300 7800 1309
rect 8024 1343 8076 1352
rect 8024 1309 8033 1343
rect 8033 1309 8067 1343
rect 8067 1309 8076 1343
rect 8024 1300 8076 1309
rect 10324 1343 10376 1352
rect 10324 1309 10333 1343
rect 10333 1309 10367 1343
rect 10367 1309 10376 1343
rect 10324 1300 10376 1309
rect 10600 1343 10652 1352
rect 10600 1309 10609 1343
rect 10609 1309 10643 1343
rect 10643 1309 10652 1343
rect 10600 1300 10652 1309
rect 11704 1343 11756 1352
rect 11704 1309 11713 1343
rect 11713 1309 11747 1343
rect 11747 1309 11756 1343
rect 11704 1300 11756 1309
rect 14280 1300 14332 1352
rect 15660 1300 15712 1352
rect 15752 1343 15804 1352
rect 15752 1309 15761 1343
rect 15761 1309 15795 1343
rect 15795 1309 15804 1343
rect 15752 1300 15804 1309
rect 17040 1343 17092 1352
rect 17040 1309 17049 1343
rect 17049 1309 17083 1343
rect 17083 1309 17092 1343
rect 17040 1300 17092 1309
rect 17316 1343 17368 1352
rect 17316 1309 17325 1343
rect 17325 1309 17359 1343
rect 17359 1309 17368 1343
rect 17316 1300 17368 1309
rect 22100 1343 22152 1352
rect 22100 1309 22109 1343
rect 22109 1309 22143 1343
rect 22143 1309 22152 1343
rect 22100 1300 22152 1309
rect 2964 1232 3016 1284
rect 13452 1275 13504 1284
rect 13452 1241 13461 1275
rect 13461 1241 13495 1275
rect 13495 1241 13504 1275
rect 13452 1232 13504 1241
rect 18604 1275 18656 1284
rect 18604 1241 18613 1275
rect 18613 1241 18647 1275
rect 18647 1241 18656 1275
rect 18604 1232 18656 1241
rect 23204 1343 23256 1352
rect 23204 1309 23213 1343
rect 23213 1309 23247 1343
rect 23247 1309 23256 1343
rect 23204 1300 23256 1309
rect 24952 1300 25004 1352
rect 25412 1343 25464 1352
rect 25412 1309 25421 1343
rect 25421 1309 25455 1343
rect 25455 1309 25464 1343
rect 25412 1300 25464 1309
rect 26056 1343 26108 1352
rect 26056 1309 26065 1343
rect 26065 1309 26099 1343
rect 26099 1309 26108 1343
rect 26056 1300 26108 1309
rect 26240 1343 26292 1352
rect 26240 1309 26249 1343
rect 26249 1309 26283 1343
rect 26283 1309 26292 1343
rect 26240 1300 26292 1309
rect 27344 1343 27396 1352
rect 27344 1309 27353 1343
rect 27353 1309 27387 1343
rect 27387 1309 27396 1343
rect 27344 1300 27396 1309
rect 27988 1343 28040 1352
rect 27988 1309 27997 1343
rect 27997 1309 28031 1343
rect 28031 1309 28040 1343
rect 27988 1300 28040 1309
rect 28816 1343 28868 1352
rect 28816 1309 28825 1343
rect 28825 1309 28859 1343
rect 28859 1309 28868 1343
rect 28816 1300 28868 1309
rect 30380 1300 30432 1352
rect 31024 1343 31076 1352
rect 31024 1309 31033 1343
rect 31033 1309 31067 1343
rect 31067 1309 31076 1343
rect 31024 1300 31076 1309
rect 32312 1343 32364 1352
rect 32312 1309 32321 1343
rect 32321 1309 32355 1343
rect 32355 1309 32364 1343
rect 32312 1300 32364 1309
rect 35624 1343 35676 1352
rect 35624 1309 35633 1343
rect 35633 1309 35667 1343
rect 35667 1309 35676 1343
rect 35624 1300 35676 1309
rect 36268 1343 36320 1352
rect 36268 1309 36277 1343
rect 36277 1309 36311 1343
rect 36311 1309 36320 1343
rect 36268 1300 36320 1309
rect 36912 1343 36964 1352
rect 36912 1309 36921 1343
rect 36921 1309 36955 1343
rect 36955 1309 36964 1343
rect 36912 1300 36964 1309
rect 38568 1300 38620 1352
rect 38844 1343 38896 1352
rect 38844 1309 38853 1343
rect 38853 1309 38887 1343
rect 38887 1309 38896 1343
rect 38844 1300 38896 1309
rect 39948 1300 40000 1352
rect 40776 1343 40828 1352
rect 40776 1309 40785 1343
rect 40785 1309 40819 1343
rect 40819 1309 40828 1343
rect 40776 1300 40828 1309
rect 41420 1343 41472 1352
rect 41420 1309 41429 1343
rect 41429 1309 41463 1343
rect 41463 1309 41472 1343
rect 41420 1300 41472 1309
rect 42064 1343 42116 1352
rect 42064 1309 42073 1343
rect 42073 1309 42107 1343
rect 42107 1309 42116 1343
rect 42064 1300 42116 1309
rect 43260 1343 43312 1352
rect 43260 1309 43269 1343
rect 43269 1309 43303 1343
rect 43303 1309 43312 1343
rect 43260 1300 43312 1309
rect 43996 1343 44048 1352
rect 43996 1309 44005 1343
rect 44005 1309 44039 1343
rect 44039 1309 44048 1343
rect 43996 1300 44048 1309
rect 44640 1343 44692 1352
rect 44640 1309 44649 1343
rect 44649 1309 44683 1343
rect 44683 1309 44692 1343
rect 44640 1300 44692 1309
rect 45928 1343 45980 1352
rect 45928 1309 45937 1343
rect 45937 1309 45971 1343
rect 45971 1309 45980 1343
rect 45928 1300 45980 1309
rect 46572 1343 46624 1352
rect 46572 1309 46581 1343
rect 46581 1309 46615 1343
rect 46615 1309 46624 1343
rect 46572 1300 46624 1309
rect 47216 1343 47268 1352
rect 47216 1309 47225 1343
rect 47225 1309 47259 1343
rect 47259 1309 47268 1343
rect 47216 1300 47268 1309
rect 48228 1300 48280 1352
rect 49148 1343 49200 1352
rect 49148 1309 49157 1343
rect 49157 1309 49191 1343
rect 49191 1309 49200 1343
rect 49148 1300 49200 1309
rect 49792 1343 49844 1352
rect 49792 1309 49801 1343
rect 49801 1309 49835 1343
rect 49835 1309 49844 1343
rect 49792 1300 49844 1309
rect 50620 1343 50672 1352
rect 50620 1309 50629 1343
rect 50629 1309 50663 1343
rect 50663 1309 50672 1343
rect 50620 1300 50672 1309
rect 51356 1343 51408 1352
rect 51356 1309 51365 1343
rect 51365 1309 51399 1343
rect 51399 1309 51408 1343
rect 51356 1300 51408 1309
rect 52092 1343 52144 1352
rect 52092 1309 52101 1343
rect 52101 1309 52135 1343
rect 52135 1309 52144 1343
rect 52092 1300 52144 1309
rect 53104 1343 53156 1352
rect 53104 1309 53113 1343
rect 53113 1309 53147 1343
rect 53147 1309 53156 1343
rect 53104 1300 53156 1309
rect 54576 1300 54628 1352
rect 54668 1343 54720 1352
rect 54668 1309 54677 1343
rect 54677 1309 54711 1343
rect 54711 1309 54720 1343
rect 54668 1300 54720 1309
rect 55036 1300 55088 1352
rect 56232 1343 56284 1352
rect 56232 1309 56241 1343
rect 56241 1309 56275 1343
rect 56275 1309 56284 1343
rect 56232 1300 56284 1309
rect 56968 1343 57020 1352
rect 56968 1309 56977 1343
rect 56977 1309 57011 1343
rect 57011 1309 57020 1343
rect 56968 1300 57020 1309
rect 58532 1343 58584 1352
rect 58532 1309 58541 1343
rect 58541 1309 58575 1343
rect 58575 1309 58584 1343
rect 58532 1300 58584 1309
rect 59820 1343 59872 1352
rect 59820 1309 59829 1343
rect 59829 1309 59863 1343
rect 59863 1309 59872 1343
rect 59820 1300 59872 1309
rect 60740 1343 60792 1352
rect 60740 1309 60749 1343
rect 60749 1309 60783 1343
rect 60783 1309 60792 1343
rect 60740 1300 60792 1309
rect 62488 1300 62540 1352
rect 63684 1343 63736 1352
rect 63684 1309 63693 1343
rect 63693 1309 63727 1343
rect 63727 1309 63736 1343
rect 63684 1300 63736 1309
rect 64420 1343 64472 1352
rect 64420 1309 64429 1343
rect 64429 1309 64463 1343
rect 64463 1309 64472 1343
rect 64420 1300 64472 1309
rect 66168 1343 66220 1352
rect 66168 1309 66177 1343
rect 66177 1309 66211 1343
rect 66211 1309 66220 1343
rect 66168 1300 66220 1309
rect 69572 1343 69624 1352
rect 69572 1309 69581 1343
rect 69581 1309 69615 1343
rect 69615 1309 69624 1343
rect 69572 1300 69624 1309
rect 43444 1232 43496 1284
rect 2044 1207 2096 1216
rect 2044 1173 2053 1207
rect 2053 1173 2087 1207
rect 2087 1173 2096 1207
rect 2044 1164 2096 1173
rect 13544 1207 13596 1216
rect 13544 1173 13553 1207
rect 13553 1173 13587 1207
rect 13587 1173 13596 1207
rect 13544 1164 13596 1173
rect 18696 1207 18748 1216
rect 18696 1173 18705 1207
rect 18705 1173 18739 1207
rect 18739 1173 18748 1207
rect 18696 1164 18748 1173
rect 21456 1164 21508 1216
rect 28172 1207 28224 1216
rect 28172 1173 28181 1207
rect 28181 1173 28215 1207
rect 28215 1173 28224 1207
rect 28172 1164 28224 1173
rect 29000 1207 29052 1216
rect 29000 1173 29009 1207
rect 29009 1173 29043 1207
rect 29043 1173 29052 1207
rect 29000 1164 29052 1173
rect 30288 1164 30340 1216
rect 31208 1207 31260 1216
rect 31208 1173 31217 1207
rect 31217 1173 31251 1207
rect 31251 1173 31260 1207
rect 31208 1164 31260 1173
rect 32496 1207 32548 1216
rect 32496 1173 32505 1207
rect 32505 1173 32539 1207
rect 32539 1173 32548 1207
rect 32496 1164 32548 1173
rect 35440 1207 35492 1216
rect 35440 1173 35449 1207
rect 35449 1173 35483 1207
rect 35483 1173 35492 1207
rect 35440 1164 35492 1173
rect 36084 1207 36136 1216
rect 36084 1173 36093 1207
rect 36093 1173 36127 1207
rect 36127 1173 36136 1207
rect 36084 1164 36136 1173
rect 36360 1164 36412 1216
rect 37832 1164 37884 1216
rect 38292 1164 38344 1216
rect 39304 1207 39356 1216
rect 39304 1173 39313 1207
rect 39313 1173 39347 1207
rect 39347 1173 39356 1207
rect 39304 1164 39356 1173
rect 40224 1164 40276 1216
rect 41236 1207 41288 1216
rect 41236 1173 41245 1207
rect 41245 1173 41279 1207
rect 41279 1173 41288 1207
rect 41236 1164 41288 1173
rect 41604 1164 41656 1216
rect 42248 1164 42300 1216
rect 43168 1164 43220 1216
rect 47584 1232 47636 1284
rect 70952 1343 71004 1352
rect 70952 1309 70961 1343
rect 70961 1309 70995 1343
rect 70995 1309 71004 1343
rect 70952 1300 71004 1309
rect 72976 1343 73028 1352
rect 72976 1309 72985 1343
rect 72985 1309 73019 1343
rect 73019 1309 73028 1343
rect 72976 1300 73028 1309
rect 74264 1343 74316 1352
rect 74264 1309 74273 1343
rect 74273 1309 74307 1343
rect 74307 1309 74316 1343
rect 74264 1300 74316 1309
rect 89076 1411 89128 1420
rect 89076 1377 89085 1411
rect 89085 1377 89119 1411
rect 89119 1377 89128 1411
rect 89076 1368 89128 1377
rect 74724 1343 74776 1352
rect 74724 1309 74733 1343
rect 74733 1309 74767 1343
rect 74767 1309 74776 1343
rect 74724 1300 74776 1309
rect 75000 1343 75052 1352
rect 75000 1309 75009 1343
rect 75009 1309 75043 1343
rect 75043 1309 75052 1343
rect 75000 1300 75052 1309
rect 77300 1343 77352 1352
rect 77300 1309 77309 1343
rect 77309 1309 77343 1343
rect 77343 1309 77352 1343
rect 77300 1300 77352 1309
rect 77576 1343 77628 1352
rect 77576 1309 77585 1343
rect 77585 1309 77619 1343
rect 77619 1309 77628 1343
rect 77576 1300 77628 1309
rect 79968 1300 80020 1352
rect 80152 1343 80204 1352
rect 80152 1309 80161 1343
rect 80161 1309 80195 1343
rect 80195 1309 80204 1343
rect 80152 1300 80204 1309
rect 82636 1300 82688 1352
rect 82728 1343 82780 1352
rect 82728 1309 82737 1343
rect 82737 1309 82771 1343
rect 82771 1309 82780 1343
rect 82728 1300 82780 1309
rect 85028 1343 85080 1352
rect 85028 1309 85037 1343
rect 85037 1309 85071 1343
rect 85071 1309 85080 1343
rect 85028 1300 85080 1309
rect 85488 1300 85540 1352
rect 86776 1343 86828 1352
rect 86776 1309 86785 1343
rect 86785 1309 86819 1343
rect 86819 1309 86828 1343
rect 86776 1300 86828 1309
rect 45376 1164 45428 1216
rect 45836 1164 45888 1216
rect 47032 1207 47084 1216
rect 47032 1173 47041 1207
rect 47041 1173 47075 1207
rect 47075 1173 47084 1207
rect 47032 1164 47084 1173
rect 47952 1164 48004 1216
rect 49516 1164 49568 1216
rect 50436 1207 50488 1216
rect 50436 1173 50445 1207
rect 50445 1173 50479 1207
rect 50479 1173 50488 1207
rect 50436 1164 50488 1173
rect 51080 1164 51132 1216
rect 51908 1207 51960 1216
rect 51908 1173 51917 1207
rect 51917 1173 51951 1207
rect 51951 1173 51960 1207
rect 51908 1164 51960 1173
rect 52000 1164 52052 1216
rect 55680 1207 55732 1216
rect 55680 1173 55689 1207
rect 55689 1173 55723 1207
rect 55723 1173 55732 1207
rect 55680 1164 55732 1173
rect 56416 1207 56468 1216
rect 56416 1173 56425 1207
rect 56425 1173 56459 1207
rect 56459 1173 56468 1207
rect 56416 1164 56468 1173
rect 57152 1207 57204 1216
rect 57152 1173 57161 1207
rect 57161 1173 57195 1207
rect 57195 1173 57204 1207
rect 57152 1164 57204 1173
rect 60004 1207 60056 1216
rect 60004 1173 60013 1207
rect 60013 1173 60047 1207
rect 60047 1173 60056 1207
rect 60004 1164 60056 1173
rect 60924 1207 60976 1216
rect 60924 1173 60933 1207
rect 60933 1173 60967 1207
rect 60967 1173 60976 1207
rect 60924 1164 60976 1173
rect 63868 1207 63920 1216
rect 63868 1173 63877 1207
rect 63877 1173 63911 1207
rect 63911 1173 63920 1207
rect 63868 1164 63920 1173
rect 64604 1207 64656 1216
rect 64604 1173 64613 1207
rect 64613 1173 64647 1207
rect 64647 1173 64656 1207
rect 64604 1164 64656 1173
rect 65892 1164 65944 1216
rect 72792 1207 72844 1216
rect 72792 1173 72801 1207
rect 72801 1173 72835 1207
rect 72835 1173 72844 1207
rect 72792 1164 72844 1173
rect 74080 1207 74132 1216
rect 74080 1173 74089 1207
rect 74089 1173 74123 1207
rect 74123 1173 74132 1207
rect 74080 1164 74132 1173
rect 84200 1232 84252 1284
rect 88800 1300 88852 1352
rect 89720 1368 89772 1420
rect 90548 1411 90600 1420
rect 90548 1377 90557 1411
rect 90557 1377 90591 1411
rect 90591 1377 90600 1411
rect 90548 1368 90600 1377
rect 94504 1368 94556 1420
rect 94964 1411 95016 1420
rect 94964 1377 94973 1411
rect 94973 1377 95007 1411
rect 95007 1377 95016 1411
rect 94964 1368 95016 1377
rect 95792 1368 95844 1420
rect 97448 1436 97500 1488
rect 99288 1504 99340 1556
rect 105176 1504 105228 1556
rect 107752 1504 107804 1556
rect 107844 1479 107896 1488
rect 107844 1445 107853 1479
rect 107853 1445 107887 1479
rect 107887 1445 107896 1479
rect 107844 1436 107896 1445
rect 109040 1479 109092 1488
rect 109040 1445 109049 1479
rect 109049 1445 109083 1479
rect 109083 1445 109092 1479
rect 109040 1436 109092 1445
rect 111340 1504 111392 1556
rect 117412 1547 117464 1556
rect 117412 1513 117421 1547
rect 117421 1513 117455 1547
rect 117455 1513 117464 1547
rect 117412 1504 117464 1513
rect 118516 1547 118568 1556
rect 118516 1513 118525 1547
rect 118525 1513 118559 1547
rect 118559 1513 118568 1547
rect 118516 1504 118568 1513
rect 120080 1504 120132 1556
rect 126060 1504 126112 1556
rect 129004 1504 129056 1556
rect 115664 1436 115716 1488
rect 117136 1436 117188 1488
rect 120724 1436 120776 1488
rect 123116 1436 123168 1488
rect 133512 1479 133564 1488
rect 133512 1445 133521 1479
rect 133521 1445 133555 1479
rect 133555 1445 133564 1479
rect 133512 1436 133564 1445
rect 138020 1436 138072 1488
rect 138296 1504 138348 1556
rect 141240 1504 141292 1556
rect 142160 1547 142212 1556
rect 142160 1513 142169 1547
rect 142169 1513 142203 1547
rect 142203 1513 142212 1547
rect 142160 1504 142212 1513
rect 143448 1504 143500 1556
rect 140872 1436 140924 1488
rect 141056 1436 141108 1488
rect 145380 1504 145432 1556
rect 146668 1504 146720 1556
rect 90732 1343 90784 1352
rect 90732 1309 90741 1343
rect 90741 1309 90775 1343
rect 90775 1309 90784 1343
rect 90732 1300 90784 1309
rect 90916 1343 90968 1352
rect 90916 1309 90925 1343
rect 90925 1309 90959 1343
rect 90959 1309 90968 1343
rect 90916 1300 90968 1309
rect 91652 1343 91704 1352
rect 91652 1309 91661 1343
rect 91661 1309 91695 1343
rect 91695 1309 91704 1343
rect 91652 1300 91704 1309
rect 80244 1164 80296 1216
rect 87512 1164 87564 1216
rect 88432 1164 88484 1216
rect 92480 1164 92532 1216
rect 92572 1207 92624 1216
rect 92572 1173 92581 1207
rect 92581 1173 92615 1207
rect 92615 1173 92624 1207
rect 92572 1164 92624 1173
rect 93216 1343 93268 1352
rect 93216 1309 93225 1343
rect 93225 1309 93259 1343
rect 93259 1309 93268 1343
rect 93216 1300 93268 1309
rect 93308 1343 93360 1352
rect 93308 1309 93317 1343
rect 93317 1309 93351 1343
rect 93351 1309 93360 1343
rect 93308 1300 93360 1309
rect 93400 1300 93452 1352
rect 93584 1300 93636 1352
rect 94412 1300 94464 1352
rect 95608 1343 95660 1352
rect 95608 1309 95617 1343
rect 95617 1309 95651 1343
rect 95651 1309 95660 1343
rect 95608 1300 95660 1309
rect 96528 1300 96580 1352
rect 98460 1368 98512 1420
rect 98920 1368 98972 1420
rect 97816 1300 97868 1352
rect 97908 1343 97960 1352
rect 97908 1309 97917 1343
rect 97917 1309 97951 1343
rect 97951 1309 97960 1343
rect 97908 1300 97960 1309
rect 98736 1300 98788 1352
rect 99380 1343 99432 1352
rect 99380 1309 99389 1343
rect 99389 1309 99423 1343
rect 99423 1309 99432 1343
rect 99380 1300 99432 1309
rect 100576 1411 100628 1420
rect 100576 1377 100585 1411
rect 100585 1377 100619 1411
rect 100619 1377 100628 1411
rect 100576 1368 100628 1377
rect 99840 1343 99892 1352
rect 99840 1309 99849 1343
rect 99849 1309 99883 1343
rect 99883 1309 99892 1343
rect 99840 1300 99892 1309
rect 100852 1343 100904 1352
rect 100852 1309 100861 1343
rect 100861 1309 100895 1343
rect 100895 1309 100904 1343
rect 100852 1300 100904 1309
rect 101496 1343 101548 1352
rect 101496 1309 101505 1343
rect 101505 1309 101539 1343
rect 101539 1309 101548 1343
rect 101496 1300 101548 1309
rect 101680 1343 101732 1352
rect 101680 1309 101689 1343
rect 101689 1309 101723 1343
rect 101723 1309 101732 1343
rect 101680 1300 101732 1309
rect 106004 1368 106056 1420
rect 109224 1368 109276 1420
rect 110696 1411 110748 1420
rect 110696 1377 110705 1411
rect 110705 1377 110739 1411
rect 110739 1377 110748 1411
rect 110696 1368 110748 1377
rect 103888 1300 103940 1352
rect 104624 1343 104676 1352
rect 104624 1309 104633 1343
rect 104633 1309 104667 1343
rect 104667 1309 104676 1343
rect 104624 1300 104676 1309
rect 105544 1343 105596 1352
rect 105544 1309 105553 1343
rect 105553 1309 105587 1343
rect 105587 1309 105596 1343
rect 105544 1300 105596 1309
rect 105728 1300 105780 1352
rect 106464 1343 106516 1352
rect 106464 1309 106473 1343
rect 106473 1309 106507 1343
rect 106507 1309 106516 1343
rect 106464 1300 106516 1309
rect 107200 1343 107252 1352
rect 107200 1309 107209 1343
rect 107209 1309 107243 1343
rect 107243 1309 107252 1343
rect 107200 1300 107252 1309
rect 107384 1343 107436 1352
rect 107384 1309 107393 1343
rect 107393 1309 107427 1343
rect 107427 1309 107436 1343
rect 107384 1300 107436 1309
rect 108120 1343 108172 1352
rect 108120 1309 108129 1343
rect 108129 1309 108163 1343
rect 108163 1309 108172 1343
rect 108120 1300 108172 1309
rect 108304 1300 108356 1352
rect 109960 1343 110012 1352
rect 109960 1309 109969 1343
rect 109969 1309 110003 1343
rect 110003 1309 110012 1343
rect 109960 1300 110012 1309
rect 110788 1343 110840 1352
rect 111340 1368 111392 1420
rect 111800 1368 111852 1420
rect 110788 1309 110822 1343
rect 110822 1309 110840 1343
rect 110788 1300 110840 1309
rect 111616 1343 111668 1352
rect 111616 1309 111625 1343
rect 111625 1309 111659 1343
rect 111659 1309 111668 1343
rect 111616 1300 111668 1309
rect 94596 1164 94648 1216
rect 97356 1164 97408 1216
rect 99288 1164 99340 1216
rect 100760 1164 100812 1216
rect 108948 1232 109000 1284
rect 112352 1343 112404 1352
rect 112352 1309 112361 1343
rect 112361 1309 112395 1343
rect 112395 1309 112404 1343
rect 112352 1300 112404 1309
rect 113088 1343 113140 1352
rect 113088 1309 113097 1343
rect 113097 1309 113131 1343
rect 113131 1309 113140 1343
rect 113088 1300 113140 1309
rect 113272 1300 113324 1352
rect 114928 1343 114980 1352
rect 114928 1309 114937 1343
rect 114937 1309 114971 1343
rect 114971 1309 114980 1343
rect 114928 1300 114980 1309
rect 115112 1343 115164 1352
rect 115112 1309 115121 1343
rect 115121 1309 115155 1343
rect 115155 1309 115164 1343
rect 115112 1300 115164 1309
rect 115848 1343 115900 1352
rect 115848 1309 115857 1343
rect 115857 1309 115891 1343
rect 115891 1309 115900 1343
rect 115848 1300 115900 1309
rect 116124 1343 116176 1352
rect 116124 1309 116133 1343
rect 116133 1309 116167 1343
rect 116167 1309 116176 1343
rect 116124 1300 116176 1309
rect 126152 1411 126204 1420
rect 126152 1377 126161 1411
rect 126161 1377 126195 1411
rect 126195 1377 126204 1411
rect 126152 1368 126204 1377
rect 128912 1411 128964 1420
rect 128912 1377 128921 1411
rect 128921 1377 128955 1411
rect 128955 1377 128964 1411
rect 128912 1368 128964 1377
rect 132776 1368 132828 1420
rect 140228 1368 140280 1420
rect 117504 1300 117556 1352
rect 118056 1343 118108 1352
rect 118056 1309 118065 1343
rect 118065 1309 118099 1343
rect 118099 1309 118108 1343
rect 118056 1300 118108 1309
rect 118700 1343 118752 1352
rect 118700 1309 118709 1343
rect 118709 1309 118743 1343
rect 118743 1309 118752 1343
rect 118700 1300 118752 1309
rect 119344 1343 119396 1352
rect 119344 1309 119353 1343
rect 119353 1309 119387 1343
rect 119387 1309 119396 1343
rect 119344 1300 119396 1309
rect 120356 1343 120408 1352
rect 120356 1309 120365 1343
rect 120365 1309 120399 1343
rect 120399 1309 120408 1343
rect 120356 1300 120408 1309
rect 121092 1343 121144 1352
rect 121092 1309 121101 1343
rect 121101 1309 121135 1343
rect 121135 1309 121144 1343
rect 121092 1300 121144 1309
rect 121644 1343 121696 1352
rect 121644 1309 121653 1343
rect 121653 1309 121687 1343
rect 121687 1309 121696 1343
rect 121644 1300 121696 1309
rect 122472 1343 122524 1352
rect 122472 1309 122481 1343
rect 122481 1309 122515 1343
rect 122515 1309 122524 1343
rect 122472 1300 122524 1309
rect 123208 1343 123260 1352
rect 123208 1309 123217 1343
rect 123217 1309 123251 1343
rect 123251 1309 123260 1343
rect 123208 1300 123260 1309
rect 125140 1300 125192 1352
rect 125784 1300 125836 1352
rect 126428 1300 126480 1352
rect 127624 1343 127676 1352
rect 127624 1309 127633 1343
rect 127633 1309 127667 1343
rect 127667 1309 127676 1343
rect 127624 1300 127676 1309
rect 129096 1343 129148 1352
rect 129096 1309 129105 1343
rect 129105 1309 129139 1343
rect 129139 1309 129148 1343
rect 129096 1300 129148 1309
rect 130660 1343 130712 1352
rect 130660 1309 130669 1343
rect 130669 1309 130703 1343
rect 130703 1309 130712 1343
rect 130660 1300 130712 1309
rect 132684 1300 132736 1352
rect 133420 1300 133472 1352
rect 134340 1343 134392 1352
rect 134340 1309 134349 1343
rect 134349 1309 134383 1343
rect 134383 1309 134392 1343
rect 134340 1300 134392 1309
rect 138756 1343 138808 1352
rect 138756 1309 138765 1343
rect 138765 1309 138799 1343
rect 138799 1309 138808 1343
rect 138756 1300 138808 1309
rect 138848 1300 138900 1352
rect 140412 1300 140464 1352
rect 141700 1368 141752 1420
rect 141240 1343 141292 1352
rect 141240 1309 141249 1343
rect 141249 1309 141283 1343
rect 141283 1309 141292 1343
rect 141240 1300 141292 1309
rect 141424 1300 141476 1352
rect 143448 1368 143500 1420
rect 146300 1436 146352 1488
rect 146392 1436 146444 1488
rect 148324 1436 148376 1488
rect 151268 1504 151320 1556
rect 151728 1504 151780 1556
rect 153292 1504 153344 1556
rect 156328 1504 156380 1556
rect 156880 1436 156932 1488
rect 144276 1411 144328 1420
rect 144276 1377 144285 1411
rect 144285 1377 144319 1411
rect 144319 1377 144328 1411
rect 144276 1368 144328 1377
rect 143080 1343 143132 1352
rect 143080 1309 143089 1343
rect 143089 1309 143123 1343
rect 143123 1309 143132 1343
rect 143080 1300 143132 1309
rect 103520 1207 103572 1216
rect 103520 1173 103529 1207
rect 103529 1173 103563 1207
rect 103563 1173 103572 1207
rect 103520 1164 103572 1173
rect 103796 1207 103848 1216
rect 103796 1173 103805 1207
rect 103805 1173 103839 1207
rect 103839 1173 103848 1207
rect 103796 1164 103848 1173
rect 107384 1164 107436 1216
rect 110328 1164 110380 1216
rect 117596 1232 117648 1284
rect 118424 1232 118476 1284
rect 112168 1164 112220 1216
rect 114928 1164 114980 1216
rect 117964 1164 118016 1216
rect 118884 1164 118936 1216
rect 121828 1207 121880 1216
rect 121828 1173 121837 1207
rect 121837 1173 121871 1207
rect 121871 1173 121880 1207
rect 121828 1164 121880 1173
rect 122656 1207 122708 1216
rect 122656 1173 122665 1207
rect 122665 1173 122699 1207
rect 122699 1173 122708 1207
rect 122656 1164 122708 1173
rect 123392 1207 123444 1216
rect 123392 1173 123401 1207
rect 123401 1173 123435 1207
rect 123435 1173 123444 1207
rect 123392 1164 123444 1173
rect 124404 1207 124456 1216
rect 124404 1173 124413 1207
rect 124413 1173 124447 1207
rect 124447 1173 124456 1207
rect 124404 1164 124456 1173
rect 125324 1164 125376 1216
rect 127808 1207 127860 1216
rect 127808 1173 127817 1207
rect 127817 1173 127851 1207
rect 127851 1173 127860 1207
rect 127808 1164 127860 1173
rect 130844 1207 130896 1216
rect 130844 1173 130853 1207
rect 130853 1173 130887 1207
rect 130887 1173 130896 1207
rect 130844 1164 130896 1173
rect 132132 1207 132184 1216
rect 132132 1173 132141 1207
rect 132141 1173 132175 1207
rect 132175 1173 132184 1207
rect 132132 1164 132184 1173
rect 134524 1207 134576 1216
rect 134524 1173 134533 1207
rect 134533 1173 134567 1207
rect 134567 1173 134576 1207
rect 134524 1164 134576 1173
rect 138388 1164 138440 1216
rect 139216 1207 139268 1216
rect 139216 1173 139225 1207
rect 139225 1173 139259 1207
rect 139259 1173 139268 1207
rect 139216 1164 139268 1173
rect 144000 1343 144052 1352
rect 144000 1309 144009 1343
rect 144009 1309 144043 1343
rect 144043 1309 144052 1343
rect 144000 1300 144052 1309
rect 144092 1343 144144 1352
rect 144092 1309 144126 1343
rect 144126 1309 144144 1343
rect 144092 1300 144144 1309
rect 144920 1300 144972 1352
rect 145840 1343 145892 1352
rect 145840 1309 145849 1343
rect 145849 1309 145883 1343
rect 145883 1309 145892 1343
rect 145840 1300 145892 1309
rect 146208 1368 146260 1420
rect 148048 1300 148100 1352
rect 144828 1164 144880 1216
rect 149152 1343 149204 1352
rect 149152 1309 149161 1343
rect 149161 1309 149195 1343
rect 149195 1309 149204 1343
rect 149152 1300 149204 1309
rect 149336 1300 149388 1352
rect 150164 1368 150216 1420
rect 150348 1368 150400 1420
rect 150900 1300 150952 1352
rect 150992 1343 151044 1352
rect 150992 1309 151001 1343
rect 151001 1309 151035 1343
rect 151035 1309 151044 1343
rect 150992 1300 151044 1309
rect 151544 1368 151596 1420
rect 154580 1368 154632 1420
rect 176936 1504 176988 1556
rect 177028 1504 177080 1556
rect 211896 1504 211948 1556
rect 216588 1504 216640 1556
rect 219440 1504 219492 1556
rect 219532 1504 219584 1556
rect 220452 1504 220504 1556
rect 223028 1504 223080 1556
rect 223396 1504 223448 1556
rect 157064 1436 157116 1488
rect 178132 1436 178184 1488
rect 196164 1436 196216 1488
rect 198280 1479 198332 1488
rect 198280 1445 198289 1479
rect 198289 1445 198323 1479
rect 198323 1445 198332 1479
rect 198280 1436 198332 1445
rect 203064 1436 203116 1488
rect 209596 1436 209648 1488
rect 210700 1479 210752 1488
rect 210700 1445 210709 1479
rect 210709 1445 210743 1479
rect 210743 1445 210752 1479
rect 210700 1436 210752 1445
rect 152280 1343 152332 1352
rect 152280 1309 152289 1343
rect 152289 1309 152323 1343
rect 152323 1309 152332 1343
rect 152280 1300 152332 1309
rect 153568 1343 153620 1352
rect 153568 1309 153577 1343
rect 153577 1309 153611 1343
rect 153611 1309 153620 1343
rect 153568 1300 153620 1309
rect 154212 1343 154264 1352
rect 154212 1309 154221 1343
rect 154221 1309 154255 1343
rect 154255 1309 154264 1343
rect 154212 1300 154264 1309
rect 154856 1343 154908 1352
rect 154856 1309 154865 1343
rect 154865 1309 154899 1343
rect 154899 1309 154908 1343
rect 154856 1300 154908 1309
rect 156420 1343 156472 1352
rect 156420 1309 156429 1343
rect 156429 1309 156463 1343
rect 156463 1309 156472 1343
rect 156420 1300 156472 1309
rect 157248 1343 157300 1352
rect 157248 1309 157257 1343
rect 157257 1309 157291 1343
rect 157291 1309 157300 1343
rect 157248 1300 157300 1309
rect 158536 1411 158588 1420
rect 158536 1377 158545 1411
rect 158545 1377 158579 1411
rect 158579 1377 158588 1411
rect 158536 1368 158588 1377
rect 159456 1368 159508 1420
rect 162584 1368 162636 1420
rect 159272 1300 159324 1352
rect 161480 1300 161532 1352
rect 163136 1368 163188 1420
rect 166908 1411 166960 1420
rect 166908 1377 166917 1411
rect 166917 1377 166951 1411
rect 166951 1377 166960 1411
rect 166908 1368 166960 1377
rect 167000 1368 167052 1420
rect 169852 1368 169904 1420
rect 171692 1411 171744 1420
rect 171692 1377 171701 1411
rect 171701 1377 171735 1411
rect 171735 1377 171744 1411
rect 171692 1368 171744 1377
rect 191380 1368 191432 1420
rect 196256 1411 196308 1420
rect 196256 1377 196265 1411
rect 196265 1377 196299 1411
rect 196299 1377 196308 1411
rect 196256 1368 196308 1377
rect 197912 1411 197964 1420
rect 197912 1377 197921 1411
rect 197921 1377 197955 1411
rect 197955 1377 197964 1411
rect 197912 1368 197964 1377
rect 201316 1411 201368 1420
rect 201316 1377 201325 1411
rect 201325 1377 201359 1411
rect 201359 1377 201368 1411
rect 201316 1368 201368 1377
rect 205824 1411 205876 1420
rect 205824 1377 205833 1411
rect 205833 1377 205867 1411
rect 205867 1377 205876 1411
rect 205824 1368 205876 1377
rect 210148 1368 210200 1420
rect 213092 1411 213144 1420
rect 213092 1377 213101 1411
rect 213101 1377 213135 1411
rect 213135 1377 213144 1411
rect 213092 1368 213144 1377
rect 217968 1436 218020 1488
rect 220636 1436 220688 1488
rect 220728 1436 220780 1488
rect 229836 1436 229888 1488
rect 213828 1368 213880 1420
rect 215576 1368 215628 1420
rect 218152 1368 218204 1420
rect 218336 1368 218388 1420
rect 222016 1368 222068 1420
rect 224408 1411 224460 1420
rect 224408 1377 224417 1411
rect 224417 1377 224451 1411
rect 224451 1377 224460 1411
rect 224408 1368 224460 1377
rect 227168 1368 227220 1420
rect 227260 1411 227312 1420
rect 227260 1377 227269 1411
rect 227269 1377 227303 1411
rect 227303 1377 227312 1411
rect 227260 1368 227312 1377
rect 162860 1343 162912 1352
rect 162860 1309 162869 1343
rect 162869 1309 162903 1343
rect 162903 1309 162912 1343
rect 162860 1300 162912 1309
rect 164424 1343 164476 1352
rect 164424 1309 164433 1343
rect 164433 1309 164467 1343
rect 164467 1309 164476 1343
rect 164424 1300 164476 1309
rect 167184 1300 167236 1352
rect 168196 1300 168248 1352
rect 172244 1343 172296 1352
rect 172244 1309 172253 1343
rect 172253 1309 172287 1343
rect 172287 1309 172296 1343
rect 172244 1300 172296 1309
rect 172520 1343 172572 1352
rect 172520 1309 172529 1343
rect 172529 1309 172563 1343
rect 172563 1309 172572 1343
rect 172520 1300 172572 1309
rect 173900 1300 173952 1352
rect 174268 1343 174320 1352
rect 174268 1309 174277 1343
rect 174277 1309 174311 1343
rect 174311 1309 174320 1343
rect 174268 1300 174320 1309
rect 175280 1300 175332 1352
rect 176844 1343 176896 1352
rect 176844 1309 176853 1343
rect 176853 1309 176887 1343
rect 176887 1309 176896 1343
rect 176844 1300 176896 1309
rect 178500 1300 178552 1352
rect 179420 1343 179472 1352
rect 179420 1309 179429 1343
rect 179429 1309 179463 1343
rect 179463 1309 179472 1343
rect 179420 1300 179472 1309
rect 180340 1300 180392 1352
rect 181996 1343 182048 1352
rect 181996 1309 182005 1343
rect 182005 1309 182039 1343
rect 182039 1309 182048 1343
rect 181996 1300 182048 1309
rect 183284 1300 183336 1352
rect 184572 1343 184624 1352
rect 184572 1309 184581 1343
rect 184581 1309 184615 1343
rect 184615 1309 184624 1343
rect 184572 1300 184624 1309
rect 185492 1300 185544 1352
rect 187148 1343 187200 1352
rect 187148 1309 187157 1343
rect 187157 1309 187191 1343
rect 187191 1309 187200 1343
rect 187148 1300 187200 1309
rect 188620 1343 188672 1352
rect 188620 1309 188629 1343
rect 188629 1309 188663 1343
rect 188663 1309 188672 1343
rect 188620 1300 188672 1309
rect 189448 1343 189500 1352
rect 189448 1309 189457 1343
rect 189457 1309 189491 1343
rect 189491 1309 189500 1343
rect 189448 1300 189500 1309
rect 189724 1343 189776 1352
rect 189724 1309 189733 1343
rect 189733 1309 189767 1343
rect 189767 1309 189776 1343
rect 189724 1300 189776 1309
rect 191012 1300 191064 1352
rect 191288 1343 191340 1352
rect 191288 1309 191297 1343
rect 191297 1309 191331 1343
rect 191331 1309 191340 1343
rect 191288 1300 191340 1309
rect 150808 1207 150860 1216
rect 150808 1173 150817 1207
rect 150817 1173 150851 1207
rect 150851 1173 150860 1207
rect 150808 1164 150860 1173
rect 152372 1232 152424 1284
rect 154948 1232 155000 1284
rect 155592 1232 155644 1284
rect 157708 1232 157760 1284
rect 194048 1300 194100 1352
rect 194600 1343 194652 1352
rect 194600 1309 194609 1343
rect 194609 1309 194643 1343
rect 194643 1309 194652 1343
rect 194600 1300 194652 1309
rect 196072 1300 196124 1352
rect 196440 1343 196492 1352
rect 196440 1309 196449 1343
rect 196449 1309 196483 1343
rect 196483 1309 196492 1343
rect 196440 1300 196492 1309
rect 198372 1300 198424 1352
rect 200580 1300 200632 1352
rect 201500 1343 201552 1352
rect 201500 1309 201509 1343
rect 201509 1309 201543 1343
rect 201543 1309 201552 1343
rect 201500 1300 201552 1309
rect 206560 1343 206612 1352
rect 206560 1309 206569 1343
rect 206569 1309 206603 1343
rect 206603 1309 206612 1343
rect 206560 1300 206612 1309
rect 207664 1343 207716 1352
rect 207664 1309 207673 1343
rect 207673 1309 207707 1343
rect 207707 1309 207716 1343
rect 207664 1300 207716 1309
rect 208308 1343 208360 1352
rect 208308 1309 208317 1343
rect 208317 1309 208351 1343
rect 208351 1309 208360 1343
rect 208308 1300 208360 1309
rect 208952 1343 209004 1352
rect 208952 1309 208961 1343
rect 208961 1309 208995 1343
rect 208995 1309 209004 1343
rect 208952 1300 209004 1309
rect 210056 1343 210108 1352
rect 210056 1309 210065 1343
rect 210065 1309 210099 1343
rect 210099 1309 210108 1343
rect 210056 1300 210108 1309
rect 210240 1343 210292 1352
rect 210240 1309 210249 1343
rect 210249 1309 210283 1343
rect 210283 1309 210292 1343
rect 210240 1300 210292 1309
rect 210976 1343 211028 1352
rect 210976 1309 210985 1343
rect 210985 1309 211019 1343
rect 211019 1309 211028 1343
rect 210976 1300 211028 1309
rect 211068 1343 211120 1352
rect 211068 1309 211102 1343
rect 211102 1309 211120 1343
rect 211068 1300 211120 1309
rect 212448 1343 212500 1352
rect 212448 1309 212457 1343
rect 212457 1309 212491 1343
rect 212491 1309 212500 1343
rect 212448 1300 212500 1309
rect 212632 1343 212684 1352
rect 212632 1309 212641 1343
rect 212641 1309 212675 1343
rect 212675 1309 212684 1343
rect 212632 1300 212684 1309
rect 213368 1343 213420 1352
rect 213368 1309 213377 1343
rect 213377 1309 213411 1343
rect 213411 1309 213420 1343
rect 213368 1300 213420 1309
rect 213552 1300 213604 1352
rect 215024 1300 215076 1352
rect 193220 1232 193272 1284
rect 201040 1232 201092 1284
rect 153936 1164 153988 1216
rect 154672 1207 154724 1216
rect 154672 1173 154681 1207
rect 154681 1173 154715 1207
rect 154715 1173 154724 1207
rect 154672 1164 154724 1173
rect 160100 1164 160152 1216
rect 161296 1207 161348 1216
rect 161296 1173 161305 1207
rect 161305 1173 161339 1207
rect 161339 1173 161348 1207
rect 161296 1164 161348 1173
rect 162124 1207 162176 1216
rect 162124 1173 162133 1207
rect 162133 1173 162167 1207
rect 162167 1173 162176 1207
rect 162124 1164 162176 1173
rect 163504 1164 163556 1216
rect 164608 1207 164660 1216
rect 164608 1173 164617 1207
rect 164617 1173 164651 1207
rect 164651 1173 164660 1207
rect 164608 1164 164660 1173
rect 167920 1207 167972 1216
rect 167920 1173 167929 1207
rect 167929 1173 167963 1207
rect 167963 1173 167972 1207
rect 167920 1164 167972 1173
rect 169024 1207 169076 1216
rect 169024 1173 169033 1207
rect 169033 1173 169067 1207
rect 169067 1173 169076 1207
rect 169024 1164 169076 1173
rect 187608 1164 187660 1216
rect 192576 1207 192628 1216
rect 192576 1173 192585 1207
rect 192585 1173 192619 1207
rect 192619 1173 192628 1207
rect 192576 1164 192628 1173
rect 192852 1164 192904 1216
rect 193588 1164 193640 1216
rect 195612 1207 195664 1216
rect 195612 1173 195621 1207
rect 195621 1173 195655 1207
rect 195655 1173 195664 1207
rect 195612 1164 195664 1173
rect 199936 1207 199988 1216
rect 199936 1173 199945 1207
rect 199945 1173 199979 1207
rect 199979 1173 199988 1207
rect 199936 1164 199988 1173
rect 202420 1164 202472 1216
rect 207112 1164 207164 1216
rect 208400 1232 208452 1284
rect 209044 1232 209096 1284
rect 207572 1164 207624 1216
rect 209136 1164 209188 1216
rect 209504 1207 209556 1216
rect 209504 1173 209513 1207
rect 209513 1173 209547 1207
rect 209547 1173 209556 1207
rect 209504 1164 209556 1173
rect 212356 1164 212408 1216
rect 214656 1207 214708 1216
rect 214656 1173 214665 1207
rect 214665 1173 214699 1207
rect 214699 1173 214708 1207
rect 214656 1164 214708 1173
rect 216128 1343 216180 1352
rect 216128 1309 216137 1343
rect 216137 1309 216171 1343
rect 216171 1309 216180 1343
rect 216128 1300 216180 1309
rect 216312 1300 216364 1352
rect 216404 1343 216456 1352
rect 216404 1309 216413 1343
rect 216413 1309 216447 1343
rect 216447 1309 216456 1343
rect 216404 1300 216456 1309
rect 217876 1343 217928 1352
rect 217876 1309 217885 1343
rect 217885 1309 217919 1343
rect 217919 1309 217928 1343
rect 217876 1300 217928 1309
rect 217968 1343 218020 1352
rect 217968 1309 217977 1343
rect 217977 1309 218011 1343
rect 218011 1309 218020 1343
rect 217968 1300 218020 1309
rect 218060 1343 218112 1352
rect 218060 1309 218069 1343
rect 218069 1309 218103 1343
rect 218103 1309 218112 1343
rect 218060 1300 218112 1309
rect 218244 1300 218296 1352
rect 219532 1343 219584 1352
rect 219532 1309 219541 1343
rect 219541 1309 219575 1343
rect 219575 1309 219584 1343
rect 219532 1300 219584 1309
rect 220544 1343 220596 1352
rect 220544 1309 220553 1343
rect 220553 1309 220587 1343
rect 220587 1309 220596 1343
rect 220544 1300 220596 1309
rect 221464 1300 221516 1352
rect 221740 1343 221792 1352
rect 221740 1309 221749 1343
rect 221749 1309 221783 1343
rect 221783 1309 221792 1343
rect 221740 1300 221792 1309
rect 217048 1207 217100 1216
rect 217048 1173 217057 1207
rect 217057 1173 217091 1207
rect 217091 1173 217100 1207
rect 217048 1164 217100 1173
rect 218428 1164 218480 1216
rect 218704 1207 218756 1216
rect 218704 1173 218713 1207
rect 218713 1173 218747 1207
rect 218747 1173 218756 1207
rect 218704 1164 218756 1173
rect 220820 1232 220872 1284
rect 223120 1343 223172 1352
rect 223120 1309 223129 1343
rect 223129 1309 223163 1343
rect 223163 1309 223172 1343
rect 223120 1300 223172 1309
rect 223948 1300 224000 1352
rect 225512 1343 225564 1352
rect 225512 1309 225521 1343
rect 225521 1309 225555 1343
rect 225555 1309 225564 1343
rect 225512 1300 225564 1309
rect 226432 1343 226484 1352
rect 226432 1309 226441 1343
rect 226441 1309 226475 1343
rect 226475 1309 226484 1343
rect 226432 1300 226484 1309
rect 227076 1343 227128 1352
rect 227076 1309 227085 1343
rect 227085 1309 227119 1343
rect 227119 1309 227128 1343
rect 227076 1300 227128 1309
rect 228548 1343 228600 1352
rect 228548 1309 228557 1343
rect 228557 1309 228591 1343
rect 228591 1309 228600 1343
rect 228548 1300 228600 1309
rect 230112 1300 230164 1352
rect 230296 1368 230348 1420
rect 243544 1504 243596 1556
rect 246580 1504 246632 1556
rect 253112 1504 253164 1556
rect 269856 1504 269908 1556
rect 231308 1411 231360 1420
rect 231308 1377 231317 1411
rect 231317 1377 231351 1411
rect 231351 1377 231360 1411
rect 231308 1368 231360 1377
rect 235908 1368 235960 1420
rect 239956 1411 240008 1420
rect 239956 1377 239965 1411
rect 239965 1377 239999 1411
rect 239999 1377 240008 1411
rect 239956 1368 240008 1377
rect 231492 1343 231544 1352
rect 231492 1309 231501 1343
rect 231501 1309 231535 1343
rect 231535 1309 231544 1343
rect 231492 1300 231544 1309
rect 233700 1343 233752 1352
rect 233700 1309 233709 1343
rect 233709 1309 233743 1343
rect 233743 1309 233752 1343
rect 233700 1300 233752 1309
rect 235264 1300 235316 1352
rect 236000 1343 236052 1352
rect 236000 1309 236009 1343
rect 236009 1309 236043 1343
rect 236043 1309 236052 1343
rect 236000 1300 236052 1309
rect 240968 1343 241020 1352
rect 240968 1309 240977 1343
rect 240977 1309 241011 1343
rect 241011 1309 241020 1343
rect 240968 1300 241020 1309
rect 241060 1300 241112 1352
rect 241980 1300 242032 1352
rect 243820 1343 243872 1352
rect 243820 1309 243829 1343
rect 243829 1309 243863 1343
rect 243863 1309 243872 1343
rect 243820 1300 243872 1309
rect 246028 1300 246080 1352
rect 225328 1232 225380 1284
rect 222936 1207 222988 1216
rect 222936 1173 222945 1207
rect 222945 1173 222979 1207
rect 222979 1173 222988 1207
rect 222936 1164 222988 1173
rect 224776 1164 224828 1216
rect 226248 1207 226300 1216
rect 226248 1173 226257 1207
rect 226257 1173 226291 1207
rect 226291 1173 226300 1207
rect 226248 1164 226300 1173
rect 226340 1164 226392 1216
rect 244372 1232 244424 1284
rect 244924 1232 244976 1284
rect 247684 1368 247736 1420
rect 250536 1436 250588 1488
rect 268844 1436 268896 1488
rect 257712 1368 257764 1420
rect 246396 1343 246448 1352
rect 246396 1309 246405 1343
rect 246405 1309 246439 1343
rect 246439 1309 246448 1343
rect 246396 1300 246448 1309
rect 247224 1300 247276 1352
rect 247592 1343 247644 1352
rect 247592 1309 247601 1343
rect 247601 1309 247635 1343
rect 247635 1309 247644 1343
rect 247592 1300 247644 1309
rect 246212 1232 246264 1284
rect 228732 1207 228784 1216
rect 228732 1173 228741 1207
rect 228741 1173 228775 1207
rect 228775 1173 228784 1207
rect 228732 1164 228784 1173
rect 229468 1207 229520 1216
rect 229468 1173 229477 1207
rect 229477 1173 229511 1207
rect 229511 1173 229520 1207
rect 229468 1164 229520 1173
rect 231860 1164 231912 1216
rect 233884 1207 233936 1216
rect 233884 1173 233893 1207
rect 233893 1173 233927 1207
rect 233927 1173 233936 1207
rect 233884 1164 233936 1173
rect 234620 1207 234672 1216
rect 234620 1173 234629 1207
rect 234629 1173 234663 1207
rect 234663 1173 234672 1207
rect 234620 1164 234672 1173
rect 235816 1164 235868 1216
rect 246304 1164 246356 1216
rect 248972 1275 249024 1284
rect 248972 1241 248981 1275
rect 248981 1241 249015 1275
rect 249015 1241 249024 1275
rect 248972 1232 249024 1241
rect 248052 1207 248104 1216
rect 248052 1173 248061 1207
rect 248061 1173 248095 1207
rect 248095 1173 248104 1207
rect 248052 1164 248104 1173
rect 248420 1164 248472 1216
rect 251548 1343 251600 1352
rect 251548 1309 251557 1343
rect 251557 1309 251591 1343
rect 251591 1309 251600 1343
rect 251548 1300 251600 1309
rect 252744 1343 252796 1352
rect 252744 1309 252753 1343
rect 252753 1309 252787 1343
rect 252787 1309 252796 1343
rect 252744 1300 252796 1309
rect 252836 1300 252888 1352
rect 254124 1343 254176 1352
rect 254124 1309 254133 1343
rect 254133 1309 254167 1343
rect 254167 1309 254176 1343
rect 254124 1300 254176 1309
rect 255596 1343 255648 1352
rect 255596 1309 255605 1343
rect 255605 1309 255639 1343
rect 255639 1309 255648 1343
rect 255596 1300 255648 1309
rect 255964 1300 256016 1352
rect 256700 1343 256752 1352
rect 256700 1309 256709 1343
rect 256709 1309 256743 1343
rect 256743 1309 256752 1343
rect 256700 1300 256752 1309
rect 256792 1300 256844 1352
rect 257988 1343 258040 1352
rect 257988 1309 257997 1343
rect 257997 1309 258031 1343
rect 258031 1309 258040 1343
rect 257988 1300 258040 1309
rect 258172 1343 258224 1352
rect 258172 1309 258181 1343
rect 258181 1309 258215 1343
rect 258215 1309 258224 1343
rect 258172 1300 258224 1309
rect 258356 1368 258408 1420
rect 261852 1368 261904 1420
rect 271052 1368 271104 1420
rect 259276 1343 259328 1352
rect 259276 1309 259285 1343
rect 259285 1309 259319 1343
rect 259319 1309 259328 1343
rect 259276 1300 259328 1309
rect 255320 1232 255372 1284
rect 255872 1232 255924 1284
rect 260656 1343 260708 1352
rect 260656 1309 260665 1343
rect 260665 1309 260699 1343
rect 260699 1309 260708 1343
rect 260656 1300 260708 1309
rect 251180 1164 251232 1216
rect 258080 1164 258132 1216
rect 258172 1164 258224 1216
rect 261484 1232 261536 1284
rect 263140 1343 263192 1352
rect 263140 1309 263149 1343
rect 263149 1309 263183 1343
rect 263183 1309 263192 1343
rect 263140 1300 263192 1309
rect 264152 1343 264204 1352
rect 264152 1309 264161 1343
rect 264161 1309 264195 1343
rect 264195 1309 264204 1343
rect 264152 1300 264204 1309
rect 264888 1343 264940 1352
rect 264888 1309 264897 1343
rect 264897 1309 264931 1343
rect 264931 1309 264940 1343
rect 264888 1300 264940 1309
rect 265624 1343 265676 1352
rect 265624 1309 265633 1343
rect 265633 1309 265667 1343
rect 265667 1309 265676 1343
rect 265624 1300 265676 1309
rect 266728 1343 266780 1352
rect 266728 1309 266737 1343
rect 266737 1309 266771 1343
rect 266771 1309 266780 1343
rect 266728 1300 266780 1309
rect 267832 1300 267884 1352
rect 268200 1343 268252 1352
rect 268200 1309 268209 1343
rect 268209 1309 268243 1343
rect 268243 1309 268252 1343
rect 268200 1300 268252 1309
rect 269120 1300 269172 1352
rect 270040 1300 270092 1352
rect 270132 1343 270184 1352
rect 270132 1309 270141 1343
rect 270141 1309 270175 1343
rect 270175 1309 270184 1343
rect 270132 1300 270184 1309
rect 261116 1164 261168 1216
rect 262864 1164 262916 1216
rect 264336 1207 264388 1216
rect 264336 1173 264345 1207
rect 264345 1173 264379 1207
rect 264379 1173 264388 1207
rect 264336 1164 264388 1173
rect 264980 1164 265032 1216
rect 265808 1207 265860 1216
rect 265808 1173 265817 1207
rect 265817 1173 265851 1207
rect 265851 1173 265860 1207
rect 265808 1164 265860 1173
rect 266360 1164 266412 1216
rect 267648 1207 267700 1216
rect 267648 1173 267657 1207
rect 267657 1173 267691 1207
rect 267691 1173 267700 1207
rect 267648 1164 267700 1173
rect 268384 1207 268436 1216
rect 268384 1173 268393 1207
rect 268393 1173 268427 1207
rect 268427 1173 268436 1207
rect 268384 1164 268436 1173
rect 270316 1207 270368 1216
rect 270316 1173 270325 1207
rect 270325 1173 270359 1207
rect 270359 1173 270368 1207
rect 270316 1164 270368 1173
rect 68546 1062 68598 1114
rect 68610 1062 68662 1114
rect 68674 1062 68726 1114
rect 68738 1062 68790 1114
rect 68802 1062 68854 1114
rect 136143 1062 136195 1114
rect 136207 1062 136259 1114
rect 136271 1062 136323 1114
rect 136335 1062 136387 1114
rect 136399 1062 136451 1114
rect 203740 1062 203792 1114
rect 203804 1062 203856 1114
rect 203868 1062 203920 1114
rect 203932 1062 203984 1114
rect 203996 1062 204048 1114
rect 271337 1062 271389 1114
rect 271401 1062 271453 1114
rect 271465 1062 271517 1114
rect 271529 1062 271581 1114
rect 271593 1062 271645 1114
rect 2044 960 2096 1012
rect 35992 960 36044 1012
rect 77484 960 77536 1012
rect 103796 960 103848 1012
rect 103980 960 104032 1012
rect 108948 960 109000 1012
rect 17316 892 17368 944
rect 51724 892 51776 944
rect 75000 892 75052 944
rect 99840 892 99892 944
rect 100852 892 100904 944
rect 10600 824 10652 876
rect 44364 824 44416 876
rect 77576 824 77628 876
rect 14280 756 14332 808
rect 45560 756 45612 808
rect 92572 824 92624 876
rect 94780 824 94832 876
rect 97816 824 97868 876
rect 103336 824 103388 876
rect 103520 892 103572 944
rect 104624 892 104676 944
rect 105636 892 105688 944
rect 108304 892 108356 944
rect 110696 960 110748 1012
rect 110788 960 110840 1012
rect 118148 960 118200 1012
rect 109132 892 109184 944
rect 105544 824 105596 876
rect 109684 824 109736 876
rect 113272 892 113324 944
rect 120540 960 120592 1012
rect 141700 960 141752 1012
rect 141792 960 141844 1012
rect 145840 960 145892 1012
rect 147680 960 147732 1012
rect 152280 960 152332 1012
rect 154028 960 154080 1012
rect 179420 960 179472 1012
rect 214932 960 214984 1012
rect 217048 960 217100 1012
rect 218060 960 218112 1012
rect 223120 960 223172 1012
rect 223304 960 223356 1012
rect 226248 960 226300 1012
rect 240048 960 240100 1012
rect 249064 960 249116 1012
rect 250076 960 250128 1012
rect 252836 960 252888 1012
rect 252928 960 252980 1012
rect 138940 892 138992 944
rect 150256 892 150308 944
rect 150440 892 150492 944
rect 154856 892 154908 944
rect 154948 892 155000 944
rect 121460 824 121512 876
rect 95240 756 95292 808
rect 96160 756 96212 808
rect 98736 756 98788 808
rect 98828 756 98880 808
rect 110880 756 110932 808
rect 18696 688 18748 740
rect 51448 688 51500 740
rect 80152 688 80204 740
rect 109960 688 110012 740
rect 110696 688 110748 740
rect 112812 688 112864 740
rect 141700 756 141752 808
rect 148324 824 148376 876
rect 148416 824 148468 876
rect 154212 824 154264 876
rect 214656 892 214708 944
rect 216128 892 216180 944
rect 216680 892 216732 944
rect 219532 892 219584 944
rect 213460 824 213512 876
rect 213552 824 213604 876
rect 246396 892 246448 944
rect 248972 892 249024 944
rect 251732 892 251784 944
rect 260748 960 260800 1012
rect 267924 960 267976 1012
rect 268016 892 268068 944
rect 144000 756 144052 808
rect 150992 756 151044 808
rect 151176 756 151228 808
rect 154672 756 154724 808
rect 162952 756 163004 808
rect 7012 620 7064 672
rect 41328 620 41380 672
rect 72792 620 72844 672
rect 92940 620 92992 672
rect 94872 620 94924 672
rect 107200 620 107252 672
rect 108120 620 108172 672
rect 112628 620 112680 672
rect 113364 620 113416 672
rect 15752 552 15804 604
rect 51632 552 51684 604
rect 82728 552 82780 604
rect 115204 552 115256 604
rect 13544 484 13596 536
rect 47860 484 47912 536
rect 78956 484 79008 536
rect 107384 484 107436 536
rect 144920 620 144972 672
rect 146208 620 146260 672
rect 147680 620 147732 672
rect 147864 688 147916 740
rect 151728 688 151780 740
rect 156420 688 156472 740
rect 160192 688 160244 740
rect 208584 688 208636 740
rect 213644 756 213696 808
rect 218704 756 218756 808
rect 220820 756 220872 808
rect 226432 756 226484 808
rect 228088 756 228140 808
rect 248788 824 248840 876
rect 259276 824 259328 876
rect 215944 688 215996 740
rect 216128 688 216180 740
rect 226892 688 226944 740
rect 243360 688 243412 740
rect 255320 756 255372 808
rect 272064 756 272116 808
rect 152464 620 152516 672
rect 144092 552 144144 604
rect 147588 484 147640 536
rect 2872 416 2924 468
rect 37372 416 37424 468
rect 74080 416 74132 468
rect 97080 416 97132 468
rect 105728 416 105780 468
rect 110972 416 111024 468
rect 146944 416 146996 468
rect 153568 552 153620 604
rect 168380 620 168432 672
rect 243544 620 243596 672
rect 243912 620 243964 672
rect 258264 688 258316 740
rect 249064 620 249116 672
rect 260196 620 260248 672
rect 177028 552 177080 604
rect 208124 552 208176 604
rect 212632 552 212684 604
rect 213460 552 213512 604
rect 216772 552 216824 604
rect 217692 552 217744 604
rect 222936 552 222988 604
rect 223028 552 223080 604
rect 254124 552 254176 604
rect 151636 484 151688 536
rect 153936 484 153988 536
rect 154304 484 154356 536
rect 187148 484 187200 536
rect 209872 484 209924 536
rect 243820 484 243872 536
rect 246856 484 246908 536
rect 256700 484 256752 536
rect 148968 416 149020 468
rect 172428 416 172480 468
rect 208676 416 208728 468
rect 214564 416 214616 468
rect 216312 416 216364 468
rect 251548 416 251600 468
rect 5448 348 5500 400
rect 40040 348 40092 400
rect 92296 348 92348 400
rect 98828 348 98880 400
rect 145012 348 145064 400
rect 150808 348 150860 400
rect 158076 348 158128 400
rect 172520 348 172572 400
rect 214472 348 214524 400
rect 220544 348 220596 400
rect 222384 348 222436 400
rect 241060 348 241112 400
rect 242992 348 243044 400
rect 256424 348 256476 400
rect 147680 280 147732 332
rect 154580 280 154632 332
rect 154764 280 154816 332
rect 184572 280 184624 332
rect 213000 280 213052 332
rect 218244 280 218296 332
rect 218796 280 218848 332
rect 228180 280 228232 332
rect 230572 280 230624 332
rect 248052 280 248104 332
rect 100484 212 100536 264
rect 144736 212 144788 264
rect 155316 212 155368 264
rect 213920 212 213972 264
rect 218612 212 218664 264
rect 223028 212 223080 264
rect 224960 212 225012 264
rect 244832 212 244884 264
rect 209504 144 209556 196
rect 211068 144 211120 196
rect 243728 144 243780 196
rect 28816 76 28868 128
rect 29000 76 29052 128
rect 149336 8 149388 60
rect 181996 8 182048 60
<< metal2 >>
rect 82084 10872 82136 10878
rect 81544 10810 81756 10826
rect 82084 10814 82136 10820
rect 94596 10872 94648 10878
rect 94596 10814 94648 10820
rect 94780 10872 94832 10878
rect 94780 10814 94832 10820
rect 100760 10872 100812 10878
rect 100760 10814 100812 10820
rect 158536 10872 158588 10878
rect 158536 10814 158588 10820
rect 166448 10872 166500 10878
rect 166448 10814 166500 10820
rect 220176 10872 220228 10878
rect 220176 10814 220228 10820
rect 224960 10872 225012 10878
rect 224960 10814 225012 10820
rect 230664 10872 230716 10878
rect 230664 10814 230716 10820
rect 257620 10872 257672 10878
rect 257620 10814 257672 10820
rect 266912 10872 266964 10878
rect 266912 10814 266964 10820
rect 69848 10804 69900 10810
rect 69848 10746 69900 10752
rect 81532 10804 81768 10810
rect 81584 10798 81716 10804
rect 81532 10746 81584 10752
rect 81716 10746 81768 10752
rect 60648 10668 60700 10674
rect 60648 10610 60700 10616
rect 53102 10568 53158 10577
rect 53102 10503 53158 10512
rect 21640 10464 21692 10470
rect 21640 10406 21692 10412
rect 30656 10464 30708 10470
rect 30656 10406 30708 10412
rect 5908 10192 5960 10198
rect 1674 10160 1730 10169
rect 1674 10095 1730 10104
rect 2410 10160 2466 10169
rect 2410 10095 2466 10104
rect 3238 10160 3294 10169
rect 3238 10095 3294 10104
rect 4342 10160 4398 10169
rect 4342 10095 4398 10104
rect 5078 10160 5134 10169
rect 5078 10095 5134 10104
rect 5814 10160 5870 10169
rect 5908 10134 5960 10140
rect 6826 10160 6882 10169
rect 5814 10095 5870 10104
rect 1688 9654 1716 10095
rect 2424 9654 2452 10095
rect 3146 9888 3202 9897
rect 3146 9823 3202 9832
rect 1676 9648 1728 9654
rect 1676 9590 1728 9596
rect 2412 9648 2464 9654
rect 2412 9590 2464 9596
rect 1398 9208 1454 9217
rect 1398 9143 1400 9152
rect 1452 9143 1454 9152
rect 1400 9114 1452 9120
rect 3160 8974 3188 9823
rect 3252 9654 3280 10095
rect 4356 9654 4384 10095
rect 5092 9654 5120 10095
rect 5828 9654 5856 10095
rect 5920 9722 5948 10134
rect 6826 10095 6882 10104
rect 7562 10160 7618 10169
rect 7562 10095 7618 10104
rect 8390 10160 8446 10169
rect 8390 10095 8446 10104
rect 9586 10160 9642 10169
rect 9586 10095 9642 10104
rect 10230 10160 10286 10169
rect 10230 10095 10286 10104
rect 10966 10160 11022 10169
rect 10966 10095 11022 10104
rect 11978 10160 12034 10169
rect 11978 10095 12034 10104
rect 12714 10160 12770 10169
rect 12714 10095 12770 10104
rect 13726 10160 13782 10169
rect 13726 10095 13782 10104
rect 14646 10160 14702 10169
rect 14646 10095 14702 10104
rect 15382 10160 15438 10169
rect 15382 10095 15438 10104
rect 16118 10160 16174 10169
rect 16118 10095 16174 10104
rect 17130 10160 17186 10169
rect 17130 10095 17186 10104
rect 17866 10160 17922 10169
rect 17866 10095 17922 10104
rect 18602 10160 18658 10169
rect 18602 10095 18658 10104
rect 5908 9716 5960 9722
rect 5908 9658 5960 9664
rect 6840 9654 6868 10095
rect 7576 9654 7604 10095
rect 8206 9888 8262 9897
rect 8206 9823 8262 9832
rect 3240 9648 3292 9654
rect 3240 9590 3292 9596
rect 4344 9648 4396 9654
rect 4344 9590 4396 9596
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 7564 9648 7616 9654
rect 7564 9590 7616 9596
rect 7564 9444 7616 9450
rect 7564 9386 7616 9392
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 3252 9178 3280 9318
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3332 8900 3384 8906
rect 3332 8842 3384 8848
rect 3344 4826 3372 8842
rect 4080 7546 4108 9318
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 4448 4214 4476 9318
rect 5184 9042 5212 9318
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 7576 8838 7604 9386
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7668 9110 7696 9318
rect 7656 9104 7708 9110
rect 7656 9046 7708 9052
rect 8220 8974 8248 9823
rect 8404 9654 8432 10095
rect 9600 9654 9628 10095
rect 10244 9654 10272 10095
rect 10980 9654 11008 10095
rect 11992 9654 12020 10095
rect 12728 9654 12756 10095
rect 13450 9888 13506 9897
rect 13450 9823 13506 9832
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 10968 9648 11020 9654
rect 10968 9590 11020 9596
rect 11980 9648 12032 9654
rect 11980 9590 12032 9596
rect 12716 9648 12768 9654
rect 12716 9590 12768 9596
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 12900 9444 12952 9450
rect 12900 9386 12952 9392
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8484 8900 8536 8906
rect 8484 8842 8536 8848
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 8496 6390 8524 8842
rect 9692 8090 9720 9386
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 10336 8634 10364 9318
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 11072 8566 11100 9318
rect 11060 8560 11112 8566
rect 11060 8502 11112 8508
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 12912 6458 12940 9386
rect 13464 8974 13492 9823
rect 13740 9654 13768 10095
rect 14660 9654 14688 10095
rect 15396 9654 15424 10095
rect 16132 9654 16160 10095
rect 17144 9654 17172 10095
rect 17880 9654 17908 10095
rect 18052 9920 18104 9926
rect 18052 9862 18104 9868
rect 18064 9654 18092 9862
rect 18616 9654 18644 10095
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 14648 9648 14700 9654
rect 14648 9590 14700 9596
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 16120 9648 16172 9654
rect 16120 9590 16172 9596
rect 17132 9648 17184 9654
rect 17132 9590 17184 9596
rect 17868 9648 17920 9654
rect 17868 9590 17920 9596
rect 18052 9648 18104 9654
rect 18052 9590 18104 9596
rect 18604 9648 18656 9654
rect 18604 9590 18656 9596
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 17224 9512 17276 9518
rect 17224 9454 17276 9460
rect 13728 9444 13780 9450
rect 13728 9386 13780 9392
rect 15568 9444 15620 9450
rect 15568 9386 15620 9392
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13636 8900 13688 8906
rect 13636 8842 13688 8848
rect 12900 6452 12952 6458
rect 12900 6394 12952 6400
rect 8484 6384 8536 6390
rect 8484 6326 8536 6332
rect 13648 6254 13676 8842
rect 13636 6248 13688 6254
rect 13636 6190 13688 6196
rect 13740 6186 13768 9386
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 14752 8974 14780 9318
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 15580 6322 15608 9386
rect 16500 7954 16528 9454
rect 17236 9042 17264 9454
rect 19156 9444 19208 9450
rect 19156 9386 19208 9392
rect 18604 9376 18656 9382
rect 18604 9318 18656 9324
rect 18696 9376 18748 9382
rect 18696 9318 18748 9324
rect 17224 9036 17276 9042
rect 17224 8978 17276 8984
rect 18420 8968 18472 8974
rect 18420 8910 18472 8916
rect 16488 7948 16540 7954
rect 16488 7890 16540 7896
rect 18432 7818 18460 8910
rect 18616 8362 18644 9318
rect 18604 8356 18656 8362
rect 18604 8298 18656 8304
rect 18420 7812 18472 7818
rect 18420 7754 18472 7760
rect 15568 6316 15620 6322
rect 15568 6258 15620 6264
rect 13728 6180 13780 6186
rect 13728 6122 13780 6128
rect 18708 6118 18736 9318
rect 19168 7750 19196 9386
rect 20260 9376 20312 9382
rect 20260 9318 20312 9324
rect 20272 8974 20300 9318
rect 21652 8974 21680 10406
rect 27712 10396 27764 10402
rect 27712 10338 27764 10344
rect 24492 10328 24544 10334
rect 24492 10270 24544 10276
rect 22652 10124 22704 10130
rect 22652 10066 22704 10072
rect 22468 10056 22520 10062
rect 22468 9998 22520 10004
rect 22480 9586 22508 9998
rect 22468 9580 22520 9586
rect 22468 9522 22520 9528
rect 21732 9036 21784 9042
rect 21732 8978 21784 8984
rect 20260 8968 20312 8974
rect 20260 8910 20312 8916
rect 21088 8968 21140 8974
rect 21088 8910 21140 8916
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21640 8968 21692 8974
rect 21640 8910 21692 8916
rect 21744 8922 21772 8978
rect 22192 8968 22244 8974
rect 22098 8936 22154 8945
rect 19340 8832 19392 8838
rect 19340 8774 19392 8780
rect 19156 7744 19208 7750
rect 19156 7686 19208 7692
rect 19246 6896 19302 6905
rect 19246 6831 19248 6840
rect 19300 6831 19302 6840
rect 19248 6802 19300 6808
rect 18696 6112 18748 6118
rect 18696 6054 18748 6060
rect 19352 5273 19380 8774
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 20720 8560 20772 8566
rect 20720 8502 20772 8508
rect 20732 6662 20760 8502
rect 20824 6730 20852 8570
rect 21100 8362 21128 8910
rect 21362 8664 21418 8673
rect 21468 8634 21496 8910
rect 21744 8894 22098 8922
rect 22192 8910 22244 8916
rect 22098 8871 22154 8880
rect 21640 8832 21692 8838
rect 21640 8774 21692 8780
rect 22100 8832 22152 8838
rect 22100 8774 22152 8780
rect 21362 8599 21364 8608
rect 21416 8599 21418 8608
rect 21456 8628 21508 8634
rect 21364 8570 21416 8576
rect 21456 8570 21508 8576
rect 21088 8356 21140 8362
rect 21088 8298 21140 8304
rect 21652 7886 21680 8774
rect 21914 8392 21970 8401
rect 21914 8327 21970 8336
rect 21928 8022 21956 8327
rect 21916 8016 21968 8022
rect 21916 7958 21968 7964
rect 21640 7880 21692 7886
rect 21640 7822 21692 7828
rect 20812 6724 20864 6730
rect 20812 6666 20864 6672
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 19338 5264 19394 5273
rect 19338 5199 19394 5208
rect 12072 5024 12124 5030
rect 12072 4966 12124 4972
rect 4436 4208 4488 4214
rect 4436 4150 4488 4156
rect 8024 4004 8076 4010
rect 8024 3946 8076 3952
rect 7380 3460 7432 3466
rect 7380 3402 7432 3408
rect 846 2816 902 2825
rect 846 2751 902 2760
rect 860 2650 888 2751
rect 848 2644 900 2650
rect 848 2586 900 2592
rect 1860 2576 1912 2582
rect 1860 2518 1912 2524
rect 4802 2544 4858 2553
rect 1872 2106 1900 2518
rect 4802 2479 4804 2488
rect 4856 2479 4858 2488
rect 5540 2508 5592 2514
rect 4804 2450 4856 2456
rect 5540 2450 5592 2456
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 1860 2100 1912 2106
rect 1860 2042 1912 2048
rect 1676 1964 1728 1970
rect 1676 1906 1728 1912
rect 1688 1057 1716 1906
rect 3792 1896 3844 1902
rect 3792 1838 3844 1844
rect 2872 1352 2924 1358
rect 2872 1294 2924 1300
rect 1952 1284 2004 1290
rect 1952 1226 2004 1232
rect 1674 1048 1730 1057
rect 1674 983 1730 992
rect 1964 649 1992 1226
rect 2044 1216 2096 1222
rect 2044 1158 2096 1164
rect 2056 1018 2084 1158
rect 2044 1012 2096 1018
rect 2044 954 2096 960
rect 1950 640 2006 649
rect 1950 575 2006 584
rect 2884 474 2912 1294
rect 2964 1284 3016 1290
rect 2964 1226 3016 1232
rect 2976 785 3004 1226
rect 3804 1057 3832 1838
rect 4540 1329 4568 2382
rect 5552 1970 5580 2450
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 5540 1964 5592 1970
rect 5540 1906 5592 1912
rect 5172 1896 5224 1902
rect 5172 1838 5224 1844
rect 4526 1320 4582 1329
rect 4526 1255 4582 1264
rect 5184 1057 5212 1838
rect 5356 1352 5408 1358
rect 5356 1294 5408 1300
rect 5448 1352 5500 1358
rect 6748 1329 6776 2382
rect 5448 1294 5500 1300
rect 6734 1320 6790 1329
rect 3790 1048 3846 1057
rect 3790 983 3846 992
rect 5170 1048 5226 1057
rect 5170 983 5226 992
rect 5368 785 5396 1294
rect 2962 776 3018 785
rect 2962 711 3018 720
rect 5354 776 5410 785
rect 5354 711 5410 720
rect 2872 468 2924 474
rect 2872 410 2924 416
rect 5460 406 5488 1294
rect 6734 1255 6790 1264
rect 7024 678 7052 2382
rect 7392 1970 7420 3402
rect 7380 1964 7432 1970
rect 7380 1906 7432 1912
rect 7104 1896 7156 1902
rect 7104 1838 7156 1844
rect 7116 1057 7144 1838
rect 8036 1358 8064 3946
rect 12084 2106 12112 4966
rect 21272 4480 21324 4486
rect 21272 4422 21324 4428
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 12820 2106 12848 4014
rect 15106 3496 15162 3505
rect 15106 3431 15162 3440
rect 14370 3224 14426 3233
rect 14370 3159 14426 3168
rect 12072 2100 12124 2106
rect 12072 2042 12124 2048
rect 12808 2100 12860 2106
rect 12808 2042 12860 2048
rect 8666 2000 8722 2009
rect 14384 1970 14412 3159
rect 15120 2446 15148 3431
rect 14832 2440 14884 2446
rect 14832 2382 14884 2388
rect 15108 2440 15160 2446
rect 15108 2382 15160 2388
rect 8666 1935 8668 1944
rect 8720 1935 8722 1944
rect 11980 1964 12032 1970
rect 8668 1906 8720 1912
rect 11980 1906 12032 1912
rect 12716 1964 12768 1970
rect 12716 1906 12768 1912
rect 14372 1964 14424 1970
rect 14372 1906 14424 1912
rect 8392 1896 8444 1902
rect 8392 1838 8444 1844
rect 9680 1896 9732 1902
rect 9680 1838 9732 1844
rect 7748 1352 7800 1358
rect 7748 1294 7800 1300
rect 8024 1352 8076 1358
rect 8024 1294 8076 1300
rect 7102 1048 7158 1057
rect 7102 983 7158 992
rect 7012 672 7064 678
rect 7012 614 7064 620
rect 7760 513 7788 1294
rect 7746 504 7802 513
rect 7746 439 7802 448
rect 5448 400 5500 406
rect 8404 377 8432 1838
rect 9692 1057 9720 1838
rect 10324 1352 10376 1358
rect 10324 1294 10376 1300
rect 10600 1352 10652 1358
rect 10600 1294 10652 1300
rect 11704 1352 11756 1358
rect 11704 1294 11756 1300
rect 9678 1048 9734 1057
rect 9678 983 9734 992
rect 10336 785 10364 1294
rect 10612 882 10640 1294
rect 10600 876 10652 882
rect 10600 818 10652 824
rect 11716 785 11744 1294
rect 11992 1057 12020 1906
rect 12728 1057 12756 1906
rect 14096 1896 14148 1902
rect 14096 1838 14148 1844
rect 13452 1284 13504 1290
rect 13452 1226 13504 1232
rect 11978 1048 12034 1057
rect 11978 983 12034 992
rect 12714 1048 12770 1057
rect 12714 983 12770 992
rect 10322 776 10378 785
rect 10322 711 10378 720
rect 11702 776 11758 785
rect 11702 711 11758 720
rect 13464 649 13492 1226
rect 13544 1216 13596 1222
rect 13544 1158 13596 1164
rect 13450 640 13506 649
rect 13450 575 13506 584
rect 13556 542 13584 1158
rect 14108 1057 14136 1838
rect 14280 1352 14332 1358
rect 14844 1329 14872 2382
rect 15844 2032 15896 2038
rect 15844 1974 15896 1980
rect 15476 1896 15528 1902
rect 15476 1838 15528 1844
rect 14280 1294 14332 1300
rect 14830 1320 14886 1329
rect 14094 1048 14150 1057
rect 14094 983 14150 992
rect 14292 814 14320 1294
rect 14830 1255 14886 1264
rect 15488 1057 15516 1838
rect 15856 1834 15884 1974
rect 18064 1970 18092 4082
rect 19248 2916 19300 2922
rect 19248 2858 19300 2864
rect 19260 2825 19288 2858
rect 19246 2816 19302 2825
rect 19246 2751 19302 2760
rect 21284 2582 21312 4422
rect 22112 3058 22140 8774
rect 22204 8634 22232 8910
rect 22192 8628 22244 8634
rect 22192 8570 22244 8576
rect 22204 8498 22232 8570
rect 22192 8492 22244 8498
rect 22192 8434 22244 8440
rect 22284 8424 22336 8430
rect 22284 8366 22336 8372
rect 22100 3052 22152 3058
rect 22100 2994 22152 3000
rect 22100 2848 22152 2854
rect 22100 2790 22152 2796
rect 21272 2576 21324 2582
rect 21272 2518 21324 2524
rect 22112 2446 22140 2790
rect 22296 2530 22324 8366
rect 22296 2502 22416 2530
rect 22480 2514 22508 9522
rect 22664 8430 22692 10066
rect 23202 9888 23258 9897
rect 23202 9823 23258 9832
rect 22928 9376 22980 9382
rect 22928 9318 22980 9324
rect 22940 8974 22968 9318
rect 23216 9042 23244 9823
rect 24400 9648 24452 9654
rect 24400 9590 24452 9596
rect 23756 9512 23808 9518
rect 23756 9454 23808 9460
rect 24308 9512 24360 9518
rect 24308 9454 24360 9460
rect 23204 9036 23256 9042
rect 23204 8978 23256 8984
rect 22928 8968 22980 8974
rect 22928 8910 22980 8916
rect 22744 8832 22796 8838
rect 22744 8774 22796 8780
rect 22652 8424 22704 8430
rect 22652 8366 22704 8372
rect 22100 2440 22152 2446
rect 22100 2382 22152 2388
rect 22284 2440 22336 2446
rect 22284 2382 22336 2388
rect 22192 2304 22244 2310
rect 22192 2246 22244 2252
rect 22204 1970 22232 2246
rect 22296 1970 22324 2382
rect 22388 2122 22416 2502
rect 22468 2508 22520 2514
rect 22468 2450 22520 2456
rect 22388 2094 22508 2122
rect 17868 1964 17920 1970
rect 17868 1906 17920 1912
rect 18052 1964 18104 1970
rect 18052 1906 18104 1912
rect 22192 1964 22244 1970
rect 22192 1906 22244 1912
rect 22284 1964 22336 1970
rect 22284 1906 22336 1912
rect 22376 1964 22428 1970
rect 22376 1906 22428 1912
rect 15844 1828 15896 1834
rect 15844 1770 15896 1776
rect 15660 1352 15712 1358
rect 15660 1294 15712 1300
rect 15752 1352 15804 1358
rect 15752 1294 15804 1300
rect 17040 1352 17092 1358
rect 17040 1294 17092 1300
rect 17316 1352 17368 1358
rect 17316 1294 17368 1300
rect 15474 1048 15530 1057
rect 15474 983 15530 992
rect 14280 808 14332 814
rect 15672 785 15700 1294
rect 14280 750 14332 756
rect 15658 776 15714 785
rect 15658 711 15714 720
rect 15764 610 15792 1294
rect 17052 785 17080 1294
rect 17328 950 17356 1294
rect 17880 1057 17908 1906
rect 22008 1760 22060 1766
rect 22006 1728 22008 1737
rect 22100 1760 22152 1766
rect 22060 1728 22062 1737
rect 22100 1702 22152 1708
rect 22006 1663 22062 1672
rect 20718 1592 20774 1601
rect 20718 1527 20720 1536
rect 20772 1527 20774 1536
rect 20720 1498 20772 1504
rect 22112 1358 22140 1702
rect 22388 1465 22416 1906
rect 22480 1902 22508 2094
rect 22468 1896 22520 1902
rect 22520 1844 22600 1850
rect 22468 1838 22600 1844
rect 22480 1822 22600 1838
rect 22572 1766 22600 1822
rect 22560 1760 22612 1766
rect 22560 1702 22612 1708
rect 22374 1456 22430 1465
rect 22664 1426 22692 8366
rect 22756 7886 22784 8774
rect 23388 8560 23440 8566
rect 23388 8502 23440 8508
rect 23112 8424 23164 8430
rect 22926 8392 22982 8401
rect 23112 8366 23164 8372
rect 22926 8327 22982 8336
rect 22940 8022 22968 8327
rect 22928 8016 22980 8022
rect 22928 7958 22980 7964
rect 22744 7880 22796 7886
rect 22744 7822 22796 7828
rect 22834 2816 22890 2825
rect 22834 2751 22890 2760
rect 22848 2650 22876 2751
rect 22836 2644 22888 2650
rect 22836 2586 22888 2592
rect 23124 2145 23152 8366
rect 23204 3528 23256 3534
rect 23204 3470 23256 3476
rect 23110 2136 23166 2145
rect 23110 2071 23166 2080
rect 23124 1902 23152 2071
rect 23112 1896 23164 1902
rect 23112 1838 23164 1844
rect 22374 1391 22430 1400
rect 22652 1420 22704 1426
rect 22652 1362 22704 1368
rect 23216 1358 23244 3470
rect 23296 3052 23348 3058
rect 23296 2994 23348 3000
rect 23308 2446 23336 2994
rect 23400 2514 23428 8502
rect 23662 8392 23718 8401
rect 23480 8356 23532 8362
rect 23662 8327 23718 8336
rect 23480 8298 23532 8304
rect 23492 7886 23520 8298
rect 23676 8022 23704 8327
rect 23664 8016 23716 8022
rect 23664 7958 23716 7964
rect 23480 7880 23532 7886
rect 23480 7822 23532 7828
rect 23572 3392 23624 3398
rect 23572 3334 23624 3340
rect 23480 3188 23532 3194
rect 23480 3130 23532 3136
rect 23492 2582 23520 3130
rect 23480 2576 23532 2582
rect 23480 2518 23532 2524
rect 23388 2508 23440 2514
rect 23388 2450 23440 2456
rect 23296 2440 23348 2446
rect 23296 2382 23348 2388
rect 23308 1970 23336 2382
rect 23296 1964 23348 1970
rect 23296 1906 23348 1912
rect 22100 1352 22152 1358
rect 22100 1294 22152 1300
rect 23204 1352 23256 1358
rect 23584 1329 23612 3334
rect 23664 3052 23716 3058
rect 23664 2994 23716 3000
rect 23676 2650 23704 2994
rect 23664 2644 23716 2650
rect 23664 2586 23716 2592
rect 23768 1465 23796 9454
rect 23938 9208 23994 9217
rect 23938 9143 23940 9152
rect 23992 9143 23994 9152
rect 23940 9114 23992 9120
rect 24032 9104 24084 9110
rect 23952 9052 24032 9058
rect 23952 9046 24084 9052
rect 23952 9030 24072 9046
rect 23952 8906 23980 9030
rect 24032 8968 24084 8974
rect 24032 8910 24084 8916
rect 23940 8900 23992 8906
rect 23940 8842 23992 8848
rect 24044 8634 24072 8910
rect 24032 8628 24084 8634
rect 24032 8570 24084 8576
rect 23848 2848 23900 2854
rect 23848 2790 23900 2796
rect 23754 1456 23810 1465
rect 23754 1391 23756 1400
rect 23808 1391 23810 1400
rect 23756 1362 23808 1368
rect 23860 1329 23888 2790
rect 24320 2582 24348 9454
rect 24412 7478 24440 9590
rect 24504 8430 24532 10270
rect 25504 9988 25556 9994
rect 25504 9930 25556 9936
rect 25516 9518 25544 9930
rect 27620 9920 27672 9926
rect 27620 9862 27672 9868
rect 25870 9752 25926 9761
rect 25870 9687 25872 9696
rect 25924 9687 25926 9696
rect 27342 9752 27398 9761
rect 27342 9687 27344 9696
rect 25872 9658 25924 9664
rect 27396 9687 27398 9696
rect 27344 9658 27396 9664
rect 26148 9648 26200 9654
rect 26148 9590 26200 9596
rect 25688 9580 25740 9586
rect 25688 9522 25740 9528
rect 25504 9512 25556 9518
rect 25504 9454 25556 9460
rect 24584 9444 24636 9450
rect 24584 9386 24636 9392
rect 25228 9444 25280 9450
rect 25228 9386 25280 9392
rect 24492 8424 24544 8430
rect 24492 8366 24544 8372
rect 24400 7472 24452 7478
rect 24400 7414 24452 7420
rect 24504 3058 24532 8366
rect 24596 6798 24624 9386
rect 24676 9376 24728 9382
rect 24676 9318 24728 9324
rect 25136 9376 25188 9382
rect 25136 9318 25188 9324
rect 24688 8974 24716 9318
rect 24676 8968 24728 8974
rect 24676 8910 24728 8916
rect 24768 8832 24820 8838
rect 24768 8774 24820 8780
rect 24780 6866 24808 8774
rect 25044 8288 25096 8294
rect 25044 8230 25096 8236
rect 25056 7886 25084 8230
rect 25044 7880 25096 7886
rect 25044 7822 25096 7828
rect 24952 7540 25004 7546
rect 24952 7482 25004 7488
rect 24768 6860 24820 6866
rect 24768 6802 24820 6808
rect 24584 6792 24636 6798
rect 24584 6734 24636 6740
rect 24964 3126 24992 7482
rect 24952 3120 25004 3126
rect 24952 3062 25004 3068
rect 24492 3052 24544 3058
rect 24492 2994 24544 3000
rect 24584 3052 24636 3058
rect 24584 2994 24636 3000
rect 24400 2848 24452 2854
rect 24400 2790 24452 2796
rect 24308 2576 24360 2582
rect 24308 2518 24360 2524
rect 24412 2446 24440 2790
rect 24596 2446 24624 2994
rect 25042 2816 25098 2825
rect 25042 2751 25098 2760
rect 25056 2650 25084 2751
rect 25044 2644 25096 2650
rect 25044 2586 25096 2592
rect 24768 2576 24820 2582
rect 24768 2518 24820 2524
rect 24400 2440 24452 2446
rect 24400 2382 24452 2388
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 24124 1964 24176 1970
rect 24124 1906 24176 1912
rect 24136 1766 24164 1906
rect 24124 1760 24176 1766
rect 24124 1702 24176 1708
rect 24780 1494 24808 2518
rect 24952 1964 25004 1970
rect 24952 1906 25004 1912
rect 24768 1488 24820 1494
rect 24768 1430 24820 1436
rect 24964 1358 24992 1906
rect 25044 1760 25096 1766
rect 25044 1702 25096 1708
rect 25056 1562 25084 1702
rect 25044 1556 25096 1562
rect 25044 1498 25096 1504
rect 25148 1426 25176 9318
rect 25240 8566 25268 9386
rect 25700 8974 25728 9522
rect 25688 8968 25740 8974
rect 25688 8910 25740 8916
rect 25700 8566 25728 8910
rect 25228 8560 25280 8566
rect 25228 8502 25280 8508
rect 25688 8560 25740 8566
rect 25688 8502 25740 8508
rect 26160 8498 26188 9590
rect 26516 9580 26568 9586
rect 26516 9522 26568 9528
rect 26528 8634 26556 9522
rect 27068 8968 27120 8974
rect 27068 8910 27120 8916
rect 27160 8968 27212 8974
rect 27160 8910 27212 8916
rect 26516 8628 26568 8634
rect 26516 8570 26568 8576
rect 27080 8566 27108 8910
rect 27068 8560 27120 8566
rect 27068 8502 27120 8508
rect 26148 8492 26200 8498
rect 26148 8434 26200 8440
rect 25688 8424 25740 8430
rect 25226 8392 25282 8401
rect 25688 8366 25740 8372
rect 25226 8327 25282 8336
rect 25240 8022 25268 8327
rect 25228 8016 25280 8022
rect 25228 7958 25280 7964
rect 25320 8016 25372 8022
rect 25320 7958 25372 7964
rect 25332 7818 25360 7958
rect 25320 7812 25372 7818
rect 25320 7754 25372 7760
rect 25412 3052 25464 3058
rect 25412 2994 25464 3000
rect 25136 1420 25188 1426
rect 25136 1362 25188 1368
rect 25424 1358 25452 2994
rect 25700 1426 25728 8366
rect 26240 3052 26292 3058
rect 26240 2994 26292 3000
rect 25964 2916 26016 2922
rect 25964 2858 26016 2864
rect 25780 2848 25832 2854
rect 25780 2790 25832 2796
rect 25688 1420 25740 1426
rect 25688 1362 25740 1368
rect 24952 1352 25004 1358
rect 23204 1294 23256 1300
rect 23570 1320 23626 1329
rect 18604 1284 18656 1290
rect 23570 1255 23626 1264
rect 23846 1320 23902 1329
rect 24952 1294 25004 1300
rect 25412 1352 25464 1358
rect 25792 1329 25820 2790
rect 25872 2304 25924 2310
rect 25872 2246 25924 2252
rect 25884 2038 25912 2246
rect 25872 2032 25924 2038
rect 25872 1974 25924 1980
rect 25976 1766 26004 2858
rect 26056 2508 26108 2514
rect 26056 2450 26108 2456
rect 25964 1760 26016 1766
rect 25964 1702 26016 1708
rect 26068 1358 26096 2450
rect 26252 1358 26280 2994
rect 26516 2848 26568 2854
rect 26516 2790 26568 2796
rect 26332 2440 26384 2446
rect 26332 2382 26384 2388
rect 26344 1970 26372 2382
rect 26332 1964 26384 1970
rect 26332 1906 26384 1912
rect 26056 1352 26108 1358
rect 25412 1294 25464 1300
rect 25778 1320 25834 1329
rect 23846 1255 23902 1264
rect 26056 1294 26108 1300
rect 26240 1352 26292 1358
rect 26528 1329 26556 2790
rect 27080 1426 27108 8502
rect 27172 8498 27200 8910
rect 27252 8832 27304 8838
rect 27252 8774 27304 8780
rect 27264 8498 27292 8774
rect 27434 8664 27490 8673
rect 27434 8599 27436 8608
rect 27488 8599 27490 8608
rect 27436 8570 27488 8576
rect 27160 8492 27212 8498
rect 27160 8434 27212 8440
rect 27252 8492 27304 8498
rect 27252 8434 27304 8440
rect 27632 7750 27660 9862
rect 27724 8974 27752 10338
rect 29552 10260 29604 10266
rect 29552 10202 29604 10208
rect 29090 9752 29146 9761
rect 29090 9687 29092 9696
rect 29144 9687 29146 9696
rect 29092 9658 29144 9664
rect 27712 8968 27764 8974
rect 27712 8910 27764 8916
rect 28540 8968 28592 8974
rect 28540 8910 28592 8916
rect 27620 7744 27672 7750
rect 27620 7686 27672 7692
rect 27526 2816 27582 2825
rect 27582 2774 27660 2802
rect 27526 2751 27582 2760
rect 27632 2650 27660 2774
rect 27620 2644 27672 2650
rect 27620 2586 27672 2592
rect 27436 2440 27488 2446
rect 27436 2382 27488 2388
rect 27344 1964 27396 1970
rect 27344 1906 27396 1912
rect 27068 1420 27120 1426
rect 27068 1362 27120 1368
rect 27356 1358 27384 1906
rect 27448 1562 27476 2382
rect 27724 1902 27752 8910
rect 27988 8832 28040 8838
rect 27988 8774 28040 8780
rect 28000 8498 28028 8774
rect 28170 8664 28226 8673
rect 28170 8599 28172 8608
rect 28224 8599 28226 8608
rect 28172 8570 28224 8576
rect 27988 8492 28040 8498
rect 27988 8434 28040 8440
rect 28552 8362 28580 8910
rect 28724 8832 28776 8838
rect 28724 8774 28776 8780
rect 28736 8498 28764 8774
rect 28906 8664 28962 8673
rect 28906 8599 28908 8608
rect 28960 8599 28962 8608
rect 28908 8570 28960 8576
rect 29564 8498 29592 10202
rect 30668 10062 30696 10406
rect 32494 10296 32550 10305
rect 32494 10231 32550 10240
rect 35162 10296 35218 10305
rect 35162 10231 35218 10240
rect 35622 10296 35678 10305
rect 35622 10231 35678 10240
rect 36266 10296 36322 10305
rect 36266 10231 36322 10240
rect 36910 10296 36966 10305
rect 36910 10231 36966 10240
rect 38106 10296 38162 10305
rect 38106 10231 38162 10240
rect 38842 10296 38898 10305
rect 38842 10231 38898 10240
rect 39486 10296 39542 10305
rect 39486 10231 39542 10240
rect 40314 10296 40370 10305
rect 40314 10231 40370 10240
rect 40774 10296 40830 10305
rect 40774 10231 40830 10240
rect 41418 10296 41474 10305
rect 41418 10231 41474 10240
rect 42062 10296 42118 10305
rect 42062 10231 42118 10240
rect 43258 10296 43314 10305
rect 43258 10231 43314 10240
rect 43994 10296 44050 10305
rect 43994 10231 44050 10240
rect 44638 10296 44694 10305
rect 44638 10231 44694 10240
rect 45466 10296 45522 10305
rect 45466 10231 45522 10240
rect 45926 10296 45982 10305
rect 45926 10231 45982 10240
rect 46570 10296 46626 10305
rect 46570 10231 46626 10240
rect 47214 10296 47270 10305
rect 47214 10231 47270 10240
rect 48226 10296 48282 10305
rect 48226 10231 48282 10240
rect 49146 10296 49202 10305
rect 49146 10231 49202 10240
rect 49790 10296 49846 10305
rect 49790 10231 49846 10240
rect 50618 10296 50674 10305
rect 50618 10231 50674 10240
rect 51354 10296 51410 10305
rect 51354 10231 51410 10240
rect 52090 10296 52146 10305
rect 52090 10231 52146 10240
rect 30564 10056 30616 10062
rect 30564 9998 30616 10004
rect 30656 10056 30708 10062
rect 30656 9998 30708 10004
rect 30104 9920 30156 9926
rect 30104 9862 30156 9868
rect 29828 9580 29880 9586
rect 29828 9522 29880 9528
rect 29840 8634 29868 9522
rect 30116 8974 30144 9862
rect 30286 9752 30342 9761
rect 30286 9687 30288 9696
rect 30340 9687 30342 9696
rect 30288 9658 30340 9664
rect 30380 9580 30432 9586
rect 30380 9522 30432 9528
rect 30392 9178 30420 9522
rect 30576 9518 30604 9998
rect 32508 9722 32536 10231
rect 32496 9716 32548 9722
rect 32496 9658 32548 9664
rect 32128 9580 32180 9586
rect 32128 9522 32180 9528
rect 30472 9512 30524 9518
rect 30472 9454 30524 9460
rect 30564 9512 30616 9518
rect 30564 9454 30616 9460
rect 30380 9172 30432 9178
rect 30380 9114 30432 9120
rect 30104 8968 30156 8974
rect 30104 8910 30156 8916
rect 29828 8628 29880 8634
rect 29828 8570 29880 8576
rect 28724 8492 28776 8498
rect 28724 8434 28776 8440
rect 29552 8492 29604 8498
rect 29552 8434 29604 8440
rect 28540 8356 28592 8362
rect 28540 8298 28592 8304
rect 28552 1902 28580 8298
rect 29000 4820 29052 4826
rect 29000 4762 29052 4768
rect 29012 3942 29040 4762
rect 29000 3936 29052 3942
rect 29000 3878 29052 3884
rect 27620 1896 27672 1902
rect 27620 1838 27672 1844
rect 27712 1896 27764 1902
rect 27712 1838 27764 1844
rect 28540 1896 28592 1902
rect 28540 1838 28592 1844
rect 29460 1896 29512 1902
rect 29564 1884 29592 8434
rect 29736 2440 29788 2446
rect 29736 2382 29788 2388
rect 29748 1902 29776 2382
rect 29920 2304 29972 2310
rect 29920 2246 29972 2252
rect 29512 1856 29592 1884
rect 29736 1896 29788 1902
rect 29460 1838 29512 1844
rect 29736 1838 29788 1844
rect 27632 1562 27660 1838
rect 27988 1760 28040 1766
rect 27988 1702 28040 1708
rect 28816 1760 28868 1766
rect 28816 1702 28868 1708
rect 27436 1556 27488 1562
rect 27436 1498 27488 1504
rect 27620 1556 27672 1562
rect 27620 1498 27672 1504
rect 28000 1358 28028 1702
rect 28828 1358 28856 1702
rect 27344 1352 27396 1358
rect 26240 1294 26292 1300
rect 26514 1320 26570 1329
rect 25778 1255 25834 1264
rect 27344 1294 27396 1300
rect 27988 1352 28040 1358
rect 27988 1294 28040 1300
rect 28816 1352 28868 1358
rect 28816 1294 28868 1300
rect 26514 1255 26570 1264
rect 18604 1226 18656 1232
rect 17866 1048 17922 1057
rect 17866 983 17922 992
rect 17316 944 17368 950
rect 17316 886 17368 892
rect 17038 776 17094 785
rect 17038 711 17094 720
rect 15752 604 15804 610
rect 15752 546 15804 552
rect 13544 536 13596 542
rect 13544 478 13596 484
rect 18616 377 18644 1226
rect 18696 1216 18748 1222
rect 18696 1158 18748 1164
rect 21456 1216 21508 1222
rect 21456 1158 21508 1164
rect 28172 1216 28224 1222
rect 28172 1158 28224 1164
rect 29000 1216 29052 1222
rect 29932 1193 29960 2246
rect 30116 1902 30144 8910
rect 30484 6866 30512 9454
rect 32140 9178 32168 9522
rect 34748 9276 35056 9285
rect 34748 9274 34754 9276
rect 34810 9274 34834 9276
rect 34890 9274 34914 9276
rect 34970 9274 34994 9276
rect 35050 9274 35056 9276
rect 34810 9222 34812 9274
rect 34992 9222 34994 9274
rect 34748 9220 34754 9222
rect 34810 9220 34834 9222
rect 34890 9220 34914 9222
rect 34970 9220 34994 9222
rect 35050 9220 35056 9222
rect 33046 9208 33102 9217
rect 34748 9211 35056 9220
rect 32128 9172 32180 9178
rect 35176 9178 35204 10231
rect 35636 9586 35664 10231
rect 36280 9586 36308 10231
rect 36924 9586 36952 10231
rect 38120 9586 38148 10231
rect 38200 9716 38252 9722
rect 38200 9658 38252 9664
rect 35624 9580 35676 9586
rect 35624 9522 35676 9528
rect 36268 9580 36320 9586
rect 36268 9522 36320 9528
rect 36912 9580 36964 9586
rect 36912 9522 36964 9528
rect 38108 9580 38160 9586
rect 38108 9522 38160 9528
rect 35624 9376 35676 9382
rect 35624 9318 35676 9324
rect 35808 9376 35860 9382
rect 35808 9318 35860 9324
rect 36636 9376 36688 9382
rect 36636 9318 36688 9324
rect 37924 9376 37976 9382
rect 37924 9318 37976 9324
rect 33046 9143 33048 9152
rect 32128 9114 32180 9120
rect 33100 9143 33102 9152
rect 35164 9172 35216 9178
rect 33048 9114 33100 9120
rect 35164 9114 35216 9120
rect 31852 9036 31904 9042
rect 31852 8978 31904 8984
rect 32772 9036 32824 9042
rect 32772 8978 32824 8984
rect 32956 9036 33008 9042
rect 32956 8978 33008 8984
rect 30748 8968 30800 8974
rect 30748 8910 30800 8916
rect 30472 6860 30524 6866
rect 30472 6802 30524 6808
rect 30760 1902 30788 8910
rect 30840 8832 30892 8838
rect 30840 8774 30892 8780
rect 30852 8498 30880 8774
rect 31022 8664 31078 8673
rect 31022 8599 31024 8608
rect 31076 8599 31078 8608
rect 31024 8570 31076 8576
rect 30840 8492 30892 8498
rect 30840 8434 30892 8440
rect 31864 1902 31892 8978
rect 31944 8968 31996 8974
rect 31944 8910 31996 8916
rect 31956 8430 31984 8910
rect 32784 8838 32812 8978
rect 32772 8832 32824 8838
rect 32772 8774 32824 8780
rect 32864 8492 32916 8498
rect 32864 8434 32916 8440
rect 31944 8424 31996 8430
rect 31944 8366 31996 8372
rect 32876 7954 32904 8434
rect 32968 8362 32996 8978
rect 33140 8968 33192 8974
rect 33140 8910 33192 8916
rect 33152 8634 33180 8910
rect 33140 8628 33192 8634
rect 33140 8570 33192 8576
rect 33692 8492 33744 8498
rect 33692 8434 33744 8440
rect 32956 8356 33008 8362
rect 32956 8298 33008 8304
rect 32864 7948 32916 7954
rect 32864 7890 32916 7896
rect 33704 7206 33732 8434
rect 34748 8188 35056 8197
rect 34748 8186 34754 8188
rect 34810 8186 34834 8188
rect 34890 8186 34914 8188
rect 34970 8186 34994 8188
rect 35050 8186 35056 8188
rect 34810 8134 34812 8186
rect 34992 8134 34994 8186
rect 34748 8132 34754 8134
rect 34810 8132 34834 8134
rect 34890 8132 34914 8134
rect 34970 8132 34994 8134
rect 35050 8132 35056 8134
rect 34748 8123 35056 8132
rect 33968 7880 34020 7886
rect 33968 7822 34020 7828
rect 33980 7750 34008 7822
rect 33968 7744 34020 7750
rect 33968 7686 34020 7692
rect 33692 7200 33744 7206
rect 33692 7142 33744 7148
rect 34748 7100 35056 7109
rect 34748 7098 34754 7100
rect 34810 7098 34834 7100
rect 34890 7098 34914 7100
rect 34970 7098 34994 7100
rect 35050 7098 35056 7100
rect 34810 7046 34812 7098
rect 34992 7046 34994 7098
rect 34748 7044 34754 7046
rect 34810 7044 34834 7046
rect 34890 7044 34914 7046
rect 34970 7044 34994 7046
rect 35050 7044 35056 7046
rect 34748 7035 35056 7044
rect 34748 6012 35056 6021
rect 34748 6010 34754 6012
rect 34810 6010 34834 6012
rect 34890 6010 34914 6012
rect 34970 6010 34994 6012
rect 35050 6010 35056 6012
rect 34810 5958 34812 6010
rect 34992 5958 34994 6010
rect 34748 5956 34754 5958
rect 34810 5956 34834 5958
rect 34890 5956 34914 5958
rect 34970 5956 34994 5958
rect 35050 5956 35056 5958
rect 34748 5947 35056 5956
rect 35532 5636 35584 5642
rect 35532 5578 35584 5584
rect 35544 5030 35572 5578
rect 35532 5024 35584 5030
rect 35532 4966 35584 4972
rect 34748 4924 35056 4933
rect 34748 4922 34754 4924
rect 34810 4922 34834 4924
rect 34890 4922 34914 4924
rect 34970 4922 34994 4924
rect 35050 4922 35056 4924
rect 34810 4870 34812 4922
rect 34992 4870 34994 4922
rect 34748 4868 34754 4870
rect 34810 4868 34834 4870
rect 34890 4868 34914 4870
rect 34970 4868 34994 4870
rect 35050 4868 35056 4870
rect 34748 4859 35056 4868
rect 35636 4622 35664 9318
rect 35820 5302 35848 9318
rect 36452 8900 36504 8906
rect 36452 8842 36504 8848
rect 36084 5364 36136 5370
rect 36084 5306 36136 5312
rect 35808 5296 35860 5302
rect 35808 5238 35860 5244
rect 35900 5228 35952 5234
rect 35900 5170 35952 5176
rect 35992 5228 36044 5234
rect 35992 5170 36044 5176
rect 35624 4616 35676 4622
rect 35624 4558 35676 4564
rect 35912 4554 35940 5170
rect 35900 4548 35952 4554
rect 35900 4490 35952 4496
rect 35440 4480 35492 4486
rect 35440 4422 35492 4428
rect 34748 3836 35056 3845
rect 34748 3834 34754 3836
rect 34810 3834 34834 3836
rect 34890 3834 34914 3836
rect 34970 3834 34994 3836
rect 35050 3834 35056 3836
rect 34810 3782 34812 3834
rect 34992 3782 34994 3834
rect 34748 3780 34754 3782
rect 34810 3780 34834 3782
rect 34890 3780 34914 3782
rect 34970 3780 34994 3782
rect 35050 3780 35056 3782
rect 34748 3771 35056 3780
rect 32770 3088 32826 3097
rect 32770 3023 32826 3032
rect 31944 2984 31996 2990
rect 31944 2926 31996 2932
rect 31956 2446 31984 2926
rect 32784 2446 32812 3023
rect 34748 2748 35056 2757
rect 34748 2746 34754 2748
rect 34810 2746 34834 2748
rect 34890 2746 34914 2748
rect 34970 2746 34994 2748
rect 35050 2746 35056 2748
rect 34810 2694 34812 2746
rect 34992 2694 34994 2746
rect 34748 2692 34754 2694
rect 34810 2692 34834 2694
rect 34890 2692 34914 2694
rect 34970 2692 34994 2694
rect 35050 2692 35056 2694
rect 34748 2683 35056 2692
rect 31944 2440 31996 2446
rect 31944 2382 31996 2388
rect 32772 2440 32824 2446
rect 32772 2382 32824 2388
rect 32496 2372 32548 2378
rect 32496 2314 32548 2320
rect 32508 1970 32536 2314
rect 32680 2304 32732 2310
rect 32680 2246 32732 2252
rect 32692 1970 32720 2246
rect 32496 1964 32548 1970
rect 32496 1906 32548 1912
rect 32680 1964 32732 1970
rect 32680 1906 32732 1912
rect 30104 1896 30156 1902
rect 30104 1838 30156 1844
rect 30748 1896 30800 1902
rect 30748 1838 30800 1844
rect 31300 1896 31352 1902
rect 31300 1838 31352 1844
rect 31852 1896 31904 1902
rect 31852 1838 31904 1844
rect 30380 1760 30432 1766
rect 30380 1702 30432 1708
rect 31024 1760 31076 1766
rect 31024 1702 31076 1708
rect 30392 1358 30420 1702
rect 31036 1358 31064 1702
rect 31312 1494 31340 1838
rect 32312 1760 32364 1766
rect 32312 1702 32364 1708
rect 33140 1760 33192 1766
rect 33140 1702 33192 1708
rect 35164 1760 35216 1766
rect 35164 1702 35216 1708
rect 31300 1488 31352 1494
rect 31300 1430 31352 1436
rect 32324 1358 32352 1702
rect 33152 1601 33180 1702
rect 34748 1660 35056 1669
rect 34748 1658 34754 1660
rect 34810 1658 34834 1660
rect 34890 1658 34914 1660
rect 34970 1658 34994 1660
rect 35050 1658 35056 1660
rect 34810 1606 34812 1658
rect 34992 1606 34994 1658
rect 34748 1604 34754 1606
rect 34810 1604 34834 1606
rect 34890 1604 34914 1606
rect 34970 1604 34994 1606
rect 35050 1604 35056 1606
rect 33138 1592 33194 1601
rect 34748 1595 35056 1604
rect 33138 1527 33194 1536
rect 30380 1352 30432 1358
rect 30380 1294 30432 1300
rect 31024 1352 31076 1358
rect 31024 1294 31076 1300
rect 32312 1352 32364 1358
rect 32312 1294 32364 1300
rect 30288 1216 30340 1222
rect 29000 1158 29052 1164
rect 29918 1184 29974 1193
rect 18708 746 18736 1158
rect 18696 740 18748 746
rect 18696 682 18748 688
rect 21468 649 21496 1158
rect 28184 649 28212 1158
rect 21454 640 21510 649
rect 21454 575 21510 584
rect 28170 640 28226 649
rect 28170 575 28226 584
rect 5448 342 5500 348
rect 8390 368 8446 377
rect 8390 303 8446 312
rect 18602 368 18658 377
rect 18602 303 18658 312
rect 28814 368 28870 377
rect 28814 303 28870 312
rect 28828 134 28856 303
rect 29012 134 29040 1158
rect 30288 1158 30340 1164
rect 31208 1216 31260 1222
rect 31208 1158 31260 1164
rect 32496 1216 32548 1222
rect 32496 1158 32548 1164
rect 29918 1119 29974 1128
rect 30300 649 30328 1158
rect 31220 649 31248 1158
rect 32508 649 32536 1158
rect 35176 649 35204 1702
rect 35452 1222 35480 4422
rect 35624 1352 35676 1358
rect 35624 1294 35676 1300
rect 35440 1216 35492 1222
rect 35440 1158 35492 1164
rect 35636 649 35664 1294
rect 36004 1018 36032 5170
rect 36096 1222 36124 5306
rect 36268 5296 36320 5302
rect 36266 5264 36268 5273
rect 36320 5264 36322 5273
rect 36266 5199 36322 5208
rect 36464 4554 36492 8842
rect 36452 4548 36504 4554
rect 36452 4490 36504 4496
rect 36544 4548 36596 4554
rect 36544 4490 36596 4496
rect 36556 4010 36584 4490
rect 36544 4004 36596 4010
rect 36544 3946 36596 3952
rect 36648 3534 36676 9318
rect 37004 5364 37056 5370
rect 37004 5306 37056 5312
rect 36728 5228 36780 5234
rect 36728 5170 36780 5176
rect 36740 4146 36768 5170
rect 36820 5024 36872 5030
rect 36818 4992 36820 5001
rect 36912 5024 36964 5030
rect 36872 4992 36874 5001
rect 36912 4966 36964 4972
rect 36818 4927 36874 4936
rect 36820 4684 36872 4690
rect 36820 4626 36872 4632
rect 36728 4140 36780 4146
rect 36728 4082 36780 4088
rect 36832 4010 36860 4626
rect 36924 4078 36952 4966
rect 37016 4826 37044 5306
rect 37096 5160 37148 5166
rect 37096 5102 37148 5108
rect 37004 4820 37056 4826
rect 37004 4762 37056 4768
rect 37108 4690 37136 5102
rect 37096 4684 37148 4690
rect 37096 4626 37148 4632
rect 37280 4616 37332 4622
rect 37280 4558 37332 4564
rect 36912 4072 36964 4078
rect 36912 4014 36964 4020
rect 36820 4004 36872 4010
rect 36820 3946 36872 3952
rect 36728 3936 36780 3942
rect 36728 3878 36780 3884
rect 36636 3528 36688 3534
rect 36740 3516 36768 3878
rect 37292 3534 37320 4558
rect 37832 4208 37884 4214
rect 37832 4150 37884 4156
rect 37372 4004 37424 4010
rect 37372 3946 37424 3952
rect 37384 3602 37412 3946
rect 37372 3596 37424 3602
rect 37372 3538 37424 3544
rect 36820 3528 36872 3534
rect 36740 3488 36820 3516
rect 36636 3470 36688 3476
rect 36820 3470 36872 3476
rect 37280 3528 37332 3534
rect 37280 3470 37332 3476
rect 36360 3392 36412 3398
rect 36360 3334 36412 3340
rect 37372 3392 37424 3398
rect 37372 3334 37424 3340
rect 36268 1352 36320 1358
rect 36268 1294 36320 1300
rect 36084 1216 36136 1222
rect 36084 1158 36136 1164
rect 35992 1012 36044 1018
rect 35992 954 36044 960
rect 36280 649 36308 1294
rect 36372 1222 36400 3334
rect 36912 1352 36964 1358
rect 36912 1294 36964 1300
rect 36360 1216 36412 1222
rect 36360 1158 36412 1164
rect 36924 649 36952 1294
rect 30286 640 30342 649
rect 30286 575 30342 584
rect 31206 640 31262 649
rect 31206 575 31262 584
rect 32494 640 32550 649
rect 32494 575 32550 584
rect 35162 640 35218 649
rect 35162 575 35218 584
rect 35622 640 35678 649
rect 35622 575 35678 584
rect 36266 640 36322 649
rect 36266 575 36322 584
rect 36910 640 36966 649
rect 36910 575 36966 584
rect 37384 474 37412 3334
rect 37648 3120 37700 3126
rect 37648 3062 37700 3068
rect 37660 2106 37688 3062
rect 37648 2100 37700 2106
rect 37648 2042 37700 2048
rect 37844 1222 37872 4150
rect 37936 3126 37964 9318
rect 38016 4616 38068 4622
rect 38016 4558 38068 4564
rect 38028 4146 38056 4558
rect 38016 4140 38068 4146
rect 38016 4082 38068 4088
rect 38028 3126 38056 4082
rect 37924 3120 37976 3126
rect 37924 3062 37976 3068
rect 38016 3120 38068 3126
rect 38016 3062 38068 3068
rect 38028 2378 38056 3062
rect 38212 2446 38240 9658
rect 38856 9586 38884 10231
rect 39500 9586 39528 10231
rect 39580 10192 39632 10198
rect 39580 10134 39632 10140
rect 38844 9580 38896 9586
rect 38844 9522 38896 9528
rect 39488 9580 39540 9586
rect 39488 9522 39540 9528
rect 38660 9376 38712 9382
rect 38660 9318 38712 9324
rect 38384 4276 38436 4282
rect 38384 4218 38436 4224
rect 38396 4146 38424 4218
rect 38672 4214 38700 9318
rect 39396 8832 39448 8838
rect 39396 8774 39448 8780
rect 39212 8084 39264 8090
rect 39212 8026 39264 8032
rect 38844 6792 38896 6798
rect 38844 6734 38896 6740
rect 39120 6792 39172 6798
rect 39120 6734 39172 6740
rect 38752 6384 38804 6390
rect 38752 6326 38804 6332
rect 38764 5098 38792 6326
rect 38752 5092 38804 5098
rect 38752 5034 38804 5040
rect 38660 4208 38712 4214
rect 38660 4150 38712 4156
rect 38752 4208 38804 4214
rect 38752 4150 38804 4156
rect 38384 4140 38436 4146
rect 38384 4082 38436 4088
rect 38476 4072 38528 4078
rect 38476 4014 38528 4020
rect 38488 3602 38516 4014
rect 38476 3596 38528 3602
rect 38476 3538 38528 3544
rect 38488 2990 38516 3538
rect 38568 3052 38620 3058
rect 38568 2994 38620 3000
rect 38476 2984 38528 2990
rect 38476 2926 38528 2932
rect 38488 2514 38516 2926
rect 38476 2508 38528 2514
rect 38476 2450 38528 2456
rect 38200 2440 38252 2446
rect 38200 2382 38252 2388
rect 38016 2372 38068 2378
rect 38016 2314 38068 2320
rect 38476 2372 38528 2378
rect 38476 2314 38528 2320
rect 38292 2304 38344 2310
rect 38292 2246 38344 2252
rect 38384 2304 38436 2310
rect 38384 2246 38436 2252
rect 38108 1964 38160 1970
rect 38108 1906 38160 1912
rect 37832 1216 37884 1222
rect 37832 1158 37884 1164
rect 38120 649 38148 1906
rect 38304 1222 38332 2246
rect 38396 1834 38424 2246
rect 38488 2106 38516 2314
rect 38476 2100 38528 2106
rect 38476 2042 38528 2048
rect 38580 2038 38608 2994
rect 38764 2553 38792 4150
rect 38856 2774 38884 6734
rect 38934 4040 38990 4049
rect 38934 3975 38936 3984
rect 38988 3975 38990 3984
rect 39028 4004 39080 4010
rect 38936 3946 38988 3952
rect 39028 3946 39080 3952
rect 38856 2746 38976 2774
rect 38750 2544 38806 2553
rect 38750 2479 38806 2488
rect 38948 2446 38976 2746
rect 38936 2440 38988 2446
rect 38936 2382 38988 2388
rect 39040 2038 39068 3946
rect 39132 3194 39160 6734
rect 39120 3188 39172 3194
rect 39120 3130 39172 3136
rect 39224 3126 39252 8026
rect 39212 3120 39264 3126
rect 39212 3062 39264 3068
rect 39408 2038 39436 8774
rect 39488 3392 39540 3398
rect 39488 3334 39540 3340
rect 39500 3194 39528 3334
rect 39488 3188 39540 3194
rect 39488 3130 39540 3136
rect 39592 2038 39620 10134
rect 39672 9716 39724 9722
rect 39672 9658 39724 9664
rect 39684 8906 39712 9658
rect 40328 8974 40356 10231
rect 40788 9586 40816 10231
rect 41432 9586 41460 10231
rect 42076 9586 42104 10231
rect 43272 9586 43300 10231
rect 44008 9586 44036 10231
rect 44652 9586 44680 10231
rect 40776 9580 40828 9586
rect 40776 9522 40828 9528
rect 41420 9580 41472 9586
rect 41420 9522 41472 9528
rect 42064 9580 42116 9586
rect 42064 9522 42116 9528
rect 43260 9580 43312 9586
rect 43260 9522 43312 9528
rect 43996 9580 44048 9586
rect 43996 9522 44048 9528
rect 44640 9580 44692 9586
rect 44640 9522 44692 9528
rect 40500 9376 40552 9382
rect 40500 9318 40552 9324
rect 41052 9376 41104 9382
rect 41052 9318 41104 9324
rect 41788 9376 41840 9382
rect 41788 9318 41840 9324
rect 42892 9376 42944 9382
rect 42892 9318 42944 9324
rect 43260 9376 43312 9382
rect 43260 9318 43312 9324
rect 43904 9376 43956 9382
rect 43904 9318 43956 9324
rect 40316 8968 40368 8974
rect 40316 8910 40368 8916
rect 39672 8900 39724 8906
rect 39672 8842 39724 8848
rect 40512 2446 40540 9318
rect 40868 6860 40920 6866
rect 40868 6802 40920 6808
rect 40592 2984 40644 2990
rect 40592 2926 40644 2932
rect 40132 2440 40184 2446
rect 40132 2382 40184 2388
rect 40500 2440 40552 2446
rect 40500 2382 40552 2388
rect 39856 2304 39908 2310
rect 39856 2246 39908 2252
rect 38568 2032 38620 2038
rect 38568 1974 38620 1980
rect 39028 2032 39080 2038
rect 39028 1974 39080 1980
rect 39304 2032 39356 2038
rect 39304 1974 39356 1980
rect 39396 2032 39448 2038
rect 39396 1974 39448 1980
rect 39580 2032 39632 2038
rect 39580 1974 39632 1980
rect 38384 1828 38436 1834
rect 38384 1770 38436 1776
rect 38568 1352 38620 1358
rect 38568 1294 38620 1300
rect 38844 1352 38896 1358
rect 38844 1294 38896 1300
rect 38292 1216 38344 1222
rect 38292 1158 38344 1164
rect 38580 649 38608 1294
rect 38106 640 38162 649
rect 38106 575 38162 584
rect 38566 640 38622 649
rect 38566 575 38622 584
rect 37372 468 37424 474
rect 37372 410 37424 416
rect 38856 377 38884 1294
rect 39316 1222 39344 1974
rect 39304 1216 39356 1222
rect 39304 1158 39356 1164
rect 39868 513 39896 2246
rect 40040 2032 40092 2038
rect 40040 1974 40092 1980
rect 39948 1352 40000 1358
rect 39948 1294 40000 1300
rect 39960 649 39988 1294
rect 39946 640 40002 649
rect 39946 575 40002 584
rect 39854 504 39910 513
rect 39854 439 39910 448
rect 40052 406 40080 1974
rect 40144 1902 40172 2382
rect 40604 2378 40632 2926
rect 40880 2774 40908 6802
rect 40960 5092 41012 5098
rect 40960 5034 41012 5040
rect 40972 4826 41000 5034
rect 40960 4820 41012 4826
rect 40960 4762 41012 4768
rect 41064 3534 41092 9318
rect 41512 9104 41564 9110
rect 41512 9046 41564 9052
rect 41144 3936 41196 3942
rect 41144 3878 41196 3884
rect 41156 3534 41184 3878
rect 41052 3528 41104 3534
rect 41052 3470 41104 3476
rect 41144 3528 41196 3534
rect 41144 3470 41196 3476
rect 41156 2990 41184 3470
rect 41524 3466 41552 9046
rect 41800 4622 41828 9318
rect 42708 6452 42760 6458
rect 42708 6394 42760 6400
rect 42614 5128 42670 5137
rect 42248 5092 42300 5098
rect 42614 5063 42670 5072
rect 42248 5034 42300 5040
rect 42260 4622 42288 5034
rect 42628 5030 42656 5063
rect 42616 5024 42668 5030
rect 42616 4966 42668 4972
rect 42720 4690 42748 6394
rect 42798 5944 42854 5953
rect 42798 5879 42854 5888
rect 42812 4826 42840 5879
rect 42800 4820 42852 4826
rect 42800 4762 42852 4768
rect 42524 4684 42576 4690
rect 42524 4626 42576 4632
rect 42708 4684 42760 4690
rect 42708 4626 42760 4632
rect 41788 4616 41840 4622
rect 41788 4558 41840 4564
rect 42248 4616 42300 4622
rect 42248 4558 42300 4564
rect 41880 4548 41932 4554
rect 41880 4490 41932 4496
rect 41604 4480 41656 4486
rect 41604 4422 41656 4428
rect 41512 3460 41564 3466
rect 41512 3402 41564 3408
rect 41236 3392 41288 3398
rect 41236 3334 41288 3340
rect 41328 3392 41380 3398
rect 41328 3334 41380 3340
rect 41144 2984 41196 2990
rect 41144 2926 41196 2932
rect 40880 2746 41000 2774
rect 40972 2446 41000 2746
rect 40960 2440 41012 2446
rect 40960 2382 41012 2388
rect 41052 2440 41104 2446
rect 41052 2382 41104 2388
rect 40592 2372 40644 2378
rect 40592 2314 40644 2320
rect 40224 2304 40276 2310
rect 40224 2246 40276 2252
rect 40132 1896 40184 1902
rect 40132 1838 40184 1844
rect 40236 1222 40264 2246
rect 40604 2106 40632 2314
rect 40592 2100 40644 2106
rect 40592 2042 40644 2048
rect 41064 1902 41092 2382
rect 41052 1896 41104 1902
rect 41052 1838 41104 1844
rect 40408 1760 40460 1766
rect 40406 1728 40408 1737
rect 40460 1728 40462 1737
rect 40406 1663 40462 1672
rect 40776 1352 40828 1358
rect 40776 1294 40828 1300
rect 40224 1216 40276 1222
rect 40224 1158 40276 1164
rect 40788 649 40816 1294
rect 41248 1222 41276 3334
rect 41340 2514 41368 3334
rect 41328 2508 41380 2514
rect 41328 2450 41380 2456
rect 41328 2304 41380 2310
rect 41328 2246 41380 2252
rect 41512 2304 41564 2310
rect 41512 2246 41564 2252
rect 41236 1216 41288 1222
rect 41236 1158 41288 1164
rect 41340 678 41368 2246
rect 41524 2106 41552 2246
rect 41512 2100 41564 2106
rect 41512 2042 41564 2048
rect 41420 1352 41472 1358
rect 41420 1294 41472 1300
rect 41328 672 41380 678
rect 40774 640 40830 649
rect 41432 649 41460 1294
rect 41616 1222 41644 4422
rect 41892 4282 41920 4490
rect 41880 4276 41932 4282
rect 41880 4218 41932 4224
rect 41892 3942 41920 4218
rect 42536 4078 42564 4626
rect 42614 4176 42670 4185
rect 42614 4111 42616 4120
rect 42668 4111 42670 4120
rect 42616 4082 42668 4088
rect 42524 4072 42576 4078
rect 42524 4014 42576 4020
rect 41880 3936 41932 3942
rect 41880 3878 41932 3884
rect 42432 3936 42484 3942
rect 42432 3878 42484 3884
rect 42064 3392 42116 3398
rect 42064 3334 42116 3340
rect 42076 2961 42104 3334
rect 42444 3194 42472 3878
rect 42536 3602 42564 4014
rect 42524 3596 42576 3602
rect 42524 3538 42576 3544
rect 42432 3188 42484 3194
rect 42432 3130 42484 3136
rect 42062 2952 42118 2961
rect 42062 2887 42118 2896
rect 42904 2446 42932 9318
rect 42984 7472 43036 7478
rect 42984 7414 43036 7420
rect 42996 2446 43024 7414
rect 43272 3126 43300 9318
rect 43534 4584 43590 4593
rect 43534 4519 43590 4528
rect 43352 4140 43404 4146
rect 43352 4082 43404 4088
rect 43364 3466 43392 4082
rect 43352 3460 43404 3466
rect 43352 3402 43404 3408
rect 43364 3126 43392 3402
rect 43444 3392 43496 3398
rect 43444 3334 43496 3340
rect 43168 3120 43220 3126
rect 43168 3062 43220 3068
rect 43260 3120 43312 3126
rect 43260 3062 43312 3068
rect 43352 3120 43404 3126
rect 43352 3062 43404 3068
rect 42892 2440 42944 2446
rect 42892 2382 42944 2388
rect 42984 2440 43036 2446
rect 42984 2382 43036 2388
rect 42248 2304 42300 2310
rect 42248 2246 42300 2252
rect 42064 1352 42116 1358
rect 42064 1294 42116 1300
rect 41604 1216 41656 1222
rect 41604 1158 41656 1164
rect 42076 649 42104 1294
rect 42260 1222 42288 2246
rect 43180 1222 43208 3062
rect 43364 2446 43392 3062
rect 43352 2440 43404 2446
rect 43352 2382 43404 2388
rect 43352 2304 43404 2310
rect 43352 2246 43404 2252
rect 43364 2009 43392 2246
rect 43350 2000 43406 2009
rect 43350 1935 43406 1944
rect 43260 1352 43312 1358
rect 43260 1294 43312 1300
rect 42248 1216 42300 1222
rect 42248 1158 42300 1164
rect 43168 1216 43220 1222
rect 43168 1158 43220 1164
rect 43272 649 43300 1294
rect 43456 1290 43484 3334
rect 43548 2650 43576 4519
rect 43916 3534 43944 9318
rect 45480 8974 45508 10231
rect 45940 9586 45968 10231
rect 46584 9586 46612 10231
rect 47228 9586 47256 10231
rect 48240 9586 48268 10231
rect 49160 9586 49188 10231
rect 49804 9586 49832 10231
rect 50632 9586 50660 10231
rect 51368 9586 51396 10231
rect 52104 9586 52132 10231
rect 53116 9586 53144 10503
rect 58532 10328 58584 10334
rect 53286 10296 53342 10305
rect 53286 10231 53342 10240
rect 53838 10296 53894 10305
rect 53838 10231 53894 10240
rect 54850 10296 54906 10305
rect 54850 10231 54906 10240
rect 55678 10296 55734 10305
rect 55678 10231 55734 10240
rect 56506 10296 56562 10305
rect 56506 10231 56562 10240
rect 57334 10296 57390 10305
rect 57334 10231 57390 10240
rect 57794 10296 57850 10305
rect 58532 10270 58584 10276
rect 58806 10296 58862 10305
rect 57794 10231 57850 10240
rect 45928 9580 45980 9586
rect 45928 9522 45980 9528
rect 46572 9580 46624 9586
rect 46572 9522 46624 9528
rect 47216 9580 47268 9586
rect 47216 9522 47268 9528
rect 48228 9580 48280 9586
rect 48228 9522 48280 9528
rect 49148 9580 49200 9586
rect 49148 9522 49200 9528
rect 49792 9580 49844 9586
rect 49792 9522 49844 9528
rect 50620 9580 50672 9586
rect 50620 9522 50672 9528
rect 51356 9580 51408 9586
rect 51356 9522 51408 9528
rect 52092 9580 52144 9586
rect 52092 9522 52144 9528
rect 53104 9580 53156 9586
rect 53104 9522 53156 9528
rect 46204 9444 46256 9450
rect 46204 9386 46256 9392
rect 48596 9444 48648 9450
rect 48596 9386 48648 9392
rect 51816 9444 51868 9450
rect 51816 9386 51868 9392
rect 45652 9376 45704 9382
rect 45652 9318 45704 9324
rect 46020 9376 46072 9382
rect 46020 9318 46072 9324
rect 45468 8968 45520 8974
rect 45468 8910 45520 8916
rect 44732 8832 44784 8838
rect 44732 8774 44784 8780
rect 43996 6724 44048 6730
rect 43996 6666 44048 6672
rect 44008 3534 44036 6666
rect 44088 5228 44140 5234
rect 44088 5170 44140 5176
rect 44100 4826 44128 5170
rect 44088 4820 44140 4826
rect 44088 4762 44140 4768
rect 44364 4616 44416 4622
rect 44364 4558 44416 4564
rect 44376 4214 44404 4558
rect 44456 4480 44508 4486
rect 44456 4422 44508 4428
rect 44468 4214 44496 4422
rect 44364 4208 44416 4214
rect 44364 4150 44416 4156
rect 44456 4208 44508 4214
rect 44456 4150 44508 4156
rect 44744 4146 44772 8774
rect 45100 6656 45152 6662
rect 45100 6598 45152 6604
rect 45112 4146 45140 6598
rect 45664 5710 45692 9318
rect 45652 5704 45704 5710
rect 45652 5646 45704 5652
rect 45744 5636 45796 5642
rect 45744 5578 45796 5584
rect 45376 5568 45428 5574
rect 45376 5510 45428 5516
rect 45284 4480 45336 4486
rect 45284 4422 45336 4428
rect 44732 4140 44784 4146
rect 44732 4082 44784 4088
rect 45100 4140 45152 4146
rect 45100 4082 45152 4088
rect 44088 4004 44140 4010
rect 44088 3946 44140 3952
rect 43904 3528 43956 3534
rect 43904 3470 43956 3476
rect 43996 3528 44048 3534
rect 43996 3470 44048 3476
rect 43812 3460 43864 3466
rect 43812 3402 43864 3408
rect 43824 2990 43852 3402
rect 44100 3194 44128 3946
rect 44456 3936 44508 3942
rect 44456 3878 44508 3884
rect 44468 3738 44496 3878
rect 44456 3732 44508 3738
rect 44456 3674 44508 3680
rect 44364 3392 44416 3398
rect 44364 3334 44416 3340
rect 44088 3188 44140 3194
rect 44088 3130 44140 3136
rect 43812 2984 43864 2990
rect 43812 2926 43864 2932
rect 44100 2938 44128 3130
rect 43824 2774 43852 2926
rect 44100 2922 44220 2938
rect 44100 2916 44232 2922
rect 44100 2910 44180 2916
rect 44180 2858 44232 2864
rect 43824 2746 44036 2774
rect 43536 2644 43588 2650
rect 43536 2586 43588 2592
rect 44008 2514 44036 2746
rect 43996 2508 44048 2514
rect 43996 2450 44048 2456
rect 43996 1352 44048 1358
rect 43996 1294 44048 1300
rect 43444 1284 43496 1290
rect 43444 1226 43496 1232
rect 44008 649 44036 1294
rect 44376 882 44404 3334
rect 45296 1834 45324 4422
rect 45284 1828 45336 1834
rect 45284 1770 45336 1776
rect 44640 1352 44692 1358
rect 44640 1294 44692 1300
rect 44364 876 44416 882
rect 44364 818 44416 824
rect 44652 649 44680 1294
rect 45388 1222 45416 5510
rect 45468 4752 45520 4758
rect 45468 4694 45520 4700
rect 45480 4078 45508 4694
rect 45756 4554 45784 5578
rect 46032 5302 46060 9318
rect 46216 9110 46244 9386
rect 47032 9376 47084 9382
rect 47032 9318 47084 9324
rect 48228 9376 48280 9382
rect 48228 9318 48280 9324
rect 48412 9376 48464 9382
rect 48412 9318 48464 9324
rect 46204 9104 46256 9110
rect 46204 9046 46256 9052
rect 46112 7948 46164 7954
rect 46112 7890 46164 7896
rect 46124 5710 46152 7890
rect 46664 6724 46716 6730
rect 46664 6666 46716 6672
rect 46676 5914 46704 6666
rect 46664 5908 46716 5914
rect 46664 5850 46716 5856
rect 46480 5772 46532 5778
rect 46480 5714 46532 5720
rect 46112 5704 46164 5710
rect 46112 5646 46164 5652
rect 45836 5296 45888 5302
rect 45836 5238 45888 5244
rect 46020 5296 46072 5302
rect 46020 5238 46072 5244
rect 45744 4548 45796 4554
rect 45744 4490 45796 4496
rect 45756 4282 45784 4490
rect 45744 4276 45796 4282
rect 45744 4218 45796 4224
rect 45560 4208 45612 4214
rect 45560 4150 45612 4156
rect 45468 4072 45520 4078
rect 45468 4014 45520 4020
rect 45480 3602 45508 4014
rect 45468 3596 45520 3602
rect 45468 3538 45520 3544
rect 45468 1964 45520 1970
rect 45468 1906 45520 1912
rect 45376 1216 45428 1222
rect 45376 1158 45428 1164
rect 45480 649 45508 1906
rect 45572 814 45600 4150
rect 45744 3936 45796 3942
rect 45744 3878 45796 3884
rect 45560 808 45612 814
rect 45756 785 45784 3878
rect 45848 1222 45876 5238
rect 46204 5228 46256 5234
rect 46204 5170 46256 5176
rect 46216 4554 46244 5170
rect 46492 5166 46520 5714
rect 46940 5704 46992 5710
rect 46940 5646 46992 5652
rect 46664 5296 46716 5302
rect 46664 5238 46716 5244
rect 46572 5228 46624 5234
rect 46572 5170 46624 5176
rect 46480 5160 46532 5166
rect 46400 5108 46480 5114
rect 46400 5102 46532 5108
rect 46400 5086 46520 5102
rect 46400 4758 46428 5086
rect 46584 4808 46612 5170
rect 46676 5137 46704 5238
rect 46756 5228 46808 5234
rect 46756 5170 46808 5176
rect 46662 5128 46718 5137
rect 46662 5063 46718 5072
rect 46768 4826 46796 5170
rect 46492 4780 46612 4808
rect 46756 4820 46808 4826
rect 46388 4752 46440 4758
rect 46388 4694 46440 4700
rect 46492 4690 46520 4780
rect 46756 4762 46808 4768
rect 46480 4684 46532 4690
rect 46480 4626 46532 4632
rect 46952 4622 46980 5646
rect 47044 4622 47072 9318
rect 47492 6248 47544 6254
rect 47492 6190 47544 6196
rect 47216 5636 47268 5642
rect 47216 5578 47268 5584
rect 47122 5128 47178 5137
rect 47122 5063 47124 5072
rect 47176 5063 47178 5072
rect 47124 5034 47176 5040
rect 46940 4616 46992 4622
rect 46940 4558 46992 4564
rect 47032 4616 47084 4622
rect 47032 4558 47084 4564
rect 46204 4548 46256 4554
rect 46204 4490 46256 4496
rect 47032 4480 47084 4486
rect 47032 4422 47084 4428
rect 45928 1352 45980 1358
rect 45928 1294 45980 1300
rect 46572 1352 46624 1358
rect 46572 1294 46624 1300
rect 45836 1216 45888 1222
rect 45836 1158 45888 1164
rect 45560 750 45612 756
rect 45742 776 45798 785
rect 45742 711 45798 720
rect 45940 649 45968 1294
rect 46584 649 46612 1294
rect 47044 1222 47072 4422
rect 47122 4176 47178 4185
rect 47228 4162 47256 5578
rect 47504 4622 47532 6190
rect 48044 6180 48096 6186
rect 48044 6122 48096 6128
rect 47952 5704 48004 5710
rect 47952 5646 48004 5652
rect 47492 4616 47544 4622
rect 47492 4558 47544 4564
rect 47964 4486 47992 5646
rect 48056 4826 48084 6122
rect 48044 4820 48096 4826
rect 48044 4762 48096 4768
rect 48136 4820 48188 4826
rect 48136 4762 48188 4768
rect 47860 4480 47912 4486
rect 47860 4422 47912 4428
rect 47952 4480 48004 4486
rect 47952 4422 48004 4428
rect 47178 4134 47256 4162
rect 47122 4111 47178 4120
rect 47136 4078 47164 4111
rect 47124 4072 47176 4078
rect 47124 4014 47176 4020
rect 47676 3936 47728 3942
rect 47676 3878 47728 3884
rect 47582 3360 47638 3369
rect 47582 3295 47638 3304
rect 47492 3188 47544 3194
rect 47492 3130 47544 3136
rect 47504 2650 47532 3130
rect 47492 2644 47544 2650
rect 47492 2586 47544 2592
rect 47216 1352 47268 1358
rect 47216 1294 47268 1300
rect 47032 1216 47084 1222
rect 47032 1158 47084 1164
rect 47228 649 47256 1294
rect 47596 1290 47624 3295
rect 47688 2990 47716 3878
rect 47768 3596 47820 3602
rect 47768 3538 47820 3544
rect 47780 2990 47808 3538
rect 47676 2984 47728 2990
rect 47676 2926 47728 2932
rect 47768 2984 47820 2990
rect 47768 2926 47820 2932
rect 47584 1284 47636 1290
rect 47584 1226 47636 1232
rect 41328 614 41380 620
rect 41418 640 41474 649
rect 40774 575 40830 584
rect 41418 575 41474 584
rect 42062 640 42118 649
rect 42062 575 42118 584
rect 43258 640 43314 649
rect 43258 575 43314 584
rect 43994 640 44050 649
rect 43994 575 44050 584
rect 44638 640 44694 649
rect 44638 575 44694 584
rect 45466 640 45522 649
rect 45466 575 45522 584
rect 45926 640 45982 649
rect 45926 575 45982 584
rect 46570 640 46626 649
rect 46570 575 46626 584
rect 47214 640 47270 649
rect 47214 575 47270 584
rect 47872 542 47900 4422
rect 47952 4072 48004 4078
rect 47952 4014 48004 4020
rect 47964 3602 47992 4014
rect 48148 3738 48176 4762
rect 48136 3732 48188 3738
rect 48136 3674 48188 3680
rect 47952 3596 48004 3602
rect 48240 3584 48268 9318
rect 48320 5568 48372 5574
rect 48320 5510 48372 5516
rect 48332 4554 48360 5510
rect 48320 4548 48372 4554
rect 48320 4490 48372 4496
rect 48424 4434 48452 9318
rect 48504 4548 48556 4554
rect 48504 4490 48556 4496
rect 47952 3538 48004 3544
rect 48148 3556 48268 3584
rect 48332 4406 48452 4434
rect 48148 3176 48176 3556
rect 48332 3482 48360 4406
rect 48412 4276 48464 4282
rect 48412 4218 48464 4224
rect 48424 3942 48452 4218
rect 48412 3936 48464 3942
rect 48412 3878 48464 3884
rect 48332 3466 48452 3482
rect 48228 3460 48280 3466
rect 48332 3460 48464 3466
rect 48332 3454 48412 3460
rect 48228 3402 48280 3408
rect 48412 3402 48464 3408
rect 48240 3369 48268 3402
rect 48226 3360 48282 3369
rect 48226 3295 48282 3304
rect 48056 3148 48176 3176
rect 47952 3120 48004 3126
rect 47952 3062 48004 3068
rect 47964 1222 47992 3062
rect 48056 3058 48084 3148
rect 48516 3058 48544 4490
rect 48608 4146 48636 9386
rect 50436 9376 50488 9382
rect 50436 9318 50488 9324
rect 51264 9376 51316 9382
rect 51264 9318 51316 9324
rect 48964 8016 49016 8022
rect 48964 7958 49016 7964
rect 48872 6248 48924 6254
rect 48872 6190 48924 6196
rect 48688 4480 48740 4486
rect 48688 4422 48740 4428
rect 48596 4140 48648 4146
rect 48596 4082 48648 4088
rect 48700 3482 48728 4422
rect 48778 3632 48834 3641
rect 48778 3567 48834 3576
rect 48792 3534 48820 3567
rect 48608 3466 48728 3482
rect 48780 3528 48832 3534
rect 48780 3470 48832 3476
rect 48596 3460 48728 3466
rect 48648 3454 48728 3460
rect 48596 3402 48648 3408
rect 48884 3380 48912 6190
rect 48976 3534 49004 7958
rect 49516 6316 49568 6322
rect 49516 6258 49568 6264
rect 49056 4480 49108 4486
rect 49056 4422 49108 4428
rect 49068 4146 49096 4422
rect 49528 4214 49556 6258
rect 49792 4548 49844 4554
rect 49792 4490 49844 4496
rect 49804 4282 49832 4490
rect 49792 4276 49844 4282
rect 49792 4218 49844 4224
rect 49148 4208 49200 4214
rect 49516 4208 49568 4214
rect 49200 4168 49464 4196
rect 49148 4150 49200 4156
rect 49056 4140 49108 4146
rect 49056 4082 49108 4088
rect 48964 3528 49016 3534
rect 48964 3470 49016 3476
rect 49330 3496 49386 3505
rect 49330 3431 49386 3440
rect 49344 3398 49372 3431
rect 48700 3352 48912 3380
rect 49332 3392 49384 3398
rect 48700 3058 48728 3352
rect 49332 3334 49384 3340
rect 49054 3224 49110 3233
rect 49054 3159 49110 3168
rect 49068 3126 49096 3159
rect 49056 3120 49108 3126
rect 49108 3068 49188 3074
rect 49056 3062 49188 3068
rect 49068 3058 49188 3062
rect 48044 3052 48096 3058
rect 48044 2994 48096 3000
rect 48504 3052 48556 3058
rect 48504 2994 48556 3000
rect 48688 3052 48740 3058
rect 49068 3052 49200 3058
rect 49068 3046 49148 3052
rect 48688 2994 48740 3000
rect 49148 2994 49200 3000
rect 49238 2952 49294 2961
rect 49238 2887 49240 2896
rect 49292 2887 49294 2896
rect 49240 2858 49292 2864
rect 49436 2774 49464 4168
rect 49516 4150 49568 4156
rect 50448 3534 50476 9318
rect 51172 8288 51224 8294
rect 51172 8230 51224 8236
rect 50988 5296 51040 5302
rect 50988 5238 51040 5244
rect 50896 4752 50948 4758
rect 50896 4694 50948 4700
rect 50908 4146 50936 4694
rect 51000 4690 51028 5238
rect 50988 4684 51040 4690
rect 50988 4626 51040 4632
rect 51080 4276 51132 4282
rect 51080 4218 51132 4224
rect 50896 4140 50948 4146
rect 50896 4082 50948 4088
rect 50908 3534 50936 4082
rect 50436 3528 50488 3534
rect 50436 3470 50488 3476
rect 50896 3528 50948 3534
rect 50896 3470 50948 3476
rect 49516 3392 49568 3398
rect 49516 3334 49568 3340
rect 50436 3392 50488 3398
rect 50436 3334 50488 3340
rect 49528 3194 49556 3334
rect 49516 3188 49568 3194
rect 49516 3130 49568 3136
rect 49436 2746 49556 2774
rect 48228 1352 48280 1358
rect 48228 1294 48280 1300
rect 49148 1352 49200 1358
rect 49148 1294 49200 1300
rect 47952 1216 48004 1222
rect 47952 1158 48004 1164
rect 48240 649 48268 1294
rect 49160 649 49188 1294
rect 49528 1222 49556 2746
rect 49792 1352 49844 1358
rect 49792 1294 49844 1300
rect 49516 1216 49568 1222
rect 49516 1158 49568 1164
rect 49804 649 49832 1294
rect 50448 1222 50476 3334
rect 50620 1352 50672 1358
rect 50620 1294 50672 1300
rect 50436 1216 50488 1222
rect 50436 1158 50488 1164
rect 50632 649 50660 1294
rect 51092 1222 51120 4218
rect 51184 4214 51212 8230
rect 51276 5234 51304 9318
rect 51724 7880 51776 7886
rect 51724 7822 51776 7828
rect 51632 7812 51684 7818
rect 51632 7754 51684 7760
rect 51448 6316 51500 6322
rect 51448 6258 51500 6264
rect 51460 5574 51488 6258
rect 51540 6112 51592 6118
rect 51540 6054 51592 6060
rect 51552 5710 51580 6054
rect 51540 5704 51592 5710
rect 51540 5646 51592 5652
rect 51448 5568 51500 5574
rect 51644 5522 51672 7754
rect 51448 5510 51500 5516
rect 51264 5228 51316 5234
rect 51264 5170 51316 5176
rect 51356 5228 51408 5234
rect 51356 5170 51408 5176
rect 51368 4758 51396 5170
rect 51356 4752 51408 4758
rect 51356 4694 51408 4700
rect 51172 4208 51224 4214
rect 51172 4150 51224 4156
rect 51356 1352 51408 1358
rect 51356 1294 51408 1300
rect 51080 1216 51132 1222
rect 51080 1158 51132 1164
rect 51368 649 51396 1294
rect 51460 746 51488 5510
rect 51552 5494 51672 5522
rect 51552 3466 51580 5494
rect 51736 5234 51764 7822
rect 51724 5228 51776 5234
rect 51724 5170 51776 5176
rect 51724 4208 51776 4214
rect 51724 4150 51776 4156
rect 51632 4072 51684 4078
rect 51632 4014 51684 4020
rect 51644 3641 51672 4014
rect 51630 3632 51686 3641
rect 51630 3567 51632 3576
rect 51684 3567 51686 3576
rect 51632 3538 51684 3544
rect 51540 3460 51592 3466
rect 51540 3402 51592 3408
rect 51632 3392 51684 3398
rect 51632 3334 51684 3340
rect 51448 740 51500 746
rect 51448 682 51500 688
rect 48226 640 48282 649
rect 48226 575 48282 584
rect 49146 640 49202 649
rect 49146 575 49202 584
rect 49790 640 49846 649
rect 49790 575 49846 584
rect 50618 640 50674 649
rect 50618 575 50674 584
rect 51354 640 51410 649
rect 51644 610 51672 3334
rect 51736 950 51764 4150
rect 51828 4146 51856 9386
rect 52276 9376 52328 9382
rect 52276 9318 52328 9324
rect 53104 9376 53156 9382
rect 53104 9318 53156 9324
rect 52182 7984 52238 7993
rect 52182 7919 52238 7928
rect 52000 5568 52052 5574
rect 52000 5510 52052 5516
rect 51908 4684 51960 4690
rect 51908 4626 51960 4632
rect 51816 4140 51868 4146
rect 51816 4082 51868 4088
rect 51814 3496 51870 3505
rect 51814 3431 51870 3440
rect 51828 3398 51856 3431
rect 51816 3392 51868 3398
rect 51816 3334 51868 3340
rect 51816 3120 51868 3126
rect 51816 3062 51868 3068
rect 51828 2650 51856 3062
rect 51816 2644 51868 2650
rect 51816 2586 51868 2592
rect 51920 1222 51948 4626
rect 52012 1222 52040 5510
rect 52092 5160 52144 5166
rect 52092 5102 52144 5108
rect 52104 4078 52132 5102
rect 52196 5098 52224 7919
rect 52288 5710 52316 9318
rect 53116 8974 53144 9318
rect 53300 9178 53328 10231
rect 53852 9178 53880 10231
rect 54864 9722 54892 10231
rect 54760 9716 54812 9722
rect 54760 9658 54812 9664
rect 54852 9716 54904 9722
rect 54852 9658 54904 9664
rect 54300 9648 54352 9654
rect 54576 9648 54628 9654
rect 54352 9596 54576 9602
rect 54300 9590 54628 9596
rect 54312 9574 54616 9590
rect 54668 9580 54720 9586
rect 54668 9522 54720 9528
rect 54300 9512 54352 9518
rect 54300 9454 54352 9460
rect 53288 9172 53340 9178
rect 53288 9114 53340 9120
rect 53840 9172 53892 9178
rect 53840 9114 53892 9120
rect 53104 8968 53156 8974
rect 53104 8910 53156 8916
rect 53656 8968 53708 8974
rect 53656 8910 53708 8916
rect 54116 8968 54168 8974
rect 54116 8910 54168 8916
rect 53668 8634 53696 8910
rect 54128 8838 54156 8910
rect 54116 8832 54168 8838
rect 54116 8774 54168 8780
rect 53656 8628 53708 8634
rect 53656 8570 53708 8576
rect 54128 8362 54156 8774
rect 54116 8356 54168 8362
rect 54116 8298 54168 8304
rect 52368 6316 52420 6322
rect 52368 6258 52420 6264
rect 52380 5794 52408 6258
rect 53104 6248 53156 6254
rect 53104 6190 53156 6196
rect 53746 6216 53802 6225
rect 52380 5766 52592 5794
rect 53116 5778 53144 6190
rect 53746 6151 53748 6160
rect 53800 6151 53802 6160
rect 53748 6122 53800 6128
rect 52276 5704 52328 5710
rect 52276 5646 52328 5652
rect 52368 5704 52420 5710
rect 52368 5646 52420 5652
rect 52380 5098 52408 5646
rect 52564 5574 52592 5766
rect 53104 5772 53156 5778
rect 53104 5714 53156 5720
rect 52552 5568 52604 5574
rect 52552 5510 52604 5516
rect 53012 5160 53064 5166
rect 53116 5148 53144 5714
rect 53286 5672 53342 5681
rect 53286 5607 53342 5616
rect 53300 5574 53328 5607
rect 53288 5568 53340 5574
rect 53288 5510 53340 5516
rect 53064 5120 53144 5148
rect 53012 5102 53064 5108
rect 52184 5092 52236 5098
rect 52184 5034 52236 5040
rect 52368 5092 52420 5098
rect 52368 5034 52420 5040
rect 52380 4758 52408 5034
rect 52368 4752 52420 4758
rect 52368 4694 52420 4700
rect 52092 4072 52144 4078
rect 52092 4014 52144 4020
rect 52092 3392 52144 3398
rect 52092 3334 52144 3340
rect 52104 2825 52132 3334
rect 52090 2816 52146 2825
rect 52090 2751 52146 2760
rect 53840 2440 53892 2446
rect 53840 2382 53892 2388
rect 53748 2304 53800 2310
rect 53748 2246 53800 2252
rect 53286 2136 53342 2145
rect 53286 2071 53342 2080
rect 53300 2038 53328 2071
rect 53288 2032 53340 2038
rect 53288 1974 53340 1980
rect 53300 1902 53328 1974
rect 53760 1970 53788 2246
rect 53748 1964 53800 1970
rect 53748 1906 53800 1912
rect 53288 1896 53340 1902
rect 53288 1838 53340 1844
rect 52920 1760 52972 1766
rect 52920 1702 52972 1708
rect 52092 1352 52144 1358
rect 52092 1294 52144 1300
rect 51908 1216 51960 1222
rect 51908 1158 51960 1164
rect 52000 1216 52052 1222
rect 52000 1158 52052 1164
rect 51724 944 51776 950
rect 51724 886 51776 892
rect 52104 649 52132 1294
rect 52932 649 52960 1702
rect 53852 1426 53880 2382
rect 54128 1902 54156 8298
rect 54312 2582 54340 9454
rect 54680 8974 54708 9522
rect 54772 9518 54800 9658
rect 54944 9580 54996 9586
rect 54944 9522 54996 9528
rect 54760 9512 54812 9518
rect 54760 9454 54812 9460
rect 54956 9178 54984 9522
rect 55692 9178 55720 10231
rect 56324 10192 56376 10198
rect 56324 10134 56376 10140
rect 56336 9450 56364 10134
rect 56416 10056 56468 10062
rect 56416 9998 56468 10004
rect 56324 9444 56376 9450
rect 56324 9386 56376 9392
rect 54944 9172 54996 9178
rect 54944 9114 54996 9120
rect 55680 9172 55732 9178
rect 55680 9114 55732 9120
rect 55680 9036 55732 9042
rect 55680 8978 55732 8984
rect 54668 8968 54720 8974
rect 54668 8910 54720 8916
rect 54680 8498 54708 8910
rect 55692 8498 55720 8978
rect 56336 8974 56364 9386
rect 55864 8968 55916 8974
rect 55864 8910 55916 8916
rect 56324 8968 56376 8974
rect 56324 8910 56376 8916
rect 55876 8634 55904 8910
rect 55864 8628 55916 8634
rect 55864 8570 55916 8576
rect 54668 8492 54720 8498
rect 54668 8434 54720 8440
rect 55588 8492 55640 8498
rect 55588 8434 55640 8440
rect 55680 8492 55732 8498
rect 55680 8434 55732 8440
rect 54392 8424 54444 8430
rect 54392 8366 54444 8372
rect 54300 2576 54352 2582
rect 54300 2518 54352 2524
rect 54208 2440 54260 2446
rect 54208 2382 54260 2388
rect 54220 1970 54248 2382
rect 54208 1964 54260 1970
rect 54208 1906 54260 1912
rect 54116 1896 54168 1902
rect 54116 1838 54168 1844
rect 54300 1760 54352 1766
rect 54300 1702 54352 1708
rect 54312 1562 54340 1702
rect 54300 1556 54352 1562
rect 54300 1498 54352 1504
rect 54298 1456 54354 1465
rect 53840 1420 53892 1426
rect 54404 1442 54432 8366
rect 54668 3052 54720 3058
rect 54668 2994 54720 3000
rect 54484 2848 54536 2854
rect 54484 2790 54536 2796
rect 54354 1414 54432 1442
rect 54298 1391 54300 1400
rect 53840 1362 53892 1368
rect 54352 1391 54354 1400
rect 54300 1362 54352 1368
rect 53104 1352 53156 1358
rect 53104 1294 53156 1300
rect 52090 640 52146 649
rect 51354 575 51410 584
rect 51632 604 51684 610
rect 52090 575 52146 584
rect 52918 640 52974 649
rect 52918 575 52974 584
rect 51632 546 51684 552
rect 47860 536 47912 542
rect 47860 478 47912 484
rect 40040 400 40092 406
rect 38842 368 38898 377
rect 53116 377 53144 1294
rect 54496 649 54524 2790
rect 54576 1964 54628 1970
rect 54576 1906 54628 1912
rect 54588 1358 54616 1906
rect 54680 1358 54708 2994
rect 55126 2816 55182 2825
rect 55182 2774 55260 2802
rect 55126 2751 55182 2760
rect 55232 2650 55260 2774
rect 55220 2644 55272 2650
rect 55220 2586 55272 2592
rect 55496 2440 55548 2446
rect 55496 2382 55548 2388
rect 55508 2038 55536 2382
rect 55496 2032 55548 2038
rect 55496 1974 55548 1980
rect 55600 1834 55628 8434
rect 55864 6792 55916 6798
rect 55864 6734 55916 6740
rect 55772 6384 55824 6390
rect 55772 6326 55824 6332
rect 55784 5914 55812 6326
rect 55772 5908 55824 5914
rect 55772 5850 55824 5856
rect 55876 5710 55904 6734
rect 55864 5704 55916 5710
rect 55864 5646 55916 5652
rect 55864 5092 55916 5098
rect 55864 5034 55916 5040
rect 55876 4826 55904 5034
rect 55864 4820 55916 4826
rect 55864 4762 55916 4768
rect 55864 4548 55916 4554
rect 55864 4490 55916 4496
rect 55876 4282 55904 4490
rect 55864 4276 55916 4282
rect 55864 4218 55916 4224
rect 56336 2774 56364 8910
rect 56428 8634 56456 9998
rect 56520 9722 56548 10231
rect 56876 10124 56928 10130
rect 56876 10066 56928 10072
rect 56508 9716 56560 9722
rect 56508 9658 56560 9664
rect 56600 9580 56652 9586
rect 56600 9522 56652 9528
rect 56612 9178 56640 9522
rect 56600 9172 56652 9178
rect 56600 9114 56652 9120
rect 56888 8974 56916 10066
rect 57348 9722 57376 10231
rect 57808 9722 57836 10231
rect 57336 9716 57388 9722
rect 57336 9658 57388 9664
rect 57796 9716 57848 9722
rect 57796 9658 57848 9664
rect 57336 9580 57388 9586
rect 57336 9522 57388 9528
rect 58072 9580 58124 9586
rect 58072 9522 58124 9528
rect 57152 9036 57204 9042
rect 57152 8978 57204 8984
rect 56876 8968 56928 8974
rect 56876 8910 56928 8916
rect 56888 8838 56916 8910
rect 56876 8832 56928 8838
rect 56876 8774 56928 8780
rect 56416 8628 56468 8634
rect 56416 8570 56468 8576
rect 56428 8430 56456 8570
rect 56416 8424 56468 8430
rect 56416 8366 56468 8372
rect 56244 2746 56364 2774
rect 56244 2038 56272 2746
rect 56232 2032 56284 2038
rect 56232 1974 56284 1980
rect 56428 1970 56456 8366
rect 56888 1970 56916 8774
rect 57164 8498 57192 8978
rect 57348 8634 57376 9522
rect 58084 9178 58112 9522
rect 58544 9178 58572 10270
rect 58806 10231 58862 10240
rect 59266 10296 59322 10305
rect 59266 10231 59322 10240
rect 60278 10296 60334 10305
rect 60278 10231 60334 10240
rect 58072 9172 58124 9178
rect 58072 9114 58124 9120
rect 58532 9172 58584 9178
rect 58532 9114 58584 9120
rect 57980 9104 58032 9110
rect 57980 9046 58032 9052
rect 57992 8974 58020 9046
rect 58544 8974 58572 9114
rect 57980 8968 58032 8974
rect 57980 8910 58032 8916
rect 58532 8968 58584 8974
rect 58532 8910 58584 8916
rect 57428 8832 57480 8838
rect 57428 8774 57480 8780
rect 57336 8628 57388 8634
rect 57336 8570 57388 8576
rect 57152 8492 57204 8498
rect 57152 8434 57204 8440
rect 57336 8492 57388 8498
rect 57336 8434 57388 8440
rect 57348 8362 57376 8434
rect 57440 8362 57468 8774
rect 57336 8356 57388 8362
rect 57336 8298 57388 8304
rect 57428 8356 57480 8362
rect 57428 8298 57480 8304
rect 57992 2774 58020 8910
rect 58256 8832 58308 8838
rect 58256 8774 58308 8780
rect 58268 8498 58296 8774
rect 58256 8492 58308 8498
rect 58256 8434 58308 8440
rect 58544 2774 58572 8910
rect 58820 8634 58848 10231
rect 59280 8634 59308 10231
rect 59728 9988 59780 9994
rect 59728 9930 59780 9936
rect 59740 9450 59768 9930
rect 59728 9444 59780 9450
rect 59728 9386 59780 9392
rect 59740 8974 59768 9386
rect 59912 9376 59964 9382
rect 59912 9318 59964 9324
rect 59924 8974 59952 9318
rect 59728 8968 59780 8974
rect 59728 8910 59780 8916
rect 59912 8968 59964 8974
rect 59912 8910 59964 8916
rect 59360 8832 59412 8838
rect 59360 8774 59412 8780
rect 58808 8628 58860 8634
rect 58808 8570 58860 8576
rect 59268 8628 59320 8634
rect 59268 8570 59320 8576
rect 59372 8498 59400 8774
rect 59360 8492 59412 8498
rect 59360 8434 59412 8440
rect 57992 2746 58204 2774
rect 58544 2746 58664 2774
rect 57520 2440 57572 2446
rect 57520 2382 57572 2388
rect 57532 2038 57560 2382
rect 57980 2304 58032 2310
rect 57980 2246 58032 2252
rect 57520 2032 57572 2038
rect 57520 1974 57572 1980
rect 56416 1964 56468 1970
rect 56416 1906 56468 1912
rect 56876 1964 56928 1970
rect 56876 1906 56928 1912
rect 55588 1828 55640 1834
rect 55588 1770 55640 1776
rect 55036 1760 55088 1766
rect 55036 1702 55088 1708
rect 56232 1760 56284 1766
rect 56232 1702 56284 1708
rect 56968 1760 57020 1766
rect 56968 1702 57020 1708
rect 55048 1358 55076 1702
rect 56244 1358 56272 1702
rect 56980 1358 57008 1702
rect 57992 1601 58020 2246
rect 58072 1964 58124 1970
rect 58072 1906 58124 1912
rect 57978 1592 58034 1601
rect 58084 1562 58112 1906
rect 57978 1527 58034 1536
rect 58072 1556 58124 1562
rect 58072 1498 58124 1504
rect 58176 1426 58204 2746
rect 58636 1970 58664 2746
rect 59176 2440 59228 2446
rect 59176 2382 59228 2388
rect 59188 2038 59216 2382
rect 59360 2304 59412 2310
rect 59360 2246 59412 2252
rect 59176 2032 59228 2038
rect 59176 1974 59228 1980
rect 58624 1964 58676 1970
rect 58624 1906 58676 1912
rect 58532 1896 58584 1902
rect 58532 1838 58584 1844
rect 58256 1760 58308 1766
rect 58256 1702 58308 1708
rect 58164 1420 58216 1426
rect 58164 1362 58216 1368
rect 54576 1352 54628 1358
rect 54576 1294 54628 1300
rect 54668 1352 54720 1358
rect 54668 1294 54720 1300
rect 55036 1352 55088 1358
rect 55036 1294 55088 1300
rect 56232 1352 56284 1358
rect 56232 1294 56284 1300
rect 56968 1352 57020 1358
rect 56968 1294 57020 1300
rect 55680 1216 55732 1222
rect 55680 1158 55732 1164
rect 56416 1216 56468 1222
rect 56416 1158 56468 1164
rect 57152 1216 57204 1222
rect 57152 1158 57204 1164
rect 54482 640 54538 649
rect 54482 575 54538 584
rect 55692 513 55720 1158
rect 56428 513 56456 1158
rect 57164 513 57192 1158
rect 58268 513 58296 1702
rect 58544 1358 58572 1838
rect 59372 1601 59400 2246
rect 59740 1970 59768 8910
rect 60096 8832 60148 8838
rect 60096 8774 60148 8780
rect 60108 8498 60136 8774
rect 60292 8634 60320 10231
rect 60660 9654 60688 10610
rect 62028 10464 62080 10470
rect 62028 10406 62080 10412
rect 61014 10296 61070 10305
rect 61014 10231 61070 10240
rect 61750 10296 61806 10305
rect 61750 10231 61806 10240
rect 60648 9648 60700 9654
rect 60648 9590 60700 9596
rect 60660 9042 60688 9590
rect 60648 9036 60700 9042
rect 60648 8978 60700 8984
rect 60660 8634 60688 8978
rect 60832 8832 60884 8838
rect 60832 8774 60884 8780
rect 60280 8628 60332 8634
rect 60280 8570 60332 8576
rect 60648 8628 60700 8634
rect 60648 8570 60700 8576
rect 60096 8492 60148 8498
rect 60096 8434 60148 8440
rect 60660 2774 60688 8570
rect 60844 8498 60872 8774
rect 60832 8492 60884 8498
rect 60832 8434 60884 8440
rect 61028 8294 61056 10231
rect 61476 10056 61528 10062
rect 61476 9998 61528 10004
rect 61488 8974 61516 9998
rect 61764 9722 61792 10231
rect 61752 9716 61804 9722
rect 61752 9658 61804 9664
rect 61476 8968 61528 8974
rect 61476 8910 61528 8916
rect 61488 8838 61516 8910
rect 61476 8832 61528 8838
rect 61476 8774 61528 8780
rect 61488 8430 61516 8774
rect 62040 8498 62068 10406
rect 63224 10328 63276 10334
rect 62486 10296 62542 10305
rect 63224 10270 63276 10276
rect 63406 10296 63462 10305
rect 62486 10231 62542 10240
rect 62500 9722 62528 10231
rect 62488 9716 62540 9722
rect 62488 9658 62540 9664
rect 62212 9580 62264 9586
rect 62212 9522 62264 9528
rect 62580 9580 62632 9586
rect 62580 9522 62632 9528
rect 62764 9580 62816 9586
rect 62764 9522 62816 9528
rect 62224 9178 62252 9522
rect 62212 9172 62264 9178
rect 62212 9114 62264 9120
rect 62304 9104 62356 9110
rect 62304 9046 62356 9052
rect 62316 8906 62344 9046
rect 62488 8968 62540 8974
rect 62488 8910 62540 8916
rect 62304 8900 62356 8906
rect 62304 8842 62356 8848
rect 62028 8492 62080 8498
rect 62028 8434 62080 8440
rect 61292 8424 61344 8430
rect 61292 8366 61344 8372
rect 61476 8424 61528 8430
rect 61476 8366 61528 8372
rect 61016 8288 61068 8294
rect 61016 8230 61068 8236
rect 60568 2746 60688 2774
rect 59820 2304 59872 2310
rect 59820 2246 59872 2252
rect 59832 1970 59860 2246
rect 60568 1970 60596 2746
rect 61304 1970 61332 8366
rect 61660 2440 61712 2446
rect 61660 2382 61712 2388
rect 61476 2304 61528 2310
rect 61476 2246 61528 2252
rect 59728 1964 59780 1970
rect 59728 1906 59780 1912
rect 59820 1964 59872 1970
rect 59820 1906 59872 1912
rect 60556 1964 60608 1970
rect 60556 1906 60608 1912
rect 61292 1964 61344 1970
rect 61292 1906 61344 1912
rect 59820 1760 59872 1766
rect 59820 1702 59872 1708
rect 60740 1760 60792 1766
rect 60740 1702 60792 1708
rect 59358 1592 59414 1601
rect 59358 1527 59414 1536
rect 59542 1592 59598 1601
rect 59542 1527 59598 1536
rect 59556 1426 59584 1527
rect 59544 1420 59596 1426
rect 59544 1362 59596 1368
rect 59832 1358 59860 1702
rect 60752 1358 60780 1702
rect 58532 1352 58584 1358
rect 58532 1294 58584 1300
rect 59820 1352 59872 1358
rect 59820 1294 59872 1300
rect 60740 1352 60792 1358
rect 60740 1294 60792 1300
rect 60004 1216 60056 1222
rect 60004 1158 60056 1164
rect 60924 1216 60976 1222
rect 60924 1158 60976 1164
rect 60016 513 60044 1158
rect 60936 513 60964 1158
rect 61488 513 61516 2246
rect 61672 2038 61700 2382
rect 61660 2032 61712 2038
rect 61660 1974 61712 1980
rect 62040 1426 62068 8434
rect 62212 2440 62264 2446
rect 62212 2382 62264 2388
rect 62224 1562 62252 2382
rect 62316 1970 62344 8842
rect 62500 8498 62528 8910
rect 62592 8634 62620 9522
rect 62776 9178 62804 9522
rect 62764 9172 62816 9178
rect 62764 9114 62816 9120
rect 63236 8974 63264 10270
rect 63406 10231 63462 10240
rect 63958 10296 64014 10305
rect 63958 10231 64014 10240
rect 64694 10296 64750 10305
rect 64694 10231 64750 10240
rect 65522 10296 65578 10305
rect 65522 10231 65578 10240
rect 65890 10296 65946 10305
rect 65890 10231 65946 10240
rect 67178 10296 67234 10305
rect 67178 10231 67234 10240
rect 63420 9722 63448 10231
rect 63408 9716 63460 9722
rect 63408 9658 63460 9664
rect 63224 8968 63276 8974
rect 63224 8910 63276 8916
rect 62672 8900 62724 8906
rect 62672 8842 62724 8848
rect 62580 8628 62632 8634
rect 62580 8570 62632 8576
rect 62488 8492 62540 8498
rect 62488 8434 62540 8440
rect 62684 8362 62712 8842
rect 62672 8356 62724 8362
rect 62672 8298 62724 8304
rect 62672 2440 62724 2446
rect 62672 2382 62724 2388
rect 62396 2304 62448 2310
rect 62396 2246 62448 2252
rect 62304 1964 62356 1970
rect 62304 1906 62356 1912
rect 62212 1556 62264 1562
rect 62212 1498 62264 1504
rect 62028 1420 62080 1426
rect 62028 1362 62080 1368
rect 62408 513 62436 2246
rect 62684 2038 62712 2382
rect 63132 2304 63184 2310
rect 63132 2246 63184 2252
rect 62672 2032 62724 2038
rect 62672 1974 62724 1980
rect 62488 1964 62540 1970
rect 62488 1906 62540 1912
rect 62500 1358 62528 1906
rect 62488 1352 62540 1358
rect 62488 1294 62540 1300
rect 63144 513 63172 2246
rect 63236 1970 63264 8910
rect 63776 8832 63828 8838
rect 63776 8774 63828 8780
rect 63788 8498 63816 8774
rect 63972 8634 64000 10231
rect 64052 9920 64104 9926
rect 64052 9862 64104 9868
rect 64064 9178 64092 9862
rect 64052 9172 64104 9178
rect 64052 9114 64104 9120
rect 64064 8974 64092 9114
rect 64052 8968 64104 8974
rect 64052 8910 64104 8916
rect 63960 8628 64012 8634
rect 63960 8570 64012 8576
rect 63776 8492 63828 8498
rect 63776 8434 63828 8440
rect 64064 1970 64092 8910
rect 64512 8832 64564 8838
rect 64512 8774 64564 8780
rect 64524 8498 64552 8774
rect 64708 8634 64736 10231
rect 64972 8968 65024 8974
rect 64972 8910 65024 8916
rect 64696 8628 64748 8634
rect 64696 8570 64748 8576
rect 64512 8492 64564 8498
rect 64512 8434 64564 8440
rect 64984 6914 65012 8910
rect 65340 8832 65392 8838
rect 65340 8774 65392 8780
rect 65352 8498 65380 8774
rect 65340 8492 65392 8498
rect 65340 8434 65392 8440
rect 65536 8362 65564 10231
rect 65904 8362 65932 10231
rect 66076 9512 66128 9518
rect 66076 9454 66128 9460
rect 65984 9036 66036 9042
rect 65984 8978 66036 8984
rect 65996 8566 66024 8978
rect 66088 8974 66116 9454
rect 66076 8968 66128 8974
rect 66352 8968 66404 8974
rect 66128 8928 66352 8956
rect 66076 8910 66128 8916
rect 66076 8832 66128 8838
rect 66076 8774 66128 8780
rect 65984 8560 66036 8566
rect 65984 8502 66036 8508
rect 66088 8498 66116 8774
rect 66076 8492 66128 8498
rect 66076 8434 66128 8440
rect 65524 8356 65576 8362
rect 65524 8298 65576 8304
rect 65892 8356 65944 8362
rect 65892 8298 65944 8304
rect 66180 6914 66208 8928
rect 66352 8910 66404 8916
rect 66996 8968 67048 8974
rect 66996 8910 67048 8916
rect 67008 8090 67036 8910
rect 67192 8838 67220 10231
rect 68546 9820 68854 9829
rect 68546 9818 68552 9820
rect 68608 9818 68632 9820
rect 68688 9818 68712 9820
rect 68768 9818 68792 9820
rect 68848 9818 68854 9820
rect 68608 9766 68610 9818
rect 68790 9766 68792 9818
rect 68546 9764 68552 9766
rect 68608 9764 68632 9766
rect 68688 9764 68712 9766
rect 68768 9764 68792 9766
rect 68848 9764 68854 9766
rect 68546 9755 68854 9764
rect 67364 9648 67416 9654
rect 67364 9590 67416 9596
rect 69110 9616 69166 9625
rect 67180 8832 67232 8838
rect 67180 8774 67232 8780
rect 67088 8560 67140 8566
rect 67088 8502 67140 8508
rect 66996 8084 67048 8090
rect 66996 8026 67048 8032
rect 67100 7886 67128 8502
rect 67376 8430 67404 9590
rect 69110 9551 69112 9560
rect 69164 9551 69166 9560
rect 69112 9522 69164 9528
rect 69860 9518 69888 10746
rect 82096 10674 82124 10814
rect 93952 10804 94004 10810
rect 93952 10746 94004 10752
rect 92388 10736 92440 10742
rect 92388 10678 92440 10684
rect 82084 10668 82136 10674
rect 82084 10610 82136 10616
rect 81622 10568 81678 10577
rect 81622 10503 81678 10512
rect 82634 10568 82690 10577
rect 82634 10503 82690 10512
rect 86774 10568 86830 10577
rect 86774 10503 86830 10512
rect 91008 10532 91060 10538
rect 74540 10464 74592 10470
rect 72054 10432 72110 10441
rect 74540 10406 74592 10412
rect 72054 10367 72110 10376
rect 71502 10160 71558 10169
rect 71502 10095 71558 10104
rect 70030 9888 70086 9897
rect 70030 9823 70086 9832
rect 69848 9512 69900 9518
rect 69848 9454 69900 9460
rect 70044 8974 70072 9823
rect 70306 9616 70362 9625
rect 71516 9586 71544 10095
rect 70306 9551 70308 9560
rect 70360 9551 70362 9560
rect 71504 9580 71556 9586
rect 70308 9522 70360 9528
rect 71504 9522 71556 9528
rect 72068 9042 72096 10367
rect 72146 9616 72202 9625
rect 72146 9551 72148 9560
rect 72200 9551 72202 9560
rect 74262 9616 74318 9625
rect 74262 9551 74318 9560
rect 72148 9522 72200 9528
rect 73712 9444 73764 9450
rect 73712 9386 73764 9392
rect 73724 9178 73752 9386
rect 73712 9172 73764 9178
rect 73712 9114 73764 9120
rect 73434 9072 73490 9081
rect 70400 9036 70452 9042
rect 70400 8978 70452 8984
rect 72056 9036 72108 9042
rect 73434 9007 73436 9016
rect 72056 8978 72108 8984
rect 73488 9007 73490 9016
rect 73436 8978 73488 8984
rect 70032 8968 70084 8974
rect 70032 8910 70084 8916
rect 68546 8732 68854 8741
rect 68546 8730 68552 8732
rect 68608 8730 68632 8732
rect 68688 8730 68712 8732
rect 68768 8730 68792 8732
rect 68848 8730 68854 8732
rect 68608 8678 68610 8730
rect 68790 8678 68792 8730
rect 68546 8676 68552 8678
rect 68608 8676 68632 8678
rect 68688 8676 68712 8678
rect 68768 8676 68792 8678
rect 68848 8676 68854 8678
rect 68546 8667 68854 8676
rect 67364 8424 67416 8430
rect 67364 8366 67416 8372
rect 70412 8294 70440 8978
rect 72332 8968 72384 8974
rect 72332 8910 72384 8916
rect 73712 8968 73764 8974
rect 73712 8910 73764 8916
rect 70400 8288 70452 8294
rect 70400 8230 70452 8236
rect 67088 7880 67140 7886
rect 67088 7822 67140 7828
rect 68546 7644 68854 7653
rect 68546 7642 68552 7644
rect 68608 7642 68632 7644
rect 68688 7642 68712 7644
rect 68768 7642 68792 7644
rect 68848 7642 68854 7644
rect 68608 7590 68610 7642
rect 68790 7590 68792 7642
rect 68546 7588 68552 7590
rect 68608 7588 68632 7590
rect 68688 7588 68712 7590
rect 68768 7588 68792 7590
rect 68848 7588 68854 7590
rect 68546 7579 68854 7588
rect 64984 6886 65104 6914
rect 65076 2417 65104 6886
rect 66088 6886 66208 6914
rect 65432 2440 65484 2446
rect 65062 2408 65118 2417
rect 65432 2382 65484 2388
rect 65062 2343 65118 2352
rect 63224 1964 63276 1970
rect 63224 1906 63276 1912
rect 64052 1964 64104 1970
rect 64052 1906 64104 1912
rect 65076 1902 65104 2343
rect 65444 2038 65472 2382
rect 65984 2304 66036 2310
rect 65984 2246 66036 2252
rect 65432 2032 65484 2038
rect 65432 1974 65484 1980
rect 65064 1896 65116 1902
rect 65064 1838 65116 1844
rect 63684 1760 63736 1766
rect 63684 1702 63736 1708
rect 64420 1760 64472 1766
rect 64420 1702 64472 1708
rect 63696 1358 63724 1702
rect 64432 1358 64460 1702
rect 65076 1494 65104 1838
rect 65064 1488 65116 1494
rect 65064 1430 65116 1436
rect 63684 1352 63736 1358
rect 63684 1294 63736 1300
rect 64420 1352 64472 1358
rect 64420 1294 64472 1300
rect 63868 1216 63920 1222
rect 63868 1158 63920 1164
rect 64604 1216 64656 1222
rect 64604 1158 64656 1164
rect 65892 1216 65944 1222
rect 65892 1158 65944 1164
rect 55678 504 55734 513
rect 55678 439 55734 448
rect 56414 504 56470 513
rect 56414 439 56470 448
rect 57150 504 57206 513
rect 57150 439 57206 448
rect 58254 504 58310 513
rect 58254 439 58310 448
rect 60002 504 60058 513
rect 60002 439 60058 448
rect 60922 504 60978 513
rect 60922 439 60978 448
rect 61474 504 61530 513
rect 61474 439 61530 448
rect 62394 504 62450 513
rect 62394 439 62450 448
rect 63130 504 63186 513
rect 63130 439 63186 448
rect 63880 377 63908 1158
rect 64616 377 64644 1158
rect 65904 513 65932 1158
rect 65890 504 65946 513
rect 65890 439 65946 448
rect 65996 377 66024 2246
rect 66088 1426 66116 6886
rect 68546 6556 68854 6565
rect 68546 6554 68552 6556
rect 68608 6554 68632 6556
rect 68688 6554 68712 6556
rect 68768 6554 68792 6556
rect 68848 6554 68854 6556
rect 68608 6502 68610 6554
rect 68790 6502 68792 6554
rect 68546 6500 68552 6502
rect 68608 6500 68632 6502
rect 68688 6500 68712 6502
rect 68768 6500 68792 6502
rect 68848 6500 68854 6502
rect 68546 6491 68854 6500
rect 72344 6458 72372 8910
rect 73724 7954 73752 8910
rect 74276 8498 74304 9551
rect 74552 8498 74580 10406
rect 80612 10396 80664 10402
rect 80612 10338 80664 10344
rect 80624 10198 80652 10338
rect 80612 10192 80664 10198
rect 79230 10160 79286 10169
rect 80612 10134 80664 10140
rect 81072 10192 81124 10198
rect 81072 10134 81124 10140
rect 79230 10095 79286 10104
rect 77206 9888 77262 9897
rect 77206 9823 77262 9832
rect 78678 9888 78734 9897
rect 78678 9823 78734 9832
rect 76380 9648 76432 9654
rect 74722 9616 74778 9625
rect 76380 9590 76432 9596
rect 76470 9616 76526 9625
rect 74722 9551 74724 9560
rect 74776 9551 74778 9560
rect 74724 9522 74776 9528
rect 75828 9512 75880 9518
rect 75828 9454 75880 9460
rect 74722 9072 74778 9081
rect 74722 9007 74778 9016
rect 74736 8974 74764 9007
rect 74724 8968 74776 8974
rect 74724 8910 74776 8916
rect 75000 8968 75052 8974
rect 75000 8910 75052 8916
rect 74264 8492 74316 8498
rect 74264 8434 74316 8440
rect 74540 8492 74592 8498
rect 74540 8434 74592 8440
rect 75012 8022 75040 8910
rect 75000 8016 75052 8022
rect 75000 7958 75052 7964
rect 73712 7948 73764 7954
rect 73712 7890 73764 7896
rect 75840 7721 75868 9454
rect 75826 7712 75882 7721
rect 75826 7647 75882 7656
rect 76392 7546 76420 9590
rect 76470 9551 76526 9560
rect 76484 8498 76512 9551
rect 77220 8974 77248 9823
rect 77298 9616 77354 9625
rect 77298 9551 77300 9560
rect 77352 9551 77354 9560
rect 77300 9522 77352 9528
rect 77576 9512 77628 9518
rect 77576 9454 77628 9460
rect 77208 8968 77260 8974
rect 77208 8910 77260 8916
rect 77484 8968 77536 8974
rect 77484 8910 77536 8916
rect 76472 8492 76524 8498
rect 76472 8434 76524 8440
rect 76380 7540 76432 7546
rect 76380 7482 76432 7488
rect 76562 7440 76618 7449
rect 76562 7375 76564 7384
rect 76616 7375 76618 7384
rect 76564 7346 76616 7352
rect 72332 6452 72384 6458
rect 72332 6394 72384 6400
rect 77496 5642 77524 8910
rect 77588 8090 77616 9454
rect 78692 8974 78720 9823
rect 79244 9654 79272 10095
rect 79232 9648 79284 9654
rect 79232 9590 79284 9596
rect 79966 9616 80022 9625
rect 79966 9551 79968 9560
rect 80020 9551 80022 9560
rect 79968 9522 80020 9528
rect 80152 9512 80204 9518
rect 80152 9454 80204 9460
rect 78680 8968 78732 8974
rect 78680 8910 78732 8916
rect 78956 8968 79008 8974
rect 78956 8910 79008 8916
rect 77576 8084 77628 8090
rect 77576 8026 77628 8032
rect 78772 7404 78824 7410
rect 78772 7346 78824 7352
rect 78784 7313 78812 7346
rect 78770 7304 78826 7313
rect 78770 7239 78826 7248
rect 78968 6361 78996 8910
rect 80164 7585 80192 9454
rect 81084 9110 81112 10134
rect 81532 9988 81584 9994
rect 81532 9930 81584 9936
rect 81254 9888 81310 9897
rect 81254 9823 81310 9832
rect 81072 9104 81124 9110
rect 81072 9046 81124 9052
rect 81268 9042 81296 9823
rect 81544 9042 81572 9930
rect 81636 9586 81664 10503
rect 81624 9580 81676 9586
rect 81624 9522 81676 9528
rect 81256 9036 81308 9042
rect 81256 8978 81308 8984
rect 81532 9036 81584 9042
rect 81532 8978 81584 8984
rect 82648 8974 82676 10503
rect 83094 10160 83150 10169
rect 83094 10095 83150 10104
rect 83922 10160 83978 10169
rect 83922 10095 83978 10104
rect 84658 10160 84714 10169
rect 84658 10095 84714 10104
rect 85394 10160 85450 10169
rect 85394 10095 85450 10104
rect 83108 9654 83136 10095
rect 83188 9716 83240 9722
rect 83188 9658 83240 9664
rect 83096 9648 83148 9654
rect 83096 9590 83148 9596
rect 82820 9036 82872 9042
rect 82820 8978 82872 8984
rect 82636 8968 82688 8974
rect 82636 8910 82688 8916
rect 82728 8424 82780 8430
rect 82728 8366 82780 8372
rect 80150 7576 80206 7585
rect 80150 7511 80206 7520
rect 82740 6633 82768 8366
rect 82832 6662 82860 8978
rect 83200 6730 83228 9658
rect 83936 9654 83964 10095
rect 84016 9920 84068 9926
rect 84016 9862 84068 9868
rect 84028 9722 84056 9862
rect 84016 9716 84068 9722
rect 84016 9658 84068 9664
rect 84672 9654 84700 10095
rect 85408 9654 85436 10095
rect 86406 9888 86462 9897
rect 86406 9823 86462 9832
rect 83924 9648 83976 9654
rect 83924 9590 83976 9596
rect 84660 9648 84712 9654
rect 84660 9590 84712 9596
rect 85396 9648 85448 9654
rect 85396 9590 85448 9596
rect 83280 9444 83332 9450
rect 83280 9386 83332 9392
rect 85488 9444 85540 9450
rect 85488 9386 85540 9392
rect 83292 7818 83320 9386
rect 84844 9172 84896 9178
rect 84844 9114 84896 9120
rect 84856 8430 84884 9114
rect 84844 8424 84896 8430
rect 84844 8366 84896 8372
rect 84108 8084 84160 8090
rect 84108 8026 84160 8032
rect 83280 7812 83332 7818
rect 83280 7754 83332 7760
rect 83188 6724 83240 6730
rect 83188 6666 83240 6672
rect 82820 6656 82872 6662
rect 82726 6624 82782 6633
rect 82820 6598 82872 6604
rect 82726 6559 82782 6568
rect 84120 6497 84148 8026
rect 85500 7857 85528 9386
rect 86420 9042 86448 9823
rect 86788 9586 86816 10503
rect 91008 10474 91060 10480
rect 91020 10402 91048 10474
rect 90732 10396 90784 10402
rect 90732 10338 90784 10344
rect 91008 10396 91060 10402
rect 91008 10338 91060 10344
rect 90362 10296 90418 10305
rect 90362 10231 90418 10240
rect 86776 9580 86828 9586
rect 86776 9522 86828 9528
rect 89444 9580 89496 9586
rect 89444 9522 89496 9528
rect 90088 9580 90140 9586
rect 90088 9522 90140 9528
rect 88984 9512 89036 9518
rect 88984 9454 89036 9460
rect 89350 9480 89406 9489
rect 88340 9376 88392 9382
rect 88340 9318 88392 9324
rect 88800 9376 88852 9382
rect 88800 9318 88852 9324
rect 88246 9208 88302 9217
rect 88246 9143 88248 9152
rect 88300 9143 88302 9152
rect 88248 9114 88300 9120
rect 86408 9036 86460 9042
rect 86408 8978 86460 8984
rect 86684 8968 86736 8974
rect 86684 8910 86736 8916
rect 86696 8090 86724 8910
rect 87510 8664 87566 8673
rect 87510 8599 87512 8608
rect 87564 8599 87566 8608
rect 87512 8570 87564 8576
rect 86684 8084 86736 8090
rect 86684 8026 86736 8032
rect 85486 7848 85542 7857
rect 85486 7783 85542 7792
rect 84200 7404 84252 7410
rect 84200 7346 84252 7352
rect 84106 6488 84162 6497
rect 84106 6423 84162 6432
rect 78954 6352 79010 6361
rect 78954 6287 79010 6296
rect 80244 6316 80296 6322
rect 80244 6258 80296 6264
rect 77484 5636 77536 5642
rect 77484 5578 77536 5584
rect 68546 5468 68854 5477
rect 68546 5466 68552 5468
rect 68608 5466 68632 5468
rect 68688 5466 68712 5468
rect 68768 5466 68792 5468
rect 68848 5466 68854 5468
rect 68608 5414 68610 5466
rect 68790 5414 68792 5466
rect 68546 5412 68552 5414
rect 68608 5412 68632 5414
rect 68688 5412 68712 5414
rect 68768 5412 68792 5414
rect 68848 5412 68854 5414
rect 68546 5403 68854 5412
rect 80058 4448 80114 4457
rect 68546 4380 68854 4389
rect 80058 4383 80114 4392
rect 68546 4378 68552 4380
rect 68608 4378 68632 4380
rect 68688 4378 68712 4380
rect 68768 4378 68792 4380
rect 68848 4378 68854 4380
rect 68608 4326 68610 4378
rect 68790 4326 68792 4378
rect 68546 4324 68552 4326
rect 68608 4324 68632 4326
rect 68688 4324 68712 4326
rect 68768 4324 68792 4326
rect 68848 4324 68854 4326
rect 68546 4315 68854 4324
rect 66720 3936 66772 3942
rect 66720 3878 66772 3884
rect 66352 2984 66404 2990
rect 66352 2926 66404 2932
rect 66168 2508 66220 2514
rect 66168 2450 66220 2456
rect 66180 2038 66208 2450
rect 66168 2032 66220 2038
rect 66168 1974 66220 1980
rect 66076 1420 66128 1426
rect 66076 1362 66128 1368
rect 66180 1358 66208 1974
rect 66364 1970 66392 2926
rect 66732 2446 66760 3878
rect 67640 3664 67692 3670
rect 67640 3606 67692 3612
rect 78586 3632 78642 3641
rect 67652 3097 67680 3606
rect 78586 3567 78642 3576
rect 68546 3292 68854 3301
rect 68546 3290 68552 3292
rect 68608 3290 68632 3292
rect 68688 3290 68712 3292
rect 68768 3290 68792 3292
rect 68848 3290 68854 3292
rect 68608 3238 68610 3290
rect 68790 3238 68792 3290
rect 68546 3236 68552 3238
rect 68608 3236 68632 3238
rect 68688 3236 68712 3238
rect 68768 3236 68792 3238
rect 68848 3236 68854 3238
rect 68546 3227 68854 3236
rect 67638 3088 67694 3097
rect 67638 3023 67694 3032
rect 66720 2440 66772 2446
rect 66720 2382 66772 2388
rect 76472 2440 76524 2446
rect 76472 2382 76524 2388
rect 68546 2204 68854 2213
rect 68546 2202 68552 2204
rect 68608 2202 68632 2204
rect 68688 2202 68712 2204
rect 68768 2202 68792 2204
rect 68848 2202 68854 2204
rect 68608 2150 68610 2202
rect 68790 2150 68792 2202
rect 68546 2148 68552 2150
rect 68608 2148 68632 2150
rect 68688 2148 68712 2150
rect 68768 2148 68792 2150
rect 68848 2148 68854 2150
rect 68546 2139 68854 2148
rect 73436 2100 73488 2106
rect 73620 2100 73672 2106
rect 73488 2060 73620 2088
rect 73436 2042 73488 2048
rect 73620 2042 73672 2048
rect 66352 1964 66404 1970
rect 66352 1906 66404 1912
rect 71504 1964 71556 1970
rect 71504 1906 71556 1912
rect 72240 1964 72292 1970
rect 73620 1964 73672 1970
rect 72240 1906 72292 1912
rect 73356 1924 73620 1952
rect 67272 1760 67324 1766
rect 67272 1702 67324 1708
rect 66168 1352 66220 1358
rect 66168 1294 66220 1300
rect 67284 513 67312 1702
rect 69112 1420 69164 1426
rect 69112 1362 69164 1368
rect 68546 1116 68854 1125
rect 68546 1114 68552 1116
rect 68608 1114 68632 1116
rect 68688 1114 68712 1116
rect 68768 1114 68792 1116
rect 68848 1114 68854 1116
rect 68608 1062 68610 1114
rect 68790 1062 68792 1114
rect 68546 1060 68552 1062
rect 68608 1060 68632 1062
rect 68688 1060 68712 1062
rect 68768 1060 68792 1062
rect 68848 1060 68854 1062
rect 68546 1051 68854 1060
rect 69124 921 69152 1362
rect 69572 1352 69624 1358
rect 69572 1294 69624 1300
rect 70952 1352 71004 1358
rect 70952 1294 71004 1300
rect 69584 921 69612 1294
rect 70964 921 70992 1294
rect 71516 1057 71544 1906
rect 72054 1864 72110 1873
rect 72054 1799 72056 1808
rect 72108 1799 72110 1808
rect 72056 1770 72108 1776
rect 72252 1057 72280 1906
rect 73356 1766 73384 1924
rect 73620 1906 73672 1912
rect 73712 1964 73764 1970
rect 73712 1906 73764 1912
rect 73436 1828 73488 1834
rect 73436 1770 73488 1776
rect 73344 1760 73396 1766
rect 73344 1702 73396 1708
rect 73448 1562 73476 1770
rect 73436 1556 73488 1562
rect 73436 1498 73488 1504
rect 72976 1352 73028 1358
rect 72976 1294 73028 1300
rect 72792 1216 72844 1222
rect 72792 1158 72844 1164
rect 71502 1048 71558 1057
rect 71502 983 71558 992
rect 72238 1048 72294 1057
rect 72238 983 72294 992
rect 69110 912 69166 921
rect 69110 847 69166 856
rect 69570 912 69626 921
rect 69570 847 69626 856
rect 70950 912 71006 921
rect 70950 847 71006 856
rect 72804 678 72832 1158
rect 72988 921 73016 1294
rect 73724 1057 73752 1906
rect 75736 1896 75788 1902
rect 74630 1864 74686 1873
rect 75736 1838 75788 1844
rect 74630 1799 74632 1808
rect 74684 1799 74686 1808
rect 74632 1770 74684 1776
rect 74264 1352 74316 1358
rect 74264 1294 74316 1300
rect 74724 1352 74776 1358
rect 74724 1294 74776 1300
rect 75000 1352 75052 1358
rect 75000 1294 75052 1300
rect 74080 1216 74132 1222
rect 74080 1158 74132 1164
rect 73710 1048 73766 1057
rect 73710 983 73766 992
rect 72974 912 73030 921
rect 72974 847 73030 856
rect 72792 672 72844 678
rect 72792 614 72844 620
rect 67270 504 67326 513
rect 74092 474 74120 1158
rect 74276 921 74304 1294
rect 74736 921 74764 1294
rect 75012 950 75040 1294
rect 75748 1057 75776 1838
rect 76484 1329 76512 2382
rect 78600 1970 78628 3567
rect 78680 2440 78732 2446
rect 78680 2382 78732 2388
rect 78956 2440 79008 2446
rect 78956 2382 79008 2388
rect 78588 1964 78640 1970
rect 78588 1906 78640 1912
rect 77208 1896 77260 1902
rect 77208 1838 77260 1844
rect 77484 1896 77536 1902
rect 77484 1838 77536 1844
rect 76470 1320 76526 1329
rect 76470 1255 76526 1264
rect 77220 1057 77248 1838
rect 77300 1352 77352 1358
rect 77300 1294 77352 1300
rect 75734 1048 75790 1057
rect 75734 983 75790 992
rect 77206 1048 77262 1057
rect 77206 983 77262 992
rect 75000 944 75052 950
rect 74262 912 74318 921
rect 74262 847 74318 856
rect 74722 912 74778 921
rect 77312 921 77340 1294
rect 77496 1018 77524 1838
rect 77576 1352 77628 1358
rect 78692 1329 78720 2382
rect 77576 1294 77628 1300
rect 78678 1320 78734 1329
rect 77484 1012 77536 1018
rect 77484 954 77536 960
rect 75000 886 75052 892
rect 77298 912 77354 921
rect 74722 847 74778 856
rect 77588 882 77616 1294
rect 78678 1255 78734 1264
rect 77298 847 77354 856
rect 77576 876 77628 882
rect 77576 818 77628 824
rect 78968 542 78996 2382
rect 80072 2106 80100 4383
rect 80060 2100 80112 2106
rect 80060 2042 80112 2048
rect 79416 1896 79468 1902
rect 79416 1838 79468 1844
rect 79428 1057 79456 1838
rect 79968 1352 80020 1358
rect 79968 1294 80020 1300
rect 80152 1352 80204 1358
rect 80152 1294 80204 1300
rect 79414 1048 79470 1057
rect 79414 983 79470 992
rect 79980 921 80008 1294
rect 79966 912 80022 921
rect 79966 847 80022 856
rect 80164 746 80192 1294
rect 80256 1222 80284 6258
rect 81440 4616 81492 4622
rect 81440 4558 81492 4564
rect 81164 2372 81216 2378
rect 81164 2314 81216 2320
rect 81176 1970 81204 2314
rect 81164 1964 81216 1970
rect 81164 1906 81216 1912
rect 80888 1896 80940 1902
rect 80888 1838 80940 1844
rect 80244 1216 80296 1222
rect 80244 1158 80296 1164
rect 80900 1057 80928 1838
rect 81452 1766 81480 4558
rect 84106 3360 84162 3369
rect 84106 3295 84162 3304
rect 84120 2514 84148 3295
rect 84108 2508 84160 2514
rect 84108 2450 84160 2456
rect 81624 2440 81676 2446
rect 81624 2382 81676 2388
rect 83832 2440 83884 2446
rect 83832 2382 83884 2388
rect 81440 1760 81492 1766
rect 81440 1702 81492 1708
rect 81636 1329 81664 2382
rect 82360 1896 82412 1902
rect 82360 1838 82412 1844
rect 82636 1896 82688 1902
rect 82636 1838 82688 1844
rect 81622 1320 81678 1329
rect 81622 1255 81678 1264
rect 82372 1057 82400 1838
rect 82648 1494 82676 1838
rect 82636 1488 82688 1494
rect 82636 1430 82688 1436
rect 82636 1352 82688 1358
rect 82636 1294 82688 1300
rect 82728 1352 82780 1358
rect 83844 1329 83872 2382
rect 82728 1294 82780 1300
rect 83830 1320 83886 1329
rect 80886 1048 80942 1057
rect 80886 983 80942 992
rect 82358 1048 82414 1057
rect 82358 983 82414 992
rect 82648 921 82676 1294
rect 82634 912 82690 921
rect 82634 847 82690 856
rect 80152 740 80204 746
rect 80152 682 80204 688
rect 82740 610 82768 1294
rect 84212 1290 84240 7346
rect 86960 4820 87012 4826
rect 86960 4762 87012 4768
rect 86972 2774 87000 4762
rect 88352 4690 88380 9318
rect 88812 8498 88840 9318
rect 88800 8492 88852 8498
rect 88800 8434 88852 8440
rect 88524 7948 88576 7954
rect 88524 7890 88576 7896
rect 88536 7546 88564 7890
rect 88524 7540 88576 7546
rect 88524 7482 88576 7488
rect 88340 4684 88392 4690
rect 88340 4626 88392 4632
rect 86880 2746 87000 2774
rect 84936 2644 84988 2650
rect 84936 2586 84988 2592
rect 84948 2446 84976 2586
rect 84936 2440 84988 2446
rect 84936 2382 84988 2388
rect 84842 2000 84898 2009
rect 86880 1970 86908 2746
rect 88996 2553 89024 9454
rect 89350 9415 89352 9424
rect 89404 9415 89406 9424
rect 89352 9386 89404 9392
rect 89456 8974 89484 9522
rect 90100 9178 90128 9522
rect 90376 9450 90404 10231
rect 90364 9444 90416 9450
rect 90364 9386 90416 9392
rect 90088 9172 90140 9178
rect 90088 9114 90140 9120
rect 90548 9172 90600 9178
rect 90548 9114 90600 9120
rect 89536 9036 89588 9042
rect 89536 8978 89588 8984
rect 89076 8968 89128 8974
rect 89076 8910 89128 8916
rect 89444 8968 89496 8974
rect 89444 8910 89496 8916
rect 89088 2774 89116 8910
rect 89548 8838 89576 8978
rect 89904 8968 89956 8974
rect 89904 8910 89956 8916
rect 89996 8968 90048 8974
rect 89996 8910 90048 8916
rect 89536 8832 89588 8838
rect 89536 8774 89588 8780
rect 89628 8560 89680 8566
rect 89628 8502 89680 8508
rect 89352 3052 89404 3058
rect 89352 2994 89404 3000
rect 89088 2746 89208 2774
rect 88982 2544 89038 2553
rect 88982 2479 89038 2488
rect 88996 2446 89024 2479
rect 88524 2440 88576 2446
rect 88524 2382 88576 2388
rect 88984 2440 89036 2446
rect 88984 2382 89036 2388
rect 89076 2440 89128 2446
rect 89076 2382 89128 2388
rect 88536 2310 88564 2382
rect 88524 2304 88576 2310
rect 88524 2246 88576 2252
rect 88800 2304 88852 2310
rect 88800 2246 88852 2252
rect 84842 1935 84844 1944
rect 84896 1935 84898 1944
rect 86868 1964 86920 1970
rect 84844 1906 84896 1912
rect 86868 1906 86920 1912
rect 88248 1964 88300 1970
rect 88248 1906 88300 1912
rect 84568 1896 84620 1902
rect 84568 1838 84620 1844
rect 86040 1896 86092 1902
rect 86040 1838 86092 1844
rect 83830 1255 83886 1264
rect 84200 1284 84252 1290
rect 84200 1226 84252 1232
rect 84580 1057 84608 1838
rect 85028 1352 85080 1358
rect 85028 1294 85080 1300
rect 85488 1352 85540 1358
rect 85488 1294 85540 1300
rect 84566 1048 84622 1057
rect 84566 983 84622 992
rect 82728 604 82780 610
rect 82728 546 82780 552
rect 78956 536 79008 542
rect 78956 478 79008 484
rect 67270 439 67326 448
rect 74080 468 74132 474
rect 74080 410 74132 416
rect 85040 377 85068 1294
rect 85500 377 85528 1294
rect 86052 1057 86080 1838
rect 86776 1352 86828 1358
rect 86776 1294 86828 1300
rect 86038 1048 86094 1057
rect 86038 983 86094 992
rect 86788 921 86816 1294
rect 87512 1216 87564 1222
rect 87512 1158 87564 1164
rect 88260 1170 88288 1906
rect 88524 1896 88576 1902
rect 88524 1838 88576 1844
rect 88340 1760 88392 1766
rect 88340 1702 88392 1708
rect 88352 1465 88380 1702
rect 88338 1456 88394 1465
rect 88338 1391 88394 1400
rect 88432 1216 88484 1222
rect 88260 1164 88432 1170
rect 88536 1193 88564 1838
rect 88812 1358 88840 2246
rect 89088 1970 89116 2382
rect 89076 1964 89128 1970
rect 89076 1906 89128 1912
rect 89074 1456 89130 1465
rect 89180 1442 89208 2746
rect 89364 2106 89392 2994
rect 89536 2848 89588 2854
rect 89536 2790 89588 2796
rect 89352 2100 89404 2106
rect 89352 2042 89404 2048
rect 89130 1414 89208 1442
rect 89074 1391 89076 1400
rect 89128 1391 89130 1400
rect 89076 1362 89128 1368
rect 88800 1352 88852 1358
rect 89548 1329 89576 2790
rect 89640 2145 89668 8502
rect 89718 8120 89774 8129
rect 89718 8055 89774 8064
rect 89732 7750 89760 8055
rect 89720 7744 89772 7750
rect 89720 7686 89772 7692
rect 89720 4004 89772 4010
rect 89720 3946 89772 3952
rect 89626 2136 89682 2145
rect 89626 2071 89682 2080
rect 89640 1902 89668 2071
rect 89628 1896 89680 1902
rect 89628 1838 89680 1844
rect 89732 1426 89760 3946
rect 89916 2038 89944 8910
rect 90008 8498 90036 8910
rect 90560 8838 90588 9114
rect 90744 8974 90772 10338
rect 91008 10124 91060 10130
rect 91008 10066 91060 10072
rect 90732 8968 90784 8974
rect 90732 8910 90784 8916
rect 90548 8832 90600 8838
rect 90548 8774 90600 8780
rect 90640 8832 90692 8838
rect 90640 8774 90692 8780
rect 90652 8498 90680 8774
rect 89996 8492 90048 8498
rect 89996 8434 90048 8440
rect 90640 8492 90692 8498
rect 90640 8434 90692 8440
rect 90088 8288 90140 8294
rect 90088 8230 90140 8236
rect 90100 7886 90128 8230
rect 90088 7880 90140 7886
rect 90088 7822 90140 7828
rect 90744 2774 90772 8910
rect 90822 8664 90878 8673
rect 90822 8599 90824 8608
rect 90876 8599 90878 8608
rect 90824 8570 90876 8576
rect 91020 8498 91048 10066
rect 91650 10024 91706 10033
rect 91650 9959 91706 9968
rect 91664 9586 91692 9959
rect 91560 9580 91612 9586
rect 91560 9522 91612 9528
rect 91652 9580 91704 9586
rect 91652 9522 91704 9528
rect 91100 8900 91152 8906
rect 91100 8842 91152 8848
rect 91008 8492 91060 8498
rect 91008 8434 91060 8440
rect 90916 3052 90968 3058
rect 90916 2994 90968 3000
rect 90824 2848 90876 2854
rect 90824 2790 90876 2796
rect 90560 2746 90772 2774
rect 90272 2440 90324 2446
rect 90272 2382 90324 2388
rect 90180 2304 90232 2310
rect 90180 2246 90232 2252
rect 89904 2032 89956 2038
rect 89904 1974 89956 1980
rect 89916 1902 89944 1974
rect 89904 1896 89956 1902
rect 89904 1838 89956 1844
rect 89916 1766 89944 1838
rect 89904 1760 89956 1766
rect 89904 1702 89956 1708
rect 89720 1420 89772 1426
rect 89720 1362 89772 1368
rect 90192 1329 90220 2246
rect 90284 2106 90312 2382
rect 90272 2100 90324 2106
rect 90272 2042 90324 2048
rect 90560 1426 90588 2746
rect 90732 1896 90784 1902
rect 90732 1838 90784 1844
rect 90548 1420 90600 1426
rect 90548 1362 90600 1368
rect 90744 1358 90772 1838
rect 90732 1352 90784 1358
rect 88800 1294 88852 1300
rect 89534 1320 89590 1329
rect 89534 1255 89590 1264
rect 90178 1320 90234 1329
rect 90836 1329 90864 2790
rect 90928 1358 90956 2994
rect 91020 2038 91048 8434
rect 91112 6254 91140 8842
rect 91572 8634 91600 9522
rect 92018 9480 92074 9489
rect 92018 9415 92020 9424
rect 92072 9415 92074 9424
rect 92020 9386 92072 9392
rect 91742 9208 91798 9217
rect 91652 9172 91704 9178
rect 91742 9143 91744 9152
rect 91652 9114 91704 9120
rect 91796 9143 91798 9152
rect 91744 9114 91796 9120
rect 91664 8974 91692 9114
rect 92400 8974 92428 10678
rect 93308 10396 93360 10402
rect 93308 10338 93360 10344
rect 92848 10328 92900 10334
rect 92848 10270 92900 10276
rect 92940 10328 92992 10334
rect 92940 10270 92992 10276
rect 92754 9752 92810 9761
rect 92754 9687 92756 9696
rect 92808 9687 92810 9696
rect 92756 9658 92808 9664
rect 92572 9580 92624 9586
rect 92572 9522 92624 9528
rect 91652 8968 91704 8974
rect 91652 8910 91704 8916
rect 92388 8968 92440 8974
rect 92388 8910 92440 8916
rect 91560 8628 91612 8634
rect 91560 8570 91612 8576
rect 91100 6248 91152 6254
rect 91100 6190 91152 6196
rect 91192 3120 91244 3126
rect 91192 3062 91244 3068
rect 91100 2440 91152 2446
rect 91204 2417 91232 3062
rect 91100 2382 91152 2388
rect 91190 2408 91246 2417
rect 91112 2106 91140 2382
rect 91190 2343 91246 2352
rect 91192 2304 91244 2310
rect 91192 2246 91244 2252
rect 91100 2100 91152 2106
rect 91100 2042 91152 2048
rect 91008 2032 91060 2038
rect 91008 1974 91060 1980
rect 91204 1601 91232 2246
rect 91664 1970 91692 8910
rect 92584 8634 92612 9522
rect 92860 8974 92888 10270
rect 92952 10198 92980 10270
rect 92940 10192 92992 10198
rect 92940 10134 92992 10140
rect 93032 10192 93084 10198
rect 93032 10134 93084 10140
rect 92848 8968 92900 8974
rect 92848 8910 92900 8916
rect 92940 8900 92992 8906
rect 92940 8842 92992 8848
rect 92572 8628 92624 8634
rect 92572 8570 92624 8576
rect 92952 8430 92980 8842
rect 93044 8430 93072 10134
rect 93124 8900 93176 8906
rect 93124 8842 93176 8848
rect 92940 8424 92992 8430
rect 92940 8366 92992 8372
rect 93032 8424 93084 8430
rect 93032 8366 93084 8372
rect 92572 7948 92624 7954
rect 92572 7890 92624 7896
rect 91928 7880 91980 7886
rect 91928 7822 91980 7828
rect 91940 3534 91968 7822
rect 92478 7032 92534 7041
rect 92478 6967 92534 6976
rect 92204 6112 92256 6118
rect 92204 6054 92256 6060
rect 92216 4758 92244 6054
rect 92388 5636 92440 5642
rect 92388 5578 92440 5584
rect 92400 5234 92428 5578
rect 92388 5228 92440 5234
rect 92388 5170 92440 5176
rect 92296 5024 92348 5030
rect 92296 4966 92348 4972
rect 92204 4752 92256 4758
rect 92204 4694 92256 4700
rect 92308 4690 92336 4966
rect 92296 4684 92348 4690
rect 92296 4626 92348 4632
rect 92388 4480 92440 4486
rect 92388 4422 92440 4428
rect 92204 3664 92256 3670
rect 92204 3606 92256 3612
rect 91928 3528 91980 3534
rect 91928 3470 91980 3476
rect 91836 3052 91888 3058
rect 91836 2994 91888 3000
rect 91848 2106 91876 2994
rect 92020 2848 92072 2854
rect 92020 2790 92072 2796
rect 91836 2100 91888 2106
rect 91836 2042 91888 2048
rect 91652 1964 91704 1970
rect 91652 1906 91704 1912
rect 91376 1760 91428 1766
rect 91376 1702 91428 1708
rect 91652 1760 91704 1766
rect 91652 1702 91704 1708
rect 91388 1601 91416 1702
rect 91190 1592 91246 1601
rect 91190 1527 91246 1536
rect 91374 1592 91430 1601
rect 91374 1527 91430 1536
rect 91664 1358 91692 1702
rect 90916 1352 90968 1358
rect 90732 1294 90784 1300
rect 90822 1320 90878 1329
rect 90178 1255 90234 1264
rect 90916 1294 90968 1300
rect 91652 1352 91704 1358
rect 92032 1329 92060 2790
rect 92216 2446 92244 3606
rect 92204 2440 92256 2446
rect 92204 2382 92256 2388
rect 92296 2372 92348 2378
rect 92296 2314 92348 2320
rect 91652 1294 91704 1300
rect 92018 1320 92074 1329
rect 90822 1255 90878 1264
rect 92018 1255 92074 1264
rect 88260 1158 88484 1164
rect 88522 1184 88578 1193
rect 86774 912 86830 921
rect 86774 847 86830 856
rect 87524 513 87552 1158
rect 88260 1142 88472 1158
rect 88522 1119 88578 1128
rect 92202 640 92258 649
rect 92202 575 92258 584
rect 87510 504 87566 513
rect 87510 439 87566 448
rect 40040 342 40092 348
rect 53102 368 53158 377
rect 38842 303 38898 312
rect 53102 303 53158 312
rect 63866 368 63922 377
rect 63866 303 63922 312
rect 64602 368 64658 377
rect 64602 303 64658 312
rect 65982 368 66038 377
rect 65982 303 66038 312
rect 85026 368 85082 377
rect 85026 303 85082 312
rect 85486 368 85542 377
rect 85486 303 85542 312
rect 28816 128 28868 134
rect 28816 70 28868 76
rect 29000 128 29052 134
rect 92216 105 92244 575
rect 92308 406 92336 2314
rect 92400 1902 92428 4422
rect 92492 3738 92520 6967
rect 92584 4146 92612 7890
rect 92940 6316 92992 6322
rect 92768 6276 92940 6304
rect 92664 6248 92716 6254
rect 92664 6190 92716 6196
rect 92676 5846 92704 6190
rect 92664 5840 92716 5846
rect 92664 5782 92716 5788
rect 92768 4622 92796 6276
rect 92940 6258 92992 6264
rect 92756 4616 92808 4622
rect 92756 4558 92808 4564
rect 92662 4312 92718 4321
rect 92662 4247 92718 4256
rect 92572 4140 92624 4146
rect 92572 4082 92624 4088
rect 92570 3768 92626 3777
rect 92480 3732 92532 3738
rect 92570 3703 92572 3712
rect 92480 3674 92532 3680
rect 92624 3703 92626 3712
rect 92572 3674 92624 3680
rect 92676 3466 92704 4247
rect 92768 4185 92796 4558
rect 93044 4486 93072 8366
rect 93032 4480 93084 4486
rect 93032 4422 93084 4428
rect 92754 4176 92810 4185
rect 92754 4111 92810 4120
rect 92940 4140 92992 4146
rect 92940 4082 92992 4088
rect 92952 4049 92980 4082
rect 92938 4040 92994 4049
rect 92938 3975 92994 3984
rect 92664 3460 92716 3466
rect 92664 3402 92716 3408
rect 93032 3188 93084 3194
rect 93032 3130 93084 3136
rect 92756 2848 92808 2854
rect 92756 2790 92808 2796
rect 92572 2372 92624 2378
rect 92572 2314 92624 2320
rect 92584 1970 92612 2314
rect 92572 1964 92624 1970
rect 92572 1906 92624 1912
rect 92388 1896 92440 1902
rect 92388 1838 92440 1844
rect 92400 1737 92428 1838
rect 92386 1728 92442 1737
rect 92386 1663 92442 1672
rect 92388 1488 92440 1494
rect 92388 1430 92440 1436
rect 92400 921 92428 1430
rect 92768 1329 92796 2790
rect 92848 2440 92900 2446
rect 92848 2382 92900 2388
rect 92860 1562 92888 2382
rect 92940 1760 92992 1766
rect 92940 1702 92992 1708
rect 92848 1556 92900 1562
rect 92848 1498 92900 1504
rect 92754 1320 92810 1329
rect 92754 1255 92810 1264
rect 92480 1216 92532 1222
rect 92480 1158 92532 1164
rect 92572 1216 92624 1222
rect 92572 1158 92624 1164
rect 92386 912 92442 921
rect 92386 847 92442 856
rect 92492 649 92520 1158
rect 92584 882 92612 1158
rect 92572 876 92624 882
rect 92572 818 92624 824
rect 92952 678 92980 1702
rect 93044 1057 93072 3130
rect 93136 1970 93164 8842
rect 93216 8288 93268 8294
rect 93216 8230 93268 8236
rect 93228 4010 93256 8230
rect 93320 5030 93348 10338
rect 93490 9752 93546 9761
rect 93490 9687 93492 9696
rect 93544 9687 93546 9696
rect 93492 9658 93544 9664
rect 93676 9580 93728 9586
rect 93676 9522 93728 9528
rect 93688 9178 93716 9522
rect 93676 9172 93728 9178
rect 93676 9114 93728 9120
rect 93400 8968 93452 8974
rect 93400 8910 93452 8916
rect 93492 8968 93544 8974
rect 93492 8910 93544 8916
rect 93412 7154 93440 8910
rect 93504 8498 93532 8910
rect 93492 8492 93544 8498
rect 93492 8434 93544 8440
rect 93964 7342 93992 10746
rect 94608 9722 94636 10814
rect 94596 9716 94648 9722
rect 94596 9658 94648 9664
rect 94228 9172 94280 9178
rect 94228 9114 94280 9120
rect 94044 9104 94096 9110
rect 94044 9046 94096 9052
rect 93952 7336 94004 7342
rect 93952 7278 94004 7284
rect 93860 7268 93912 7274
rect 93860 7210 93912 7216
rect 93412 7126 93532 7154
rect 93308 5024 93360 5030
rect 93308 4966 93360 4972
rect 93504 4554 93532 7126
rect 93584 6996 93636 7002
rect 93584 6938 93636 6944
rect 93492 4548 93544 4554
rect 93492 4490 93544 4496
rect 93216 4004 93268 4010
rect 93216 3946 93268 3952
rect 93308 3936 93360 3942
rect 93308 3878 93360 3884
rect 93216 3528 93268 3534
rect 93216 3470 93268 3476
rect 93228 2106 93256 3470
rect 93320 3194 93348 3878
rect 93308 3188 93360 3194
rect 93308 3130 93360 3136
rect 93504 3074 93532 4490
rect 93596 4146 93624 6938
rect 93768 6724 93820 6730
rect 93768 6666 93820 6672
rect 93780 5930 93808 6666
rect 93872 6118 93900 7210
rect 93952 6452 94004 6458
rect 93952 6394 94004 6400
rect 93860 6112 93912 6118
rect 93860 6054 93912 6060
rect 93780 5902 93900 5930
rect 93584 4140 93636 4146
rect 93584 4082 93636 4088
rect 93320 3046 93532 3074
rect 93216 2100 93268 2106
rect 93216 2042 93268 2048
rect 93320 1986 93348 3046
rect 93400 2984 93452 2990
rect 93400 2926 93452 2932
rect 93124 1964 93176 1970
rect 93124 1906 93176 1912
rect 93228 1958 93348 1986
rect 93228 1358 93256 1958
rect 93412 1358 93440 2926
rect 93872 2514 93900 5902
rect 93964 3534 93992 6394
rect 94056 5846 94084 9046
rect 94240 6905 94268 9114
rect 94608 9042 94636 9658
rect 94792 9586 94820 10814
rect 99196 10804 99248 10810
rect 99196 10746 99248 10752
rect 94964 10668 95016 10674
rect 94964 10610 95016 10616
rect 94780 9580 94832 9586
rect 94780 9522 94832 9528
rect 94872 9580 94924 9586
rect 94872 9522 94924 9528
rect 94596 9036 94648 9042
rect 94516 8996 94596 9024
rect 94412 8832 94464 8838
rect 94412 8774 94464 8780
rect 94424 8498 94452 8774
rect 94412 8492 94464 8498
rect 94412 8434 94464 8440
rect 94318 8120 94374 8129
rect 94318 8055 94374 8064
rect 94332 7721 94360 8055
rect 94318 7712 94374 7721
rect 94516 7698 94544 8996
rect 94596 8978 94648 8984
rect 94884 8974 94912 9522
rect 94872 8968 94924 8974
rect 94872 8910 94924 8916
rect 94872 8832 94924 8838
rect 94872 8774 94924 8780
rect 94594 8664 94650 8673
rect 94594 8599 94596 8608
rect 94648 8599 94650 8608
rect 94596 8570 94648 8576
rect 94884 8498 94912 8774
rect 94872 8492 94924 8498
rect 94872 8434 94924 8440
rect 94318 7647 94374 7656
rect 94424 7670 94544 7698
rect 94226 6896 94282 6905
rect 94226 6831 94282 6840
rect 94228 6656 94280 6662
rect 94228 6598 94280 6604
rect 94136 6112 94188 6118
rect 94136 6054 94188 6060
rect 94044 5840 94096 5846
rect 94044 5782 94096 5788
rect 94148 3670 94176 6054
rect 94136 3664 94188 3670
rect 94136 3606 94188 3612
rect 93952 3528 94004 3534
rect 93952 3470 94004 3476
rect 94044 3528 94096 3534
rect 94044 3470 94096 3476
rect 93952 3392 94004 3398
rect 93952 3334 94004 3340
rect 93964 3097 93992 3334
rect 93950 3088 94006 3097
rect 93950 3023 94006 3032
rect 93860 2508 93912 2514
rect 93860 2450 93912 2456
rect 93768 2304 93820 2310
rect 93674 2272 93730 2281
rect 93768 2246 93820 2252
rect 93674 2207 93730 2216
rect 93492 1896 93544 1902
rect 93688 1873 93716 2207
rect 93780 2038 93808 2246
rect 93768 2032 93820 2038
rect 93768 1974 93820 1980
rect 93492 1838 93544 1844
rect 93674 1864 93730 1873
rect 93216 1352 93268 1358
rect 93216 1294 93268 1300
rect 93308 1352 93360 1358
rect 93308 1294 93360 1300
rect 93400 1352 93452 1358
rect 93400 1294 93452 1300
rect 93504 1340 93532 1838
rect 94056 1834 94084 3470
rect 94136 3052 94188 3058
rect 94136 2994 94188 3000
rect 94148 2106 94176 2994
rect 94240 2774 94268 6598
rect 94424 5658 94452 7670
rect 94502 7576 94558 7585
rect 94502 7511 94558 7520
rect 94516 7177 94544 7511
rect 94502 7168 94558 7177
rect 94502 7103 94558 7112
rect 94976 7018 95004 10610
rect 96436 10600 96488 10606
rect 96436 10542 96488 10548
rect 98644 10600 98696 10606
rect 98644 10542 98696 10548
rect 95516 10328 95568 10334
rect 95516 10270 95568 10276
rect 95608 10328 95660 10334
rect 95608 10270 95660 10276
rect 95528 10062 95556 10270
rect 95424 10056 95476 10062
rect 95424 9998 95476 10004
rect 95516 10056 95568 10062
rect 95516 9998 95568 10004
rect 95240 9036 95292 9042
rect 95240 8978 95292 8984
rect 95054 8664 95110 8673
rect 95054 8599 95056 8608
rect 95108 8599 95110 8608
rect 95056 8570 95108 8576
rect 95252 8537 95280 8978
rect 95436 8634 95464 9998
rect 95424 8628 95476 8634
rect 95424 8570 95476 8576
rect 95238 8528 95294 8537
rect 95056 8492 95108 8498
rect 95436 8498 95464 8570
rect 95238 8463 95294 8472
rect 95424 8492 95476 8498
rect 95056 8434 95108 8440
rect 95424 8434 95476 8440
rect 94884 6990 95004 7018
rect 94504 6792 94556 6798
rect 94504 6734 94556 6740
rect 94516 6361 94544 6734
rect 94688 6724 94740 6730
rect 94688 6666 94740 6672
rect 94502 6352 94558 6361
rect 94502 6287 94558 6296
rect 94504 5908 94556 5914
rect 94504 5850 94556 5856
rect 94516 5817 94544 5850
rect 94502 5808 94558 5817
rect 94502 5743 94558 5752
rect 94700 5710 94728 6666
rect 94780 6112 94832 6118
rect 94780 6054 94832 6060
rect 94596 5704 94648 5710
rect 94424 5630 94544 5658
rect 94596 5646 94648 5652
rect 94688 5704 94740 5710
rect 94688 5646 94740 5652
rect 94412 5568 94464 5574
rect 94410 5536 94412 5545
rect 94464 5536 94466 5545
rect 94410 5471 94466 5480
rect 94516 5114 94544 5630
rect 94320 5092 94372 5098
rect 94320 5034 94372 5040
rect 94424 5086 94544 5114
rect 94332 4622 94360 5034
rect 94320 4616 94372 4622
rect 94320 4558 94372 4564
rect 94424 4162 94452 5086
rect 94504 5024 94556 5030
rect 94504 4966 94556 4972
rect 94516 4690 94544 4966
rect 94608 4690 94636 5646
rect 94688 5024 94740 5030
rect 94688 4966 94740 4972
rect 94504 4684 94556 4690
rect 94504 4626 94556 4632
rect 94596 4684 94648 4690
rect 94596 4626 94648 4632
rect 94700 4554 94728 4966
rect 94688 4548 94740 4554
rect 94688 4490 94740 4496
rect 94596 4480 94648 4486
rect 94596 4422 94648 4428
rect 94332 4134 94452 4162
rect 94504 4208 94556 4214
rect 94504 4150 94556 4156
rect 94332 3058 94360 4134
rect 94412 4072 94464 4078
rect 94412 4014 94464 4020
rect 94320 3052 94372 3058
rect 94320 2994 94372 3000
rect 94240 2746 94360 2774
rect 94226 2136 94282 2145
rect 94136 2100 94188 2106
rect 94226 2071 94282 2080
rect 94136 2042 94188 2048
rect 94240 1970 94268 2071
rect 94228 1964 94280 1970
rect 94228 1906 94280 1912
rect 93674 1799 93730 1808
rect 94044 1828 94096 1834
rect 94044 1770 94096 1776
rect 93584 1352 93636 1358
rect 93504 1312 93584 1340
rect 93320 1170 93348 1294
rect 93504 1170 93532 1312
rect 93584 1294 93636 1300
rect 93320 1142 93532 1170
rect 93030 1048 93086 1057
rect 93030 983 93086 992
rect 92940 672 92992 678
rect 92478 640 92534 649
rect 92940 614 92992 620
rect 92478 575 92534 584
rect 92296 400 92348 406
rect 92296 342 92348 348
rect 94332 241 94360 2746
rect 94424 2689 94452 4014
rect 94516 3602 94544 4150
rect 94608 4146 94636 4422
rect 94596 4140 94648 4146
rect 94596 4082 94648 4088
rect 94792 4078 94820 6054
rect 94780 4072 94832 4078
rect 94780 4014 94832 4020
rect 94688 3664 94740 3670
rect 94688 3606 94740 3612
rect 94504 3596 94556 3602
rect 94504 3538 94556 3544
rect 94504 3052 94556 3058
rect 94504 2994 94556 3000
rect 94410 2680 94466 2689
rect 94410 2615 94466 2624
rect 94412 2440 94464 2446
rect 94412 2382 94464 2388
rect 94424 1358 94452 2382
rect 94516 1426 94544 2994
rect 94700 2774 94728 3606
rect 94884 3602 94912 6990
rect 95068 6916 95096 8434
rect 95148 8016 95200 8022
rect 95148 7958 95200 7964
rect 94976 6888 95096 6916
rect 94872 3596 94924 3602
rect 94872 3538 94924 3544
rect 94870 3224 94926 3233
rect 94870 3159 94926 3168
rect 94700 2746 94820 2774
rect 94792 2582 94820 2746
rect 94688 2576 94740 2582
rect 94688 2518 94740 2524
rect 94780 2576 94832 2582
rect 94780 2518 94832 2524
rect 94596 2508 94648 2514
rect 94596 2450 94648 2456
rect 94608 1766 94636 2450
rect 94700 2106 94728 2518
rect 94688 2100 94740 2106
rect 94688 2042 94740 2048
rect 94792 1834 94820 2518
rect 94780 1828 94832 1834
rect 94780 1770 94832 1776
rect 94596 1760 94648 1766
rect 94596 1702 94648 1708
rect 94504 1420 94556 1426
rect 94504 1362 94556 1368
rect 94412 1352 94464 1358
rect 94412 1294 94464 1300
rect 94596 1216 94648 1222
rect 94596 1158 94648 1164
rect 94608 1057 94636 1158
rect 94594 1048 94650 1057
rect 94594 983 94650 992
rect 94780 876 94832 882
rect 94780 818 94832 824
rect 94792 649 94820 818
rect 94884 678 94912 3159
rect 94976 3058 95004 6888
rect 95054 6080 95110 6089
rect 95054 6015 95110 6024
rect 95068 3602 95096 6015
rect 95160 5370 95188 7958
rect 95516 6928 95568 6934
rect 95516 6870 95568 6876
rect 95240 6860 95292 6866
rect 95240 6802 95292 6808
rect 95252 6322 95280 6802
rect 95332 6452 95384 6458
rect 95332 6394 95384 6400
rect 95240 6316 95292 6322
rect 95240 6258 95292 6264
rect 95240 5636 95292 5642
rect 95240 5578 95292 5584
rect 95148 5364 95200 5370
rect 95148 5306 95200 5312
rect 95252 5302 95280 5578
rect 95240 5296 95292 5302
rect 95240 5238 95292 5244
rect 95344 5098 95372 6394
rect 95332 5092 95384 5098
rect 95332 5034 95384 5040
rect 95332 4480 95384 4486
rect 95332 4422 95384 4428
rect 95148 4072 95200 4078
rect 95148 4014 95200 4020
rect 95056 3596 95108 3602
rect 95056 3538 95108 3544
rect 95160 3482 95188 4014
rect 95240 3936 95292 3942
rect 95240 3878 95292 3884
rect 95252 3777 95280 3878
rect 95238 3768 95294 3777
rect 95238 3703 95294 3712
rect 95068 3454 95188 3482
rect 94964 3052 95016 3058
rect 94964 2994 95016 3000
rect 95068 2938 95096 3454
rect 95238 3224 95294 3233
rect 95238 3159 95294 3168
rect 94976 2910 95096 2938
rect 94976 1426 95004 2910
rect 95252 2774 95280 3159
rect 95160 2746 95280 2774
rect 95056 1896 95108 1902
rect 95054 1864 95056 1873
rect 95108 1864 95110 1873
rect 95160 1850 95188 2746
rect 95240 2508 95292 2514
rect 95344 2496 95372 4422
rect 95528 4185 95556 6870
rect 95620 4486 95648 10270
rect 95792 10056 95844 10062
rect 95792 9998 95844 10004
rect 95700 8492 95752 8498
rect 95700 8434 95752 8440
rect 95712 8362 95740 8434
rect 95700 8356 95752 8362
rect 95700 8298 95752 8304
rect 95700 7540 95752 7546
rect 95700 7482 95752 7488
rect 95608 4480 95660 4486
rect 95608 4422 95660 4428
rect 95514 4176 95570 4185
rect 95514 4111 95570 4120
rect 95528 3602 95556 4111
rect 95516 3596 95568 3602
rect 95568 3556 95648 3584
rect 95516 3538 95568 3544
rect 95424 2916 95476 2922
rect 95424 2858 95476 2864
rect 95436 2825 95464 2858
rect 95422 2816 95478 2825
rect 95422 2751 95478 2760
rect 95292 2468 95372 2496
rect 95240 2450 95292 2456
rect 95516 2440 95568 2446
rect 95620 2428 95648 3556
rect 95712 2922 95740 7482
rect 95700 2916 95752 2922
rect 95700 2858 95752 2864
rect 95568 2400 95648 2428
rect 95516 2382 95568 2388
rect 95330 2136 95386 2145
rect 95330 2071 95386 2080
rect 95110 1822 95188 1850
rect 95238 1864 95294 1873
rect 95054 1799 95110 1808
rect 95238 1799 95294 1808
rect 94964 1420 95016 1426
rect 94964 1362 95016 1368
rect 95252 814 95280 1799
rect 95344 1601 95372 2071
rect 95330 1592 95386 1601
rect 95528 1562 95556 2382
rect 95608 1896 95660 1902
rect 95608 1838 95660 1844
rect 95330 1527 95386 1536
rect 95516 1556 95568 1562
rect 95516 1498 95568 1504
rect 95620 1358 95648 1838
rect 95804 1426 95832 9998
rect 96066 9752 96122 9761
rect 95976 9716 96028 9722
rect 96066 9687 96068 9696
rect 95976 9658 96028 9664
rect 96120 9687 96122 9696
rect 96342 9752 96398 9761
rect 96342 9687 96344 9696
rect 96068 9658 96120 9664
rect 96396 9687 96398 9696
rect 96344 9658 96396 9664
rect 95988 9042 96016 9658
rect 96160 9580 96212 9586
rect 96160 9522 96212 9528
rect 96068 9172 96120 9178
rect 96068 9114 96120 9120
rect 95976 9036 96028 9042
rect 95976 8978 96028 8984
rect 95882 8528 95938 8537
rect 95882 8463 95884 8472
rect 95936 8463 95938 8472
rect 95884 8434 95936 8440
rect 95988 8265 96016 8978
rect 96080 8838 96108 9114
rect 96068 8832 96120 8838
rect 96068 8774 96120 8780
rect 96172 8634 96200 9522
rect 96252 9172 96304 9178
rect 96252 9114 96304 9120
rect 96160 8628 96212 8634
rect 96160 8570 96212 8576
rect 95974 8256 96030 8265
rect 95974 8191 96030 8200
rect 95976 7744 96028 7750
rect 95976 7686 96028 7692
rect 95884 7540 95936 7546
rect 95884 7482 95936 7488
rect 95896 7410 95924 7482
rect 95884 7404 95936 7410
rect 95884 7346 95936 7352
rect 95988 6746 96016 7686
rect 96160 7336 96212 7342
rect 96160 7278 96212 7284
rect 96172 6934 96200 7278
rect 96160 6928 96212 6934
rect 96160 6870 96212 6876
rect 95896 6718 96016 6746
rect 96160 6792 96212 6798
rect 96160 6734 96212 6740
rect 95896 1970 95924 6718
rect 95976 6656 96028 6662
rect 95976 6598 96028 6604
rect 95988 5166 96016 6598
rect 96068 6112 96120 6118
rect 96068 6054 96120 6060
rect 96080 5914 96108 6054
rect 96172 5914 96200 6734
rect 96068 5908 96120 5914
rect 96068 5850 96120 5856
rect 96160 5908 96212 5914
rect 96160 5850 96212 5856
rect 96068 5704 96120 5710
rect 96068 5646 96120 5652
rect 96080 5545 96108 5646
rect 96160 5568 96212 5574
rect 96066 5536 96122 5545
rect 96160 5510 96212 5516
rect 96066 5471 96122 5480
rect 96172 5370 96200 5510
rect 96068 5364 96120 5370
rect 96068 5306 96120 5312
rect 96160 5364 96212 5370
rect 96160 5306 96212 5312
rect 95976 5160 96028 5166
rect 95976 5102 96028 5108
rect 95976 3664 96028 3670
rect 95976 3606 96028 3612
rect 95988 2281 96016 3606
rect 96080 2836 96108 5306
rect 96160 4548 96212 4554
rect 96160 4490 96212 4496
rect 96172 4078 96200 4490
rect 96160 4072 96212 4078
rect 96160 4014 96212 4020
rect 96172 3097 96200 4014
rect 96158 3088 96214 3097
rect 96158 3023 96214 3032
rect 96160 2984 96212 2990
rect 96264 2972 96292 9114
rect 96448 8430 96476 10542
rect 96620 10464 96672 10470
rect 96618 10432 96620 10441
rect 96672 10432 96674 10441
rect 96618 10367 96674 10376
rect 96528 10260 96580 10266
rect 96528 10202 96580 10208
rect 96540 9178 96568 10202
rect 98656 10062 98684 10542
rect 98828 10464 98880 10470
rect 98828 10406 98880 10412
rect 98552 10056 98604 10062
rect 98552 9998 98604 10004
rect 98644 10056 98696 10062
rect 98644 9998 98696 10004
rect 96896 9580 96948 9586
rect 96896 9522 96948 9528
rect 96528 9172 96580 9178
rect 96528 9114 96580 9120
rect 96528 9036 96580 9042
rect 96528 8978 96580 8984
rect 96540 8945 96568 8978
rect 96620 8968 96672 8974
rect 96526 8936 96582 8945
rect 96620 8910 96672 8916
rect 96526 8871 96582 8880
rect 96632 8430 96660 8910
rect 96908 8634 96936 9522
rect 97724 9172 97776 9178
rect 97724 9114 97776 9120
rect 96986 9072 97042 9081
rect 96986 9007 97042 9016
rect 97000 8974 97028 9007
rect 97736 8974 97764 9114
rect 98564 8974 98592 9998
rect 96988 8968 97040 8974
rect 96988 8910 97040 8916
rect 97724 8968 97776 8974
rect 97724 8910 97776 8916
rect 98092 8968 98144 8974
rect 98552 8968 98604 8974
rect 98092 8910 98144 8916
rect 98550 8936 98552 8945
rect 98604 8936 98606 8945
rect 97356 8900 97408 8906
rect 97356 8842 97408 8848
rect 97540 8900 97592 8906
rect 97540 8842 97592 8848
rect 97264 8832 97316 8838
rect 97264 8774 97316 8780
rect 97368 8786 97396 8842
rect 97552 8786 97580 8842
rect 97276 8634 97304 8774
rect 97368 8758 97580 8786
rect 96896 8628 96948 8634
rect 96896 8570 96948 8576
rect 97264 8628 97316 8634
rect 97264 8570 97316 8576
rect 97172 8560 97224 8566
rect 97170 8528 97172 8537
rect 97224 8528 97226 8537
rect 97170 8463 97226 8472
rect 97264 8492 97316 8498
rect 97460 8480 97488 8758
rect 97538 8664 97594 8673
rect 97538 8599 97540 8608
rect 97592 8599 97594 8608
rect 97998 8664 98054 8673
rect 97998 8599 98000 8608
rect 97540 8570 97592 8576
rect 98052 8599 98054 8608
rect 98000 8570 98052 8576
rect 98104 8498 98132 8910
rect 98550 8871 98606 8880
rect 97316 8452 97488 8480
rect 98092 8492 98144 8498
rect 97264 8434 97316 8440
rect 98092 8434 98144 8440
rect 96436 8424 96488 8430
rect 96356 8384 96436 8412
rect 96356 4146 96384 8384
rect 96436 8366 96488 8372
rect 96620 8424 96672 8430
rect 96620 8366 96672 8372
rect 98000 8424 98052 8430
rect 98000 8366 98052 8372
rect 96620 7948 96672 7954
rect 96620 7890 96672 7896
rect 96632 7857 96660 7890
rect 96618 7848 96674 7857
rect 96618 7783 96674 7792
rect 98012 7750 98040 8366
rect 98000 7744 98052 7750
rect 98000 7686 98052 7692
rect 97264 7472 97316 7478
rect 97264 7414 97316 7420
rect 96528 7336 96580 7342
rect 96528 7278 96580 7284
rect 96540 7002 96568 7278
rect 97080 7200 97132 7206
rect 97080 7142 97132 7148
rect 96528 6996 96580 7002
rect 96528 6938 96580 6944
rect 96988 6860 97040 6866
rect 96988 6802 97040 6808
rect 96712 6656 96764 6662
rect 96712 6598 96764 6604
rect 96724 6390 96752 6598
rect 96712 6384 96764 6390
rect 96712 6326 96764 6332
rect 96804 6384 96856 6390
rect 96804 6326 96856 6332
rect 96436 5908 96488 5914
rect 96436 5850 96488 5856
rect 96448 5692 96476 5850
rect 96620 5840 96672 5846
rect 96816 5794 96844 6326
rect 96896 6248 96948 6254
rect 96896 6190 96948 6196
rect 96672 5788 96844 5794
rect 96620 5782 96844 5788
rect 96632 5766 96844 5782
rect 96804 5704 96856 5710
rect 96448 5664 96568 5692
rect 96540 5624 96568 5664
rect 96804 5646 96856 5652
rect 96908 5658 96936 6190
rect 97000 5778 97028 6802
rect 97092 5778 97120 7142
rect 97172 6928 97224 6934
rect 97172 6870 97224 6876
rect 96988 5772 97040 5778
rect 96988 5714 97040 5720
rect 97080 5772 97132 5778
rect 97080 5714 97132 5720
rect 96540 5596 96660 5624
rect 96436 5568 96488 5574
rect 96436 5510 96488 5516
rect 96448 5370 96476 5510
rect 96632 5370 96660 5596
rect 96436 5364 96488 5370
rect 96436 5306 96488 5312
rect 96620 5364 96672 5370
rect 96620 5306 96672 5312
rect 96620 5160 96672 5166
rect 96620 5102 96672 5108
rect 96632 5001 96660 5102
rect 96618 4992 96674 5001
rect 96618 4927 96674 4936
rect 96436 4616 96488 4622
rect 96436 4558 96488 4564
rect 96344 4140 96396 4146
rect 96344 4082 96396 4088
rect 96448 3194 96476 4558
rect 96526 4448 96582 4457
rect 96526 4383 96582 4392
rect 96540 3194 96568 4383
rect 96712 4004 96764 4010
rect 96712 3946 96764 3952
rect 96618 3904 96674 3913
rect 96618 3839 96674 3848
rect 96436 3188 96488 3194
rect 96436 3130 96488 3136
rect 96528 3188 96580 3194
rect 96528 3130 96580 3136
rect 96632 3058 96660 3839
rect 96344 3052 96396 3058
rect 96344 2994 96396 3000
rect 96620 3052 96672 3058
rect 96620 2994 96672 3000
rect 96212 2944 96292 2972
rect 96160 2926 96212 2932
rect 96080 2808 96200 2836
rect 96068 2372 96120 2378
rect 96068 2314 96120 2320
rect 95974 2272 96030 2281
rect 95974 2207 96030 2216
rect 96080 2106 96108 2314
rect 96068 2100 96120 2106
rect 96068 2042 96120 2048
rect 95884 1964 95936 1970
rect 95884 1906 95936 1912
rect 95792 1420 95844 1426
rect 95792 1362 95844 1368
rect 95608 1352 95660 1358
rect 95608 1294 95660 1300
rect 96172 814 96200 2808
rect 96252 2304 96304 2310
rect 96252 2246 96304 2252
rect 96264 1601 96292 2246
rect 96356 1970 96384 2994
rect 96436 2916 96488 2922
rect 96488 2876 96568 2904
rect 96436 2858 96488 2864
rect 96434 2408 96490 2417
rect 96434 2343 96490 2352
rect 96448 2310 96476 2343
rect 96436 2304 96488 2310
rect 96436 2246 96488 2252
rect 96434 2136 96490 2145
rect 96434 2071 96436 2080
rect 96488 2071 96490 2080
rect 96436 2042 96488 2048
rect 96344 1964 96396 1970
rect 96344 1906 96396 1912
rect 96250 1592 96306 1601
rect 96250 1527 96306 1536
rect 96540 1358 96568 2876
rect 96724 2514 96752 3946
rect 96816 3618 96844 5646
rect 96908 5630 97028 5658
rect 97000 5556 97028 5630
rect 96908 5528 97028 5556
rect 96908 5098 96936 5528
rect 96988 5364 97040 5370
rect 96988 5306 97040 5312
rect 96896 5092 96948 5098
rect 96896 5034 96948 5040
rect 96896 4072 96948 4078
rect 96896 4014 96948 4020
rect 96908 3738 96936 4014
rect 97000 3738 97028 5306
rect 97184 4554 97212 6870
rect 97172 4548 97224 4554
rect 97172 4490 97224 4496
rect 96896 3732 96948 3738
rect 96896 3674 96948 3680
rect 96988 3732 97040 3738
rect 96988 3674 97040 3680
rect 96816 3590 96936 3618
rect 96908 3534 96936 3590
rect 96804 3528 96856 3534
rect 96804 3470 96856 3476
rect 96896 3528 96948 3534
rect 96896 3470 96948 3476
rect 96712 2508 96764 2514
rect 96712 2450 96764 2456
rect 96816 1737 96844 3470
rect 97276 3194 97304 7414
rect 97356 7404 97408 7410
rect 97356 7346 97408 7352
rect 97540 7404 97592 7410
rect 97540 7346 97592 7352
rect 98736 7404 98788 7410
rect 98736 7346 98788 7352
rect 97368 6798 97396 7346
rect 97448 7200 97500 7206
rect 97448 7142 97500 7148
rect 97460 6905 97488 7142
rect 97446 6896 97502 6905
rect 97552 6866 97580 7346
rect 98552 7336 98604 7342
rect 98552 7278 98604 7284
rect 97724 7200 97776 7206
rect 97724 7142 97776 7148
rect 97816 7200 97868 7206
rect 97816 7142 97868 7148
rect 97446 6831 97502 6840
rect 97540 6860 97592 6866
rect 97356 6792 97408 6798
rect 97356 6734 97408 6740
rect 97356 6248 97408 6254
rect 97356 6190 97408 6196
rect 97368 5710 97396 6190
rect 97460 6118 97488 6831
rect 97540 6802 97592 6808
rect 97448 6112 97500 6118
rect 97448 6054 97500 6060
rect 97356 5704 97408 5710
rect 97356 5646 97408 5652
rect 97368 3534 97396 5646
rect 97448 5568 97500 5574
rect 97448 5510 97500 5516
rect 97460 5166 97488 5510
rect 97552 5409 97580 6802
rect 97736 6458 97764 7142
rect 97724 6452 97776 6458
rect 97724 6394 97776 6400
rect 97724 6112 97776 6118
rect 97724 6054 97776 6060
rect 97632 5840 97684 5846
rect 97632 5782 97684 5788
rect 97538 5400 97594 5409
rect 97538 5335 97594 5344
rect 97448 5160 97500 5166
rect 97448 5102 97500 5108
rect 97540 4480 97592 4486
rect 97540 4422 97592 4428
rect 97552 3777 97580 4422
rect 97644 4049 97672 5782
rect 97736 5778 97764 6054
rect 97724 5772 97776 5778
rect 97724 5714 97776 5720
rect 97724 5160 97776 5166
rect 97724 5102 97776 5108
rect 97630 4040 97686 4049
rect 97630 3975 97686 3984
rect 97538 3768 97594 3777
rect 97538 3703 97594 3712
rect 97736 3670 97764 5102
rect 97828 4010 97856 7142
rect 98000 6996 98052 7002
rect 98000 6938 98052 6944
rect 97908 6928 97960 6934
rect 97906 6896 97908 6905
rect 97960 6896 97962 6905
rect 97906 6831 97962 6840
rect 97908 6316 97960 6322
rect 97908 6258 97960 6264
rect 97920 5846 97948 6258
rect 98012 6118 98040 6938
rect 98276 6792 98328 6798
rect 98276 6734 98328 6740
rect 98460 6792 98512 6798
rect 98460 6734 98512 6740
rect 98092 6724 98144 6730
rect 98092 6666 98144 6672
rect 98000 6112 98052 6118
rect 98000 6054 98052 6060
rect 97908 5840 97960 5846
rect 97908 5782 97960 5788
rect 98012 5370 98040 6054
rect 98104 5370 98132 6666
rect 98288 6322 98316 6734
rect 98368 6452 98420 6458
rect 98368 6394 98420 6400
rect 98276 6316 98328 6322
rect 98276 6258 98328 6264
rect 98000 5364 98052 5370
rect 98000 5306 98052 5312
rect 98092 5364 98144 5370
rect 98092 5306 98144 5312
rect 98380 4690 98408 6394
rect 98472 6254 98500 6734
rect 98564 6390 98592 7278
rect 98644 6656 98696 6662
rect 98644 6598 98696 6604
rect 98552 6384 98604 6390
rect 98552 6326 98604 6332
rect 98460 6248 98512 6254
rect 98512 6208 98592 6236
rect 98460 6190 98512 6196
rect 98564 5778 98592 6208
rect 98460 5772 98512 5778
rect 98460 5714 98512 5720
rect 98552 5772 98604 5778
rect 98552 5714 98604 5720
rect 98472 5409 98500 5714
rect 98656 5642 98684 6598
rect 98748 6458 98776 7346
rect 98736 6452 98788 6458
rect 98736 6394 98788 6400
rect 98644 5636 98696 5642
rect 98644 5578 98696 5584
rect 98458 5400 98514 5409
rect 98458 5335 98514 5344
rect 98472 5234 98500 5335
rect 98460 5228 98512 5234
rect 98460 5170 98512 5176
rect 98840 5166 98868 10406
rect 98920 9580 98972 9586
rect 98920 9522 98972 9528
rect 98932 9178 98960 9522
rect 98920 9172 98972 9178
rect 98920 9114 98972 9120
rect 99208 9042 99236 10746
rect 100024 10600 100076 10606
rect 100024 10542 100076 10548
rect 99378 9752 99434 9761
rect 99378 9687 99380 9696
rect 99432 9687 99434 9696
rect 99380 9658 99432 9664
rect 99286 9072 99342 9081
rect 99196 9036 99248 9042
rect 99286 9007 99288 9016
rect 99196 8978 99248 8984
rect 99340 9007 99342 9016
rect 99288 8978 99340 8984
rect 99470 8936 99526 8945
rect 99470 8871 99526 8880
rect 99378 8664 99434 8673
rect 99378 8599 99380 8608
rect 99432 8599 99434 8608
rect 99380 8570 99432 8576
rect 99484 8566 99512 8871
rect 99656 8832 99708 8838
rect 99656 8774 99708 8780
rect 99472 8560 99524 8566
rect 98918 8528 98974 8537
rect 99472 8502 99524 8508
rect 99668 8498 99696 8774
rect 98918 8463 98974 8472
rect 99656 8492 99708 8498
rect 98828 5160 98880 5166
rect 98828 5102 98880 5108
rect 98368 4684 98420 4690
rect 98368 4626 98420 4632
rect 98644 4684 98696 4690
rect 98644 4626 98696 4632
rect 98656 4214 98684 4626
rect 98644 4208 98696 4214
rect 98644 4150 98696 4156
rect 98276 4072 98328 4078
rect 98276 4014 98328 4020
rect 97816 4004 97868 4010
rect 97816 3946 97868 3952
rect 97724 3664 97776 3670
rect 97724 3606 97776 3612
rect 97356 3528 97408 3534
rect 97356 3470 97408 3476
rect 97264 3188 97316 3194
rect 97264 3130 97316 3136
rect 97632 3188 97684 3194
rect 97632 3130 97684 3136
rect 97908 3188 97960 3194
rect 97908 3130 97960 3136
rect 96988 2848 97040 2854
rect 96986 2816 96988 2825
rect 97356 2848 97408 2854
rect 97040 2816 97042 2825
rect 97356 2790 97408 2796
rect 96986 2751 97042 2760
rect 96894 2408 96950 2417
rect 96894 2343 96950 2352
rect 96908 1970 96936 2343
rect 96896 1964 96948 1970
rect 96896 1906 96948 1912
rect 97080 1896 97132 1902
rect 97080 1838 97132 1844
rect 96802 1728 96858 1737
rect 96802 1663 96858 1672
rect 96986 1728 97042 1737
rect 96986 1663 97042 1672
rect 97000 1562 97028 1663
rect 96988 1556 97040 1562
rect 96988 1498 97040 1504
rect 96528 1352 96580 1358
rect 96528 1294 96580 1300
rect 95240 808 95292 814
rect 95240 750 95292 756
rect 96160 808 96212 814
rect 96160 750 96212 756
rect 94872 672 94924 678
rect 94778 640 94834 649
rect 94872 614 94924 620
rect 94778 575 94834 584
rect 97092 474 97120 1838
rect 97368 1222 97396 2790
rect 97644 2582 97672 3130
rect 97722 2680 97778 2689
rect 97722 2615 97778 2624
rect 97736 2582 97764 2615
rect 97632 2576 97684 2582
rect 97632 2518 97684 2524
rect 97724 2576 97776 2582
rect 97724 2518 97776 2524
rect 97920 2378 97948 3130
rect 97908 2372 97960 2378
rect 97908 2314 97960 2320
rect 97814 2136 97870 2145
rect 97814 2071 97870 2080
rect 97908 2100 97960 2106
rect 97828 1970 97856 2071
rect 97908 2042 97960 2048
rect 97828 1964 97886 1970
rect 97828 1924 97834 1964
rect 97834 1906 97886 1912
rect 97448 1828 97500 1834
rect 97448 1770 97500 1776
rect 97460 1494 97488 1770
rect 97920 1601 97948 2042
rect 98092 1964 98144 1970
rect 98012 1924 98092 1952
rect 98012 1737 98040 1924
rect 98092 1906 98144 1912
rect 97998 1728 98054 1737
rect 97998 1663 98054 1672
rect 97906 1592 97962 1601
rect 97906 1527 97962 1536
rect 97448 1488 97500 1494
rect 97448 1430 97500 1436
rect 97816 1352 97868 1358
rect 97816 1294 97868 1300
rect 97908 1352 97960 1358
rect 98012 1340 98040 1663
rect 97960 1312 98040 1340
rect 97908 1294 97960 1300
rect 97356 1216 97408 1222
rect 97356 1158 97408 1164
rect 97828 882 97856 1294
rect 97816 876 97868 882
rect 97816 818 97868 824
rect 97080 468 97132 474
rect 97080 410 97132 416
rect 94318 232 94374 241
rect 94318 167 94374 176
rect 98288 105 98316 4014
rect 98460 3392 98512 3398
rect 98460 3334 98512 3340
rect 98472 1426 98500 3334
rect 98736 2440 98788 2446
rect 98736 2382 98788 2388
rect 98748 2106 98776 2382
rect 98828 2304 98880 2310
rect 98828 2246 98880 2252
rect 98840 2106 98868 2246
rect 98736 2100 98788 2106
rect 98736 2042 98788 2048
rect 98828 2100 98880 2106
rect 98828 2042 98880 2048
rect 98932 1426 98960 8463
rect 99656 8434 99708 8440
rect 99102 8392 99158 8401
rect 99102 8327 99158 8336
rect 99012 7336 99064 7342
rect 99012 7278 99064 7284
rect 99024 5574 99052 7278
rect 99116 7274 99144 8327
rect 99288 7880 99340 7886
rect 99288 7822 99340 7828
rect 99300 7478 99328 7822
rect 99196 7472 99248 7478
rect 99196 7414 99248 7420
rect 99288 7472 99340 7478
rect 99288 7414 99340 7420
rect 99208 7290 99236 7414
rect 99208 7274 99512 7290
rect 99104 7268 99156 7274
rect 99208 7268 99524 7274
rect 99208 7262 99472 7268
rect 99104 7210 99156 7216
rect 99472 7210 99524 7216
rect 99288 7200 99340 7206
rect 99288 7142 99340 7148
rect 99932 7200 99984 7206
rect 99932 7142 99984 7148
rect 99196 6860 99248 6866
rect 99196 6802 99248 6808
rect 99102 6488 99158 6497
rect 99102 6423 99158 6432
rect 99012 5568 99064 5574
rect 99012 5510 99064 5516
rect 99012 2984 99064 2990
rect 99012 2926 99064 2932
rect 99024 2378 99052 2926
rect 99012 2372 99064 2378
rect 99012 2314 99064 2320
rect 99116 2310 99144 6423
rect 99208 5030 99236 6802
rect 99196 5024 99248 5030
rect 99196 4966 99248 4972
rect 99196 4208 99248 4214
rect 99196 4150 99248 4156
rect 99104 2304 99156 2310
rect 99104 2246 99156 2252
rect 98460 1420 98512 1426
rect 98460 1362 98512 1368
rect 98920 1420 98972 1426
rect 98920 1362 98972 1368
rect 98736 1352 98788 1358
rect 99208 1329 99236 4150
rect 99300 3602 99328 7142
rect 99380 6792 99432 6798
rect 99380 6734 99432 6740
rect 99840 6792 99892 6798
rect 99840 6734 99892 6740
rect 99392 6254 99420 6734
rect 99852 6662 99880 6734
rect 99656 6656 99708 6662
rect 99656 6598 99708 6604
rect 99840 6656 99892 6662
rect 99840 6598 99892 6604
rect 99564 6316 99616 6322
rect 99564 6258 99616 6264
rect 99380 6248 99432 6254
rect 99380 6190 99432 6196
rect 99472 6112 99524 6118
rect 99472 6054 99524 6060
rect 99380 5704 99432 5710
rect 99380 5646 99432 5652
rect 99392 5234 99420 5646
rect 99484 5284 99512 6054
rect 99576 5710 99604 6258
rect 99564 5704 99616 5710
rect 99564 5646 99616 5652
rect 99564 5296 99616 5302
rect 99484 5256 99564 5284
rect 99564 5238 99616 5244
rect 99380 5228 99432 5234
rect 99380 5170 99432 5176
rect 99392 4622 99420 5170
rect 99564 5160 99616 5166
rect 99564 5102 99616 5108
rect 99470 4856 99526 4865
rect 99470 4791 99472 4800
rect 99524 4791 99526 4800
rect 99472 4762 99524 4768
rect 99380 4616 99432 4622
rect 99380 4558 99432 4564
rect 99576 4554 99604 5102
rect 99564 4548 99616 4554
rect 99564 4490 99616 4496
rect 99288 3596 99340 3602
rect 99288 3538 99340 3544
rect 99380 3460 99432 3466
rect 99380 3402 99432 3408
rect 99392 2922 99420 3402
rect 99380 2916 99432 2922
rect 99380 2858 99432 2864
rect 99288 1896 99340 1902
rect 99288 1838 99340 1844
rect 99300 1562 99328 1838
rect 99288 1556 99340 1562
rect 99288 1498 99340 1504
rect 99392 1358 99420 2858
rect 99668 2514 99696 6598
rect 99748 6112 99800 6118
rect 99748 6054 99800 6060
rect 99760 3126 99788 6054
rect 99840 5092 99892 5098
rect 99840 5034 99892 5040
rect 99852 4457 99880 5034
rect 99838 4448 99894 4457
rect 99838 4383 99894 4392
rect 99748 3120 99800 3126
rect 99748 3062 99800 3068
rect 99656 2508 99708 2514
rect 99656 2450 99708 2456
rect 99944 2038 99972 7142
rect 100036 6866 100064 10542
rect 100482 9752 100538 9761
rect 100482 9687 100484 9696
rect 100536 9687 100538 9696
rect 100668 9716 100720 9722
rect 100484 9658 100536 9664
rect 100668 9658 100720 9664
rect 100208 9580 100260 9586
rect 100208 9522 100260 9528
rect 100576 9580 100628 9586
rect 100576 9522 100628 9528
rect 100220 8838 100248 9522
rect 100588 9178 100616 9522
rect 100576 9172 100628 9178
rect 100576 9114 100628 9120
rect 100300 8968 100352 8974
rect 100300 8910 100352 8916
rect 100208 8832 100260 8838
rect 100208 8774 100260 8780
rect 100312 8566 100340 8910
rect 100300 8560 100352 8566
rect 100298 8528 100300 8537
rect 100352 8528 100354 8537
rect 100298 8463 100354 8472
rect 100680 8401 100708 9658
rect 100772 8430 100800 10814
rect 132776 10804 132828 10810
rect 132776 10746 132828 10752
rect 133788 10804 133840 10810
rect 133788 10746 133840 10752
rect 146576 10804 146628 10810
rect 146576 10746 146628 10752
rect 125876 10736 125928 10742
rect 125876 10678 125928 10684
rect 106188 10668 106240 10674
rect 106188 10610 106240 10616
rect 105452 10396 105504 10402
rect 105452 10338 105504 10344
rect 103242 10296 103298 10305
rect 103242 10231 103298 10240
rect 103886 10296 103942 10305
rect 103886 10231 103942 10240
rect 104714 10296 104770 10305
rect 104714 10231 104770 10240
rect 103060 9648 103112 9654
rect 103060 9590 103112 9596
rect 100852 9580 100904 9586
rect 100852 9522 100904 9528
rect 100760 8424 100812 8430
rect 100666 8392 100722 8401
rect 100760 8366 100812 8372
rect 100666 8327 100722 8336
rect 100484 8084 100536 8090
rect 100484 8026 100536 8032
rect 100024 6860 100076 6866
rect 100024 6802 100076 6808
rect 100496 6497 100524 8026
rect 100668 8016 100720 8022
rect 100668 7958 100720 7964
rect 100576 7540 100628 7546
rect 100576 7482 100628 7488
rect 100588 7206 100616 7482
rect 100576 7200 100628 7206
rect 100576 7142 100628 7148
rect 100680 7041 100708 7958
rect 100772 7546 100800 8366
rect 100760 7540 100812 7546
rect 100760 7482 100812 7488
rect 100666 7032 100722 7041
rect 100666 6967 100722 6976
rect 100482 6488 100538 6497
rect 100482 6423 100538 6432
rect 100392 6316 100444 6322
rect 100392 6258 100444 6264
rect 100668 6316 100720 6322
rect 100668 6258 100720 6264
rect 100206 6216 100262 6225
rect 100206 6151 100262 6160
rect 100116 5908 100168 5914
rect 100116 5850 100168 5856
rect 100128 5574 100156 5850
rect 100024 5568 100076 5574
rect 100024 5510 100076 5516
rect 100116 5568 100168 5574
rect 100116 5510 100168 5516
rect 100036 5370 100064 5510
rect 100024 5364 100076 5370
rect 100024 5306 100076 5312
rect 100024 5092 100076 5098
rect 100024 5034 100076 5040
rect 100036 4865 100064 5034
rect 100128 5030 100156 5510
rect 100116 5024 100168 5030
rect 100116 4966 100168 4972
rect 100022 4856 100078 4865
rect 100128 4826 100156 4966
rect 100022 4791 100078 4800
rect 100116 4820 100168 4826
rect 100116 4762 100168 4768
rect 100022 4584 100078 4593
rect 100022 4519 100078 4528
rect 100036 2514 100064 4519
rect 100220 3942 100248 6151
rect 100404 5710 100432 6258
rect 100392 5704 100444 5710
rect 100298 5672 100354 5681
rect 100392 5646 100444 5652
rect 100298 5607 100300 5616
rect 100352 5607 100354 5616
rect 100300 5578 100352 5584
rect 100312 5234 100340 5578
rect 100404 5522 100432 5646
rect 100680 5642 100708 6258
rect 100864 6066 100892 9522
rect 101496 9512 101548 9518
rect 101496 9454 101548 9460
rect 101218 9208 101274 9217
rect 101218 9143 101220 9152
rect 101272 9143 101274 9152
rect 101220 9114 101272 9120
rect 101508 8974 101536 9454
rect 102345 9276 102653 9285
rect 102345 9274 102351 9276
rect 102407 9274 102431 9276
rect 102487 9274 102511 9276
rect 102567 9274 102591 9276
rect 102647 9274 102653 9276
rect 102407 9222 102409 9274
rect 102589 9222 102591 9274
rect 102345 9220 102351 9222
rect 102407 9220 102431 9222
rect 102487 9220 102511 9222
rect 102567 9220 102591 9222
rect 102647 9220 102653 9222
rect 102345 9211 102653 9220
rect 100944 8968 100996 8974
rect 100944 8910 100996 8916
rect 101036 8968 101088 8974
rect 101036 8910 101088 8916
rect 101496 8968 101548 8974
rect 101496 8910 101548 8916
rect 100956 8430 100984 8910
rect 100944 8424 100996 8430
rect 100944 8366 100996 8372
rect 100956 7886 100984 8366
rect 101048 8090 101076 8910
rect 102048 8492 102100 8498
rect 102048 8434 102100 8440
rect 101956 8424 102008 8430
rect 101956 8366 102008 8372
rect 101036 8084 101088 8090
rect 101036 8026 101088 8032
rect 101496 8016 101548 8022
rect 101496 7958 101548 7964
rect 100944 7880 100996 7886
rect 100944 7822 100996 7828
rect 101508 7410 101536 7958
rect 101968 7954 101996 8366
rect 102060 8265 102088 8434
rect 102046 8256 102102 8265
rect 102046 8191 102102 8200
rect 102345 8188 102653 8197
rect 102345 8186 102351 8188
rect 102407 8186 102431 8188
rect 102487 8186 102511 8188
rect 102567 8186 102591 8188
rect 102647 8186 102653 8188
rect 102407 8134 102409 8186
rect 102589 8134 102591 8186
rect 102345 8132 102351 8134
rect 102407 8132 102431 8134
rect 102487 8132 102511 8134
rect 102567 8132 102591 8134
rect 102647 8132 102653 8134
rect 102345 8123 102653 8132
rect 101956 7948 102008 7954
rect 101956 7890 102008 7896
rect 102874 7712 102930 7721
rect 102874 7647 102930 7656
rect 101404 7404 101456 7410
rect 101404 7346 101456 7352
rect 101496 7404 101548 7410
rect 101496 7346 101548 7352
rect 100944 6996 100996 7002
rect 100944 6938 100996 6944
rect 100956 6118 100984 6938
rect 101220 6724 101272 6730
rect 101220 6666 101272 6672
rect 101128 6656 101180 6662
rect 101128 6598 101180 6604
rect 101036 6452 101088 6458
rect 101036 6394 101088 6400
rect 101048 6322 101076 6394
rect 101036 6316 101088 6322
rect 101036 6258 101088 6264
rect 100772 6038 100892 6066
rect 100944 6112 100996 6118
rect 100944 6054 100996 6060
rect 100668 5636 100720 5642
rect 100668 5578 100720 5584
rect 100404 5494 100616 5522
rect 100392 5296 100444 5302
rect 100392 5238 100444 5244
rect 100300 5228 100352 5234
rect 100300 5170 100352 5176
rect 100312 4622 100340 5170
rect 100404 5030 100432 5238
rect 100588 5166 100616 5494
rect 100576 5160 100628 5166
rect 100576 5102 100628 5108
rect 100392 5024 100444 5030
rect 100392 4966 100444 4972
rect 100404 4826 100432 4966
rect 100392 4820 100444 4826
rect 100392 4762 100444 4768
rect 100300 4616 100352 4622
rect 100300 4558 100352 4564
rect 100588 4554 100616 5102
rect 100666 4720 100722 4729
rect 100666 4655 100722 4664
rect 100576 4548 100628 4554
rect 100576 4490 100628 4496
rect 100680 4282 100708 4655
rect 100668 4276 100720 4282
rect 100668 4218 100720 4224
rect 100298 4040 100354 4049
rect 100298 3975 100354 3984
rect 100208 3936 100260 3942
rect 100208 3878 100260 3884
rect 100312 3505 100340 3975
rect 100772 3754 100800 6038
rect 100850 5944 100906 5953
rect 100956 5914 100984 6054
rect 100850 5879 100906 5888
rect 100944 5908 100996 5914
rect 100864 4690 100892 5879
rect 100944 5850 100996 5856
rect 100944 5704 100996 5710
rect 101048 5692 101076 6258
rect 100996 5664 101076 5692
rect 100944 5646 100996 5652
rect 100852 4684 100904 4690
rect 100852 4626 100904 4632
rect 100772 3726 100892 3754
rect 100760 3664 100812 3670
rect 100760 3606 100812 3612
rect 100298 3496 100354 3505
rect 100298 3431 100354 3440
rect 100482 3496 100538 3505
rect 100482 3431 100538 3440
rect 100496 3233 100524 3431
rect 100772 3233 100800 3606
rect 100482 3224 100538 3233
rect 100482 3159 100538 3168
rect 100758 3224 100814 3233
rect 100758 3159 100814 3168
rect 100864 2774 100892 3726
rect 100944 3460 100996 3466
rect 100944 3402 100996 3408
rect 100772 2746 100892 2774
rect 100024 2508 100076 2514
rect 100024 2450 100076 2456
rect 100484 2372 100536 2378
rect 100484 2314 100536 2320
rect 99932 2032 99984 2038
rect 99932 1974 99984 1980
rect 99380 1352 99432 1358
rect 98736 1294 98788 1300
rect 99194 1320 99250 1329
rect 98748 814 98776 1294
rect 99380 1294 99432 1300
rect 99840 1352 99892 1358
rect 99840 1294 99892 1300
rect 99194 1255 99250 1264
rect 99288 1216 99340 1222
rect 99288 1158 99340 1164
rect 98736 808 98788 814
rect 98736 750 98788 756
rect 98828 808 98880 814
rect 98828 750 98880 756
rect 98840 406 98868 750
rect 99300 649 99328 1158
rect 99852 950 99880 1294
rect 99840 944 99892 950
rect 99840 886 99892 892
rect 99286 640 99342 649
rect 99286 575 99342 584
rect 98828 400 98880 406
rect 98828 342 98880 348
rect 100496 270 100524 2314
rect 100576 1420 100628 1426
rect 100772 1408 100800 2746
rect 100956 2446 100984 3402
rect 101034 3224 101090 3233
rect 101034 3159 101090 3168
rect 100944 2440 100996 2446
rect 100944 2382 100996 2388
rect 101048 2038 101076 3159
rect 101036 2032 101088 2038
rect 101036 1974 101088 1980
rect 101140 1902 101168 6598
rect 101232 4826 101260 6666
rect 101310 6216 101366 6225
rect 101310 6151 101366 6160
rect 101324 5681 101352 6151
rect 101310 5672 101366 5681
rect 101310 5607 101366 5616
rect 101324 5234 101352 5607
rect 101416 5370 101444 7346
rect 102138 7168 102194 7177
rect 102138 7103 102194 7112
rect 102152 6984 102180 7103
rect 102345 7100 102653 7109
rect 102345 7098 102351 7100
rect 102407 7098 102431 7100
rect 102487 7098 102511 7100
rect 102567 7098 102591 7100
rect 102647 7098 102653 7100
rect 102407 7046 102409 7098
rect 102589 7046 102591 7098
rect 102345 7044 102351 7046
rect 102407 7044 102431 7046
rect 102487 7044 102511 7046
rect 102567 7044 102591 7046
rect 102647 7044 102653 7046
rect 102345 7035 102653 7044
rect 102152 6956 102824 6984
rect 102232 6860 102284 6866
rect 102232 6802 102284 6808
rect 101680 6792 101732 6798
rect 101680 6734 101732 6740
rect 101770 6760 101826 6769
rect 101588 6656 101640 6662
rect 101588 6598 101640 6604
rect 101496 6316 101548 6322
rect 101496 6258 101548 6264
rect 101508 5953 101536 6258
rect 101494 5944 101550 5953
rect 101494 5879 101550 5888
rect 101508 5778 101536 5879
rect 101496 5772 101548 5778
rect 101496 5714 101548 5720
rect 101404 5364 101456 5370
rect 101404 5306 101456 5312
rect 101312 5228 101364 5234
rect 101312 5170 101364 5176
rect 101404 5024 101456 5030
rect 101404 4966 101456 4972
rect 101220 4820 101272 4826
rect 101220 4762 101272 4768
rect 101416 4486 101444 4966
rect 101404 4480 101456 4486
rect 101404 4422 101456 4428
rect 101508 4298 101536 5714
rect 101416 4270 101536 4298
rect 101220 4072 101272 4078
rect 101220 4014 101272 4020
rect 101232 3233 101260 4014
rect 101416 3602 101444 4270
rect 101496 4208 101548 4214
rect 101496 4150 101548 4156
rect 101404 3596 101456 3602
rect 101404 3538 101456 3544
rect 101218 3224 101274 3233
rect 101218 3159 101274 3168
rect 101508 2990 101536 4150
rect 101600 3126 101628 6598
rect 101692 6186 101720 6734
rect 102244 6746 102272 6802
rect 102692 6792 102744 6798
rect 101770 6695 101826 6704
rect 101968 6718 102272 6746
rect 102690 6760 102692 6769
rect 102744 6760 102746 6769
rect 102324 6724 102376 6730
rect 101680 6180 101732 6186
rect 101680 6122 101732 6128
rect 101784 6066 101812 6695
rect 101864 6452 101916 6458
rect 101864 6394 101916 6400
rect 101876 6322 101904 6394
rect 101864 6316 101916 6322
rect 101864 6258 101916 6264
rect 101692 6038 101812 6066
rect 101864 6112 101916 6118
rect 101968 6089 101996 6718
rect 102690 6695 102746 6704
rect 102324 6666 102376 6672
rect 102140 6656 102192 6662
rect 102140 6598 102192 6604
rect 102048 6316 102100 6322
rect 102048 6258 102100 6264
rect 101864 6054 101916 6060
rect 101954 6080 102010 6089
rect 101692 5846 101720 6038
rect 101772 5908 101824 5914
rect 101876 5896 101904 6054
rect 101954 6015 102010 6024
rect 102060 5953 102088 6258
rect 101824 5868 101904 5896
rect 102046 5944 102102 5953
rect 102046 5879 102102 5888
rect 101772 5850 101824 5856
rect 101680 5840 101732 5846
rect 101680 5782 101732 5788
rect 101678 5672 101734 5681
rect 101678 5607 101734 5616
rect 101692 5234 101720 5607
rect 101680 5228 101732 5234
rect 101680 5170 101732 5176
rect 101784 5030 101812 5850
rect 101956 5636 102008 5642
rect 101956 5578 102008 5584
rect 101864 5228 101916 5234
rect 101864 5170 101916 5176
rect 101772 5024 101824 5030
rect 101772 4966 101824 4972
rect 101784 3738 101812 4966
rect 101772 3732 101824 3738
rect 101772 3674 101824 3680
rect 101876 3534 101904 5170
rect 101968 3738 101996 5578
rect 102046 4312 102102 4321
rect 102046 4247 102102 4256
rect 102060 4146 102088 4247
rect 102048 4140 102100 4146
rect 102048 4082 102100 4088
rect 101956 3732 102008 3738
rect 101956 3674 102008 3680
rect 101864 3528 101916 3534
rect 101864 3470 101916 3476
rect 101588 3120 101640 3126
rect 101588 3062 101640 3068
rect 101496 2984 101548 2990
rect 101496 2926 101548 2932
rect 102152 2514 102180 6598
rect 102336 6458 102364 6666
rect 102324 6452 102376 6458
rect 102324 6394 102376 6400
rect 102345 6012 102653 6021
rect 102345 6010 102351 6012
rect 102407 6010 102431 6012
rect 102487 6010 102511 6012
rect 102567 6010 102591 6012
rect 102647 6010 102653 6012
rect 102407 5958 102409 6010
rect 102589 5958 102591 6010
rect 102345 5956 102351 5958
rect 102407 5956 102431 5958
rect 102487 5956 102511 5958
rect 102567 5956 102591 5958
rect 102647 5956 102653 5958
rect 102345 5947 102653 5956
rect 102416 5772 102468 5778
rect 102416 5714 102468 5720
rect 102324 5704 102376 5710
rect 102324 5646 102376 5652
rect 102336 5234 102364 5646
rect 102324 5228 102376 5234
rect 102324 5170 102376 5176
rect 102428 5166 102456 5714
rect 102416 5160 102468 5166
rect 102416 5102 102468 5108
rect 102345 4924 102653 4933
rect 102345 4922 102351 4924
rect 102407 4922 102431 4924
rect 102487 4922 102511 4924
rect 102567 4922 102591 4924
rect 102647 4922 102653 4924
rect 102407 4870 102409 4922
rect 102589 4870 102591 4922
rect 102345 4868 102351 4870
rect 102407 4868 102431 4870
rect 102487 4868 102511 4870
rect 102567 4868 102591 4870
rect 102647 4868 102653 4870
rect 102345 4859 102653 4868
rect 102796 4826 102824 6956
rect 102784 4820 102836 4826
rect 102784 4762 102836 4768
rect 102230 4176 102286 4185
rect 102230 4111 102286 4120
rect 102244 3534 102272 4111
rect 102888 4010 102916 7647
rect 102968 5840 103020 5846
rect 102968 5782 103020 5788
rect 102980 5710 103008 5782
rect 102968 5704 103020 5710
rect 102968 5646 103020 5652
rect 102968 5568 103020 5574
rect 102968 5510 103020 5516
rect 102980 4078 103008 5510
rect 102968 4072 103020 4078
rect 102968 4014 103020 4020
rect 102876 4004 102928 4010
rect 102876 3946 102928 3952
rect 102345 3836 102653 3845
rect 102345 3834 102351 3836
rect 102407 3834 102431 3836
rect 102487 3834 102511 3836
rect 102567 3834 102591 3836
rect 102647 3834 102653 3836
rect 102407 3782 102409 3834
rect 102589 3782 102591 3834
rect 102345 3780 102351 3782
rect 102407 3780 102431 3782
rect 102487 3780 102511 3782
rect 102567 3780 102591 3782
rect 102647 3780 102653 3782
rect 102345 3771 102653 3780
rect 102232 3528 102284 3534
rect 102232 3470 102284 3476
rect 103072 3398 103100 9590
rect 103256 9586 103284 10231
rect 103900 9586 103928 10231
rect 104728 9586 104756 10231
rect 105464 9722 105492 10338
rect 105634 10296 105690 10305
rect 105634 10231 105690 10240
rect 105452 9716 105504 9722
rect 105452 9658 105504 9664
rect 105648 9586 105676 10231
rect 106200 9722 106228 10610
rect 124220 10532 124272 10538
rect 124220 10474 124272 10480
rect 124680 10532 124732 10538
rect 124680 10474 124732 10480
rect 122840 10464 122892 10470
rect 122840 10406 122892 10412
rect 107016 10328 107068 10334
rect 106278 10296 106334 10305
rect 107016 10270 107068 10276
rect 107198 10296 107254 10305
rect 106278 10231 106334 10240
rect 106188 9716 106240 9722
rect 106188 9658 106240 9664
rect 106292 9586 106320 10231
rect 103244 9580 103296 9586
rect 103244 9522 103296 9528
rect 103888 9580 103940 9586
rect 103888 9522 103940 9528
rect 104716 9580 104768 9586
rect 104716 9522 104768 9528
rect 105636 9580 105688 9586
rect 105636 9522 105688 9528
rect 106280 9580 106332 9586
rect 106280 9522 106332 9528
rect 103428 9376 103480 9382
rect 103428 9318 103480 9324
rect 103704 9376 103756 9382
rect 103704 9318 103756 9324
rect 104072 9376 104124 9382
rect 104072 9318 104124 9324
rect 103440 8265 103468 9318
rect 103716 9110 103744 9318
rect 103704 9104 103756 9110
rect 103704 9046 103756 9052
rect 103426 8256 103482 8265
rect 103426 8191 103482 8200
rect 103428 7200 103480 7206
rect 103428 7142 103480 7148
rect 103888 7200 103940 7206
rect 103888 7142 103940 7148
rect 103336 6656 103388 6662
rect 103336 6598 103388 6604
rect 103152 5024 103204 5030
rect 103152 4966 103204 4972
rect 103244 5024 103296 5030
rect 103244 4966 103296 4972
rect 103164 4690 103192 4966
rect 103152 4684 103204 4690
rect 103152 4626 103204 4632
rect 103150 3496 103206 3505
rect 103150 3431 103152 3440
rect 103204 3431 103206 3440
rect 103152 3402 103204 3408
rect 103060 3392 103112 3398
rect 103060 3334 103112 3340
rect 102345 2748 102653 2757
rect 102345 2746 102351 2748
rect 102407 2746 102431 2748
rect 102487 2746 102511 2748
rect 102567 2746 102591 2748
rect 102647 2746 102653 2748
rect 102407 2694 102409 2746
rect 102589 2694 102591 2746
rect 102345 2692 102351 2694
rect 102407 2692 102431 2694
rect 102487 2692 102511 2694
rect 102567 2692 102591 2694
rect 102647 2692 102653 2694
rect 102345 2683 102653 2692
rect 102140 2508 102192 2514
rect 102140 2450 102192 2456
rect 101312 2440 101364 2446
rect 101310 2408 101312 2417
rect 101364 2408 101366 2417
rect 101310 2343 101366 2352
rect 101496 2372 101548 2378
rect 101496 2314 101548 2320
rect 101128 1896 101180 1902
rect 101128 1838 101180 1844
rect 100850 1728 100906 1737
rect 100850 1663 100906 1672
rect 100628 1380 100800 1408
rect 100576 1362 100628 1368
rect 100864 1358 100892 1663
rect 101508 1358 101536 2314
rect 103256 1834 103284 4966
rect 103244 1828 103296 1834
rect 103244 1770 103296 1776
rect 101680 1760 101732 1766
rect 101680 1702 101732 1708
rect 101692 1358 101720 1702
rect 102345 1660 102653 1669
rect 102345 1658 102351 1660
rect 102407 1658 102431 1660
rect 102487 1658 102511 1660
rect 102567 1658 102591 1660
rect 102647 1658 102653 1660
rect 102407 1606 102409 1658
rect 102589 1606 102591 1658
rect 102345 1604 102351 1606
rect 102407 1604 102431 1606
rect 102487 1604 102511 1606
rect 102567 1604 102591 1606
rect 102647 1604 102653 1606
rect 102345 1595 102653 1604
rect 100852 1352 100904 1358
rect 100852 1294 100904 1300
rect 101496 1352 101548 1358
rect 101496 1294 101548 1300
rect 101680 1352 101732 1358
rect 101680 1294 101732 1300
rect 100760 1216 100812 1222
rect 100760 1158 100812 1164
rect 100772 921 100800 1158
rect 100864 950 100892 1294
rect 100852 944 100904 950
rect 100758 912 100814 921
rect 100852 886 100904 892
rect 103348 882 103376 6598
rect 103440 5914 103468 7142
rect 103610 6624 103666 6633
rect 103610 6559 103666 6568
rect 103520 6112 103572 6118
rect 103520 6054 103572 6060
rect 103428 5908 103480 5914
rect 103428 5850 103480 5856
rect 103426 4040 103482 4049
rect 103532 4026 103560 6054
rect 103482 3998 103560 4026
rect 103426 3975 103482 3984
rect 103624 3058 103652 6559
rect 103796 6112 103848 6118
rect 103796 6054 103848 6060
rect 103808 4758 103836 6054
rect 103796 4752 103848 4758
rect 103796 4694 103848 4700
rect 103702 3632 103758 3641
rect 103702 3567 103704 3576
rect 103756 3567 103758 3576
rect 103704 3538 103756 3544
rect 103704 3392 103756 3398
rect 103704 3334 103756 3340
rect 103716 3126 103744 3334
rect 103704 3120 103756 3126
rect 103704 3062 103756 3068
rect 103612 3052 103664 3058
rect 103612 2994 103664 3000
rect 103900 1358 103928 7142
rect 103980 4820 104032 4826
rect 103980 4762 104032 4768
rect 103888 1352 103940 1358
rect 103888 1294 103940 1300
rect 103520 1216 103572 1222
rect 103520 1158 103572 1164
rect 103796 1216 103848 1222
rect 103796 1158 103848 1164
rect 103532 950 103560 1158
rect 103808 1018 103836 1158
rect 103992 1018 104020 4762
rect 104084 2145 104112 9318
rect 107028 9178 107056 10270
rect 107198 10231 107254 10240
rect 107750 10296 107806 10305
rect 107750 10231 107806 10240
rect 108394 10296 108450 10305
rect 108394 10231 108450 10240
rect 109038 10296 109094 10305
rect 109038 10231 109094 10240
rect 110050 10296 110106 10305
rect 110050 10231 110106 10240
rect 110786 10296 110842 10305
rect 110786 10231 110842 10240
rect 111522 10296 111578 10305
rect 111522 10231 111578 10240
rect 112350 10296 112406 10305
rect 112350 10231 112406 10240
rect 112902 10296 112958 10305
rect 112902 10231 112958 10240
rect 113546 10296 113602 10305
rect 113546 10231 113602 10240
rect 114190 10296 114246 10305
rect 114190 10231 114246 10240
rect 115202 10296 115258 10305
rect 115202 10231 115258 10240
rect 115754 10296 115810 10305
rect 115754 10231 115810 10240
rect 116674 10296 116730 10305
rect 116674 10231 116730 10240
rect 117226 10296 117282 10305
rect 117226 10231 117282 10240
rect 118054 10296 118110 10305
rect 118054 10231 118110 10240
rect 118698 10296 118754 10305
rect 118698 10231 118754 10240
rect 119342 10296 119398 10305
rect 119342 10231 119398 10240
rect 120354 10296 120410 10305
rect 120354 10231 120410 10240
rect 121090 10296 121146 10305
rect 121090 10231 121146 10240
rect 121734 10296 121790 10305
rect 121734 10231 121790 10240
rect 122378 10296 122434 10305
rect 122378 10231 122434 10240
rect 107016 9172 107068 9178
rect 107016 9114 107068 9120
rect 104992 9104 105044 9110
rect 104992 9046 105044 9052
rect 104440 7948 104492 7954
rect 104440 7890 104492 7896
rect 104164 7812 104216 7818
rect 104164 7754 104216 7760
rect 104176 7478 104204 7754
rect 104164 7472 104216 7478
rect 104164 7414 104216 7420
rect 104346 4992 104402 5001
rect 104346 4927 104402 4936
rect 104360 4486 104388 4927
rect 104348 4480 104400 4486
rect 104348 4422 104400 4428
rect 104360 3942 104388 4422
rect 104164 3936 104216 3942
rect 104164 3878 104216 3884
rect 104348 3936 104400 3942
rect 104452 3924 104480 7890
rect 104624 6316 104676 6322
rect 104624 6258 104676 6264
rect 104532 6180 104584 6186
rect 104532 6122 104584 6128
rect 104544 5846 104572 6122
rect 104532 5840 104584 5846
rect 104532 5782 104584 5788
rect 104532 5704 104584 5710
rect 104532 5646 104584 5652
rect 104544 4049 104572 5646
rect 104530 4040 104586 4049
rect 104530 3975 104586 3984
rect 104452 3896 104572 3924
rect 104636 3913 104664 6258
rect 104900 5840 104952 5846
rect 104900 5782 104952 5788
rect 104808 5568 104860 5574
rect 104808 5510 104860 5516
rect 104716 4480 104768 4486
rect 104716 4422 104768 4428
rect 104348 3878 104400 3884
rect 104176 3670 104204 3878
rect 104438 3768 104494 3777
rect 104438 3703 104494 3712
rect 104544 3720 104572 3896
rect 104622 3904 104678 3913
rect 104622 3839 104678 3848
rect 104164 3664 104216 3670
rect 104164 3606 104216 3612
rect 104070 2136 104126 2145
rect 104070 2071 104126 2080
rect 104176 1834 104204 3606
rect 104452 3602 104480 3703
rect 104544 3692 104597 3720
rect 104569 3602 104597 3692
rect 104440 3596 104492 3602
rect 104440 3538 104492 3544
rect 104557 3596 104609 3602
rect 104557 3538 104609 3544
rect 104728 2854 104756 4422
rect 104348 2848 104400 2854
rect 104254 2816 104310 2825
rect 104348 2790 104400 2796
rect 104716 2848 104768 2854
rect 104716 2790 104768 2796
rect 104254 2751 104310 2760
rect 104268 2650 104296 2751
rect 104360 2650 104388 2790
rect 104256 2644 104308 2650
rect 104256 2586 104308 2592
rect 104348 2644 104400 2650
rect 104348 2586 104400 2592
rect 104820 2514 104848 5510
rect 104912 4622 104940 5782
rect 104900 4616 104952 4622
rect 104900 4558 104952 4564
rect 104898 3904 104954 3913
rect 104898 3839 104954 3848
rect 104912 3233 104940 3839
rect 105004 3777 105032 9046
rect 107212 8974 107240 10231
rect 107764 9586 107792 10231
rect 108120 9716 108172 9722
rect 108120 9658 108172 9664
rect 107752 9580 107804 9586
rect 107752 9522 107804 9528
rect 108132 9450 108160 9658
rect 108408 9586 108436 10231
rect 109052 9586 109080 10231
rect 110064 9586 110092 10231
rect 110512 9988 110564 9994
rect 110512 9930 110564 9936
rect 108396 9580 108448 9586
rect 108396 9522 108448 9528
rect 109040 9580 109092 9586
rect 109040 9522 109092 9528
rect 110052 9580 110104 9586
rect 110052 9522 110104 9528
rect 108120 9444 108172 9450
rect 108120 9386 108172 9392
rect 109040 9444 109092 9450
rect 109040 9386 109092 9392
rect 109684 9444 109736 9450
rect 109684 9386 109736 9392
rect 108948 9376 109000 9382
rect 108948 9318 109000 9324
rect 108960 9110 108988 9318
rect 108948 9104 109000 9110
rect 108948 9046 109000 9052
rect 106372 8968 106424 8974
rect 106372 8910 106424 8916
rect 107200 8968 107252 8974
rect 107200 8910 107252 8916
rect 105084 8900 105136 8906
rect 105084 8842 105136 8848
rect 104990 3768 105046 3777
rect 104990 3703 105046 3712
rect 105096 3482 105124 8842
rect 106278 8256 106334 8265
rect 106278 8191 106334 8200
rect 106292 6866 106320 8191
rect 106384 7002 106412 8910
rect 107752 7880 107804 7886
rect 107752 7822 107804 7828
rect 107108 7404 107160 7410
rect 107108 7346 107160 7352
rect 106372 6996 106424 7002
rect 106372 6938 106424 6944
rect 106280 6860 106332 6866
rect 106280 6802 106332 6808
rect 106188 6792 106240 6798
rect 106188 6734 106240 6740
rect 106004 6384 106056 6390
rect 106004 6326 106056 6332
rect 105636 6316 105688 6322
rect 105636 6258 105688 6264
rect 105268 5704 105320 5710
rect 105268 5646 105320 5652
rect 105176 4752 105228 4758
rect 105176 4694 105228 4700
rect 105188 4078 105216 4694
rect 105176 4072 105228 4078
rect 105176 4014 105228 4020
rect 105188 3670 105216 4014
rect 105280 4010 105308 5646
rect 105452 5568 105504 5574
rect 105452 5510 105504 5516
rect 105464 4593 105492 5510
rect 105544 4616 105596 4622
rect 105450 4584 105506 4593
rect 105544 4558 105596 4564
rect 105450 4519 105506 4528
rect 105556 4214 105584 4558
rect 105544 4208 105596 4214
rect 105544 4150 105596 4156
rect 105360 4072 105412 4078
rect 105360 4014 105412 4020
rect 105268 4004 105320 4010
rect 105268 3946 105320 3952
rect 105372 3738 105400 4014
rect 105452 3936 105504 3942
rect 105452 3878 105504 3884
rect 105360 3732 105412 3738
rect 105360 3674 105412 3680
rect 105176 3664 105228 3670
rect 105176 3606 105228 3612
rect 105096 3454 105400 3482
rect 104898 3224 104954 3233
rect 104898 3159 104954 3168
rect 104992 3188 105044 3194
rect 104992 3130 105044 3136
rect 105004 2922 105032 3130
rect 105372 3058 105400 3454
rect 105360 3052 105412 3058
rect 105360 2994 105412 3000
rect 105464 2990 105492 3878
rect 105556 3534 105584 4150
rect 105648 4049 105676 6258
rect 105912 6112 105964 6118
rect 105912 6054 105964 6060
rect 105820 5160 105872 5166
rect 105820 5102 105872 5108
rect 105728 5024 105780 5030
rect 105728 4966 105780 4972
rect 105634 4040 105690 4049
rect 105634 3975 105690 3984
rect 105636 3596 105688 3602
rect 105740 3584 105768 4966
rect 105832 4282 105860 5102
rect 105820 4276 105872 4282
rect 105820 4218 105872 4224
rect 105924 4078 105952 6054
rect 106016 5953 106044 6326
rect 106002 5944 106058 5953
rect 106002 5879 106058 5888
rect 106004 5024 106056 5030
rect 106002 4992 106004 5001
rect 106056 4992 106058 5001
rect 106002 4927 106058 4936
rect 106016 4826 106044 4927
rect 106200 4865 106228 6734
rect 107016 6724 107068 6730
rect 107016 6666 107068 6672
rect 106464 6316 106516 6322
rect 106464 6258 106516 6264
rect 106372 5704 106424 5710
rect 106372 5646 106424 5652
rect 106186 4856 106242 4865
rect 106004 4820 106056 4826
rect 106004 4762 106056 4768
rect 106096 4820 106148 4826
rect 106186 4791 106242 4800
rect 106096 4762 106148 4768
rect 106108 4690 106136 4762
rect 106096 4684 106148 4690
rect 106096 4626 106148 4632
rect 106094 4584 106150 4593
rect 106094 4519 106150 4528
rect 106004 4208 106056 4214
rect 106004 4150 106056 4156
rect 106016 4078 106044 4150
rect 105912 4072 105964 4078
rect 105912 4014 105964 4020
rect 106004 4072 106056 4078
rect 106004 4014 106056 4020
rect 105818 3768 105874 3777
rect 105818 3703 105874 3712
rect 105688 3556 105768 3584
rect 105636 3538 105688 3544
rect 105544 3528 105596 3534
rect 105544 3470 105596 3476
rect 105648 3058 105676 3538
rect 105728 3460 105780 3466
rect 105728 3402 105780 3408
rect 105636 3052 105688 3058
rect 105636 2994 105688 3000
rect 105452 2984 105504 2990
rect 105452 2926 105504 2932
rect 104992 2916 105044 2922
rect 104992 2858 105044 2864
rect 105176 2916 105228 2922
rect 105176 2858 105228 2864
rect 104808 2508 104860 2514
rect 104808 2450 104860 2456
rect 104900 2304 104952 2310
rect 104900 2246 104952 2252
rect 104912 1970 104940 2246
rect 104900 1964 104952 1970
rect 104900 1906 104952 1912
rect 105084 1896 105136 1902
rect 105082 1864 105084 1873
rect 105136 1864 105138 1873
rect 104164 1828 104216 1834
rect 105082 1799 105138 1808
rect 104164 1770 104216 1776
rect 105188 1562 105216 2858
rect 105176 1556 105228 1562
rect 105176 1498 105228 1504
rect 104624 1352 104676 1358
rect 104070 1320 104126 1329
rect 104624 1294 104676 1300
rect 105544 1352 105596 1358
rect 105544 1294 105596 1300
rect 104070 1255 104126 1264
rect 103796 1012 103848 1018
rect 103796 954 103848 960
rect 103980 1012 104032 1018
rect 103980 954 104032 960
rect 103520 944 103572 950
rect 103520 886 103572 892
rect 100758 847 100814 856
rect 103336 876 103388 882
rect 103336 818 103388 824
rect 103532 377 103560 886
rect 104084 649 104112 1255
rect 104636 950 104664 1294
rect 104624 944 104676 950
rect 104162 912 104218 921
rect 104624 886 104676 892
rect 105556 882 105584 1294
rect 105648 950 105676 2994
rect 105740 2825 105768 3402
rect 105726 2816 105782 2825
rect 105726 2751 105782 2760
rect 105832 1970 105860 3703
rect 106108 3602 106136 4519
rect 106234 4480 106286 4486
rect 106286 4428 106320 4434
rect 106234 4422 106320 4428
rect 106246 4406 106320 4422
rect 106292 4321 106320 4406
rect 106278 4312 106334 4321
rect 106278 4247 106334 4256
rect 106280 4208 106332 4214
rect 106280 4150 106332 4156
rect 106292 3924 106320 4150
rect 106200 3896 106320 3924
rect 106200 3738 106228 3896
rect 106384 3738 106412 5646
rect 106476 4758 106504 6258
rect 106924 5908 106976 5914
rect 106924 5850 106976 5856
rect 106936 5030 106964 5850
rect 107028 5234 107056 6666
rect 107016 5228 107068 5234
rect 107016 5170 107068 5176
rect 106924 5024 106976 5030
rect 106924 4966 106976 4972
rect 106936 4826 106964 4966
rect 106924 4820 106976 4826
rect 106924 4762 106976 4768
rect 106464 4752 106516 4758
rect 106464 4694 106516 4700
rect 106556 4548 106608 4554
rect 106556 4490 106608 4496
rect 106188 3732 106240 3738
rect 106188 3674 106240 3680
rect 106372 3732 106424 3738
rect 106372 3674 106424 3680
rect 106568 3670 106596 4490
rect 106936 4214 106964 4762
rect 106924 4208 106976 4214
rect 106924 4150 106976 4156
rect 107120 4049 107148 7346
rect 107200 6928 107252 6934
rect 107200 6870 107252 6876
rect 107212 5914 107240 6870
rect 107568 6792 107620 6798
rect 107568 6734 107620 6740
rect 107476 6656 107528 6662
rect 107476 6598 107528 6604
rect 107384 6180 107436 6186
rect 107384 6122 107436 6128
rect 107200 5908 107252 5914
rect 107200 5850 107252 5856
rect 107292 5908 107344 5914
rect 107292 5850 107344 5856
rect 107200 5704 107252 5710
rect 107200 5646 107252 5652
rect 107212 5166 107240 5646
rect 107304 5642 107332 5850
rect 107396 5710 107424 6122
rect 107384 5704 107436 5710
rect 107384 5646 107436 5652
rect 107292 5636 107344 5642
rect 107292 5578 107344 5584
rect 107200 5160 107252 5166
rect 107200 5102 107252 5108
rect 107212 4622 107240 5102
rect 107396 4690 107424 5646
rect 107384 4684 107436 4690
rect 107384 4626 107436 4632
rect 107200 4616 107252 4622
rect 107200 4558 107252 4564
rect 107198 4312 107254 4321
rect 107198 4247 107254 4256
rect 107106 4040 107162 4049
rect 107106 3975 107162 3984
rect 106556 3664 106608 3670
rect 106556 3606 106608 3612
rect 106096 3596 106148 3602
rect 106096 3538 106148 3544
rect 106188 3528 106240 3534
rect 106186 3496 106188 3505
rect 106280 3528 106332 3534
rect 106240 3496 106242 3505
rect 106280 3470 106332 3476
rect 106186 3431 106242 3440
rect 106292 3194 106320 3470
rect 106188 3188 106240 3194
rect 106188 3130 106240 3136
rect 106280 3188 106332 3194
rect 106280 3130 106332 3136
rect 106200 2854 106228 3130
rect 106464 2984 106516 2990
rect 106464 2926 106516 2932
rect 106372 2916 106424 2922
rect 106372 2858 106424 2864
rect 106188 2848 106240 2854
rect 106188 2790 106240 2796
rect 106002 2544 106058 2553
rect 106200 2514 106228 2790
rect 106002 2479 106058 2488
rect 106188 2508 106240 2514
rect 106016 1970 106044 2479
rect 106188 2450 106240 2456
rect 106384 2378 106412 2858
rect 106372 2372 106424 2378
rect 106372 2314 106424 2320
rect 105820 1964 105872 1970
rect 105820 1906 105872 1912
rect 106004 1964 106056 1970
rect 106004 1906 106056 1912
rect 106096 1964 106148 1970
rect 106096 1906 106148 1912
rect 106004 1420 106056 1426
rect 106108 1408 106136 1906
rect 106056 1380 106136 1408
rect 106004 1362 106056 1368
rect 106476 1358 106504 2926
rect 107212 2514 107240 4247
rect 107396 3505 107424 4626
rect 107488 4486 107516 6598
rect 107476 4480 107528 4486
rect 107476 4422 107528 4428
rect 107580 4049 107608 6734
rect 107660 5636 107712 5642
rect 107660 5578 107712 5584
rect 107672 5234 107700 5578
rect 107660 5228 107712 5234
rect 107660 5170 107712 5176
rect 107764 5114 107792 7822
rect 109052 7750 109080 9386
rect 109592 8084 109644 8090
rect 109592 8026 109644 8032
rect 109604 7886 109632 8026
rect 109316 7880 109368 7886
rect 109316 7822 109368 7828
rect 109592 7880 109644 7886
rect 109592 7822 109644 7828
rect 109040 7744 109092 7750
rect 109040 7686 109092 7692
rect 107844 7540 107896 7546
rect 107844 7482 107896 7488
rect 107672 5086 107792 5114
rect 107566 4040 107622 4049
rect 107566 3975 107622 3984
rect 107382 3496 107438 3505
rect 107672 3482 107700 5086
rect 107856 3942 107884 7482
rect 108856 7472 108908 7478
rect 108856 7414 108908 7420
rect 108396 6996 108448 7002
rect 108396 6938 108448 6944
rect 108764 6996 108816 7002
rect 108764 6938 108816 6944
rect 107936 6656 107988 6662
rect 107936 6598 107988 6604
rect 108028 6656 108080 6662
rect 108028 6598 108080 6604
rect 107844 3936 107896 3942
rect 107844 3878 107896 3884
rect 107672 3454 107792 3482
rect 107382 3431 107438 3440
rect 107660 3392 107712 3398
rect 107660 3334 107712 3340
rect 107672 2650 107700 3334
rect 107764 2774 107792 3454
rect 107764 2746 107884 2774
rect 107568 2644 107620 2650
rect 107568 2586 107620 2592
rect 107660 2644 107712 2650
rect 107660 2586 107712 2592
rect 107200 2508 107252 2514
rect 107200 2450 107252 2456
rect 107580 2258 107608 2586
rect 107672 2514 107700 2586
rect 107660 2508 107712 2514
rect 107660 2450 107712 2456
rect 107856 2310 107884 2746
rect 107844 2304 107896 2310
rect 107580 2230 107792 2258
rect 107844 2246 107896 2252
rect 107764 2106 107792 2230
rect 107660 2100 107712 2106
rect 107660 2042 107712 2048
rect 107752 2100 107804 2106
rect 107752 2042 107804 2048
rect 107672 1902 107700 2042
rect 107948 2038 107976 6598
rect 108040 6458 108068 6598
rect 108028 6452 108080 6458
rect 108028 6394 108080 6400
rect 108210 6216 108266 6225
rect 108210 6151 108212 6160
rect 108264 6151 108266 6160
rect 108212 6122 108264 6128
rect 108224 5846 108252 6122
rect 108212 5840 108264 5846
rect 108212 5782 108264 5788
rect 108120 5568 108172 5574
rect 108120 5510 108172 5516
rect 108028 5296 108080 5302
rect 108028 5238 108080 5244
rect 108040 4049 108068 5238
rect 108132 4842 108160 5510
rect 108132 4826 108252 4842
rect 108132 4820 108264 4826
rect 108132 4814 108212 4820
rect 108212 4762 108264 4768
rect 108120 4616 108172 4622
rect 108120 4558 108172 4564
rect 108132 4214 108160 4558
rect 108120 4208 108172 4214
rect 108120 4150 108172 4156
rect 108120 4072 108172 4078
rect 108026 4040 108082 4049
rect 108120 4014 108172 4020
rect 108026 3975 108082 3984
rect 108132 3505 108160 4014
rect 108118 3496 108174 3505
rect 108118 3431 108174 3440
rect 108408 2774 108436 6938
rect 108580 6792 108632 6798
rect 108580 6734 108632 6740
rect 108672 6792 108724 6798
rect 108672 6734 108724 6740
rect 108592 6322 108620 6734
rect 108580 6316 108632 6322
rect 108580 6258 108632 6264
rect 108592 5234 108620 6258
rect 108684 6254 108712 6734
rect 108672 6248 108724 6254
rect 108672 6190 108724 6196
rect 108684 5574 108712 6190
rect 108776 6118 108804 6938
rect 108764 6112 108816 6118
rect 108764 6054 108816 6060
rect 108776 5846 108804 6054
rect 108764 5840 108816 5846
rect 108764 5782 108816 5788
rect 108672 5568 108724 5574
rect 108672 5510 108724 5516
rect 108684 5234 108712 5510
rect 108580 5228 108632 5234
rect 108580 5170 108632 5176
rect 108672 5228 108724 5234
rect 108672 5170 108724 5176
rect 108776 5030 108804 5782
rect 108868 5370 108896 7414
rect 109040 7404 109092 7410
rect 109040 7346 109092 7352
rect 109052 7002 109080 7346
rect 109132 7336 109184 7342
rect 109132 7278 109184 7284
rect 109040 6996 109092 7002
rect 109040 6938 109092 6944
rect 108948 6112 109000 6118
rect 108948 6054 109000 6060
rect 108960 5778 108988 6054
rect 109038 5808 109094 5817
rect 108948 5772 109000 5778
rect 109038 5743 109040 5752
rect 108948 5714 109000 5720
rect 109092 5743 109094 5752
rect 109040 5714 109092 5720
rect 109144 5658 109172 7278
rect 109224 7200 109276 7206
rect 109224 7142 109276 7148
rect 109236 5778 109264 7142
rect 109328 6458 109356 7822
rect 109500 7744 109552 7750
rect 109500 7686 109552 7692
rect 109408 6724 109460 6730
rect 109408 6666 109460 6672
rect 109316 6452 109368 6458
rect 109316 6394 109368 6400
rect 109316 6248 109368 6254
rect 109316 6190 109368 6196
rect 109224 5772 109276 5778
rect 109224 5714 109276 5720
rect 109144 5630 109264 5658
rect 108856 5364 108908 5370
rect 108856 5306 108908 5312
rect 109130 5128 109186 5137
rect 109130 5063 109186 5072
rect 108764 5024 108816 5030
rect 108670 4992 108726 5001
rect 108764 4966 108816 4972
rect 108670 4927 108726 4936
rect 108316 2746 108436 2774
rect 108316 2038 108344 2746
rect 108684 2650 108712 4927
rect 109144 4622 109172 5063
rect 108764 4616 108816 4622
rect 108764 4558 108816 4564
rect 109132 4616 109184 4622
rect 109132 4558 109184 4564
rect 108776 4146 108804 4558
rect 108764 4140 108816 4146
rect 108764 4082 108816 4088
rect 108856 4072 108908 4078
rect 109236 4049 109264 5630
rect 108856 4014 108908 4020
rect 109222 4040 109278 4049
rect 108764 4004 108816 4010
rect 108764 3946 108816 3952
rect 108776 3738 108804 3946
rect 108868 3942 108896 4014
rect 109222 3975 109278 3984
rect 109328 3942 109356 6190
rect 108856 3936 108908 3942
rect 108856 3878 108908 3884
rect 109316 3936 109368 3942
rect 109316 3878 109368 3884
rect 108854 3768 108910 3777
rect 108764 3732 108816 3738
rect 108854 3703 108910 3712
rect 108764 3674 108816 3680
rect 108868 3602 108896 3703
rect 109420 3602 109448 6666
rect 108856 3596 108908 3602
rect 108856 3538 108908 3544
rect 109408 3596 109460 3602
rect 109408 3538 109460 3544
rect 108946 3224 109002 3233
rect 108946 3159 109002 3168
rect 108960 2990 108988 3159
rect 108948 2984 109000 2990
rect 108948 2926 109000 2932
rect 108672 2644 108724 2650
rect 108672 2586 108724 2592
rect 108764 2644 108816 2650
rect 108764 2586 108816 2592
rect 108488 2440 108540 2446
rect 108488 2382 108540 2388
rect 107936 2032 107988 2038
rect 107936 1974 107988 1980
rect 108304 2032 108356 2038
rect 108304 1974 108356 1980
rect 107660 1896 107712 1902
rect 107660 1838 107712 1844
rect 107764 1822 107976 1850
rect 107764 1562 107792 1822
rect 107948 1766 107976 1822
rect 107844 1760 107896 1766
rect 107844 1702 107896 1708
rect 107936 1760 107988 1766
rect 107936 1702 107988 1708
rect 107752 1556 107804 1562
rect 107752 1498 107804 1504
rect 107856 1494 107884 1702
rect 107844 1488 107896 1494
rect 107844 1430 107896 1436
rect 105728 1352 105780 1358
rect 105728 1294 105780 1300
rect 106464 1352 106516 1358
rect 106464 1294 106516 1300
rect 107200 1352 107252 1358
rect 107200 1294 107252 1300
rect 107384 1352 107436 1358
rect 107384 1294 107436 1300
rect 108120 1352 108172 1358
rect 108120 1294 108172 1300
rect 108304 1352 108356 1358
rect 108304 1294 108356 1300
rect 105636 944 105688 950
rect 105636 886 105688 892
rect 104162 847 104218 856
rect 105544 876 105596 882
rect 104070 640 104126 649
rect 104070 575 104126 584
rect 103518 368 103574 377
rect 103518 303 103574 312
rect 100484 264 100536 270
rect 104176 241 104204 847
rect 105544 818 105596 824
rect 105740 474 105768 1294
rect 107212 678 107240 1294
rect 107396 1222 107424 1294
rect 107384 1216 107436 1222
rect 107384 1158 107436 1164
rect 107200 672 107252 678
rect 107200 614 107252 620
rect 107396 542 107424 1158
rect 108132 678 108160 1294
rect 108316 950 108344 1294
rect 108304 944 108356 950
rect 108304 886 108356 892
rect 108500 785 108528 2382
rect 108580 2304 108632 2310
rect 108580 2246 108632 2252
rect 108592 1834 108620 2246
rect 108776 2106 108804 2586
rect 109512 2514 109540 7686
rect 109590 6352 109646 6361
rect 109590 6287 109592 6296
rect 109644 6287 109646 6296
rect 109592 6258 109644 6264
rect 109592 2848 109644 2854
rect 109590 2816 109592 2825
rect 109644 2816 109646 2825
rect 109590 2751 109646 2760
rect 109040 2508 109092 2514
rect 109040 2450 109092 2456
rect 109500 2508 109552 2514
rect 109500 2450 109552 2456
rect 108764 2100 108816 2106
rect 108764 2042 108816 2048
rect 108580 1828 108632 1834
rect 108580 1770 108632 1776
rect 109052 1494 109080 2450
rect 109132 1896 109184 1902
rect 109132 1838 109184 1844
rect 109040 1488 109092 1494
rect 109040 1430 109092 1436
rect 108948 1284 109000 1290
rect 108948 1226 109000 1232
rect 108960 1018 108988 1226
rect 108948 1012 109000 1018
rect 108948 954 109000 960
rect 109144 950 109172 1838
rect 109222 1456 109278 1465
rect 109222 1391 109224 1400
rect 109276 1391 109278 1400
rect 109224 1362 109276 1368
rect 109132 944 109184 950
rect 109132 886 109184 892
rect 109696 882 109724 9386
rect 110524 8786 110552 9930
rect 110800 9586 110828 10231
rect 111536 9586 111564 10231
rect 110788 9580 110840 9586
rect 110788 9522 110840 9528
rect 111524 9580 111576 9586
rect 111524 9522 111576 9528
rect 112076 9444 112128 9450
rect 112076 9386 112128 9392
rect 110604 9376 110656 9382
rect 110604 9318 110656 9324
rect 110616 8906 110644 9318
rect 111892 9172 111944 9178
rect 111892 9114 111944 9120
rect 111156 9104 111208 9110
rect 111156 9046 111208 9052
rect 110604 8900 110656 8906
rect 110604 8842 110656 8848
rect 110524 8758 110644 8786
rect 110052 7880 110104 7886
rect 110052 7822 110104 7828
rect 109776 7268 109828 7274
rect 109776 7210 109828 7216
rect 109788 6390 109816 7210
rect 109960 6792 110012 6798
rect 109960 6734 110012 6740
rect 109972 6662 110000 6734
rect 109960 6656 110012 6662
rect 109960 6598 110012 6604
rect 109776 6384 109828 6390
rect 109776 6326 109828 6332
rect 109972 5846 110000 6598
rect 109960 5840 110012 5846
rect 109960 5782 110012 5788
rect 109776 5024 109828 5030
rect 109776 4966 109828 4972
rect 109960 5024 110012 5030
rect 109960 4966 110012 4972
rect 109788 3942 109816 4966
rect 109972 4146 110000 4966
rect 109960 4140 110012 4146
rect 109960 4082 110012 4088
rect 110064 4049 110092 7822
rect 110236 6996 110288 7002
rect 110236 6938 110288 6944
rect 110144 6860 110196 6866
rect 110144 6802 110196 6808
rect 110050 4040 110106 4049
rect 110050 3975 110106 3984
rect 109776 3936 109828 3942
rect 109776 3878 109828 3884
rect 110156 2553 110184 6802
rect 110248 5642 110276 6938
rect 110420 6792 110472 6798
rect 110420 6734 110472 6740
rect 110432 6458 110460 6734
rect 110420 6452 110472 6458
rect 110420 6394 110472 6400
rect 110432 5710 110460 6394
rect 110420 5704 110472 5710
rect 110420 5646 110472 5652
rect 110236 5636 110288 5642
rect 110236 5578 110288 5584
rect 110512 5228 110564 5234
rect 110512 5170 110564 5176
rect 110236 5160 110288 5166
rect 110236 5102 110288 5108
rect 110248 4146 110276 5102
rect 110236 4140 110288 4146
rect 110236 4082 110288 4088
rect 110248 3058 110276 4082
rect 110524 4078 110552 5170
rect 110512 4072 110564 4078
rect 110512 4014 110564 4020
rect 110328 3936 110380 3942
rect 110328 3878 110380 3884
rect 110236 3052 110288 3058
rect 110236 2994 110288 3000
rect 110340 2904 110368 3878
rect 110420 3596 110472 3602
rect 110420 3538 110472 3544
rect 110432 3398 110460 3538
rect 110420 3392 110472 3398
rect 110420 3334 110472 3340
rect 110524 2990 110552 4014
rect 110512 2984 110564 2990
rect 110512 2926 110564 2932
rect 110420 2916 110472 2922
rect 110340 2876 110420 2904
rect 110420 2858 110472 2864
rect 110616 2774 110644 8758
rect 110696 7404 110748 7410
rect 110696 7346 110748 7352
rect 110708 4049 110736 7346
rect 111064 7200 111116 7206
rect 111064 7142 111116 7148
rect 110972 6928 111024 6934
rect 110972 6870 111024 6876
rect 110984 6798 111012 6870
rect 110972 6792 111024 6798
rect 110972 6734 111024 6740
rect 110972 6656 111024 6662
rect 110972 6598 111024 6604
rect 110880 5636 110932 5642
rect 110880 5578 110932 5584
rect 110786 5264 110842 5273
rect 110786 5199 110788 5208
rect 110840 5199 110842 5208
rect 110788 5170 110840 5176
rect 110892 4690 110920 5578
rect 110984 5302 111012 6598
rect 110972 5296 111024 5302
rect 110972 5238 111024 5244
rect 110880 4684 110932 4690
rect 110880 4626 110932 4632
rect 110788 4072 110840 4078
rect 110694 4040 110750 4049
rect 110788 4014 110840 4020
rect 110694 3975 110750 3984
rect 110800 3890 110828 4014
rect 110708 3862 110828 3890
rect 110708 3602 110736 3862
rect 110696 3596 110748 3602
rect 110696 3538 110748 3544
rect 110880 3528 110932 3534
rect 110880 3470 110932 3476
rect 110524 2746 110644 2774
rect 110142 2544 110198 2553
rect 110326 2544 110382 2553
rect 110142 2479 110198 2488
rect 110248 2502 110326 2530
rect 110248 2310 110276 2502
rect 110326 2479 110382 2488
rect 110236 2304 110288 2310
rect 110236 2246 110288 2252
rect 110248 1970 110276 2246
rect 110328 2032 110380 2038
rect 110328 1974 110380 1980
rect 110236 1964 110288 1970
rect 110236 1906 110288 1912
rect 109960 1352 110012 1358
rect 109960 1294 110012 1300
rect 109684 876 109736 882
rect 109684 818 109736 824
rect 108486 776 108542 785
rect 109972 746 110000 1294
rect 110340 1222 110368 1974
rect 110524 1970 110552 2746
rect 110696 2440 110748 2446
rect 110696 2382 110748 2388
rect 110512 1964 110564 1970
rect 110512 1906 110564 1912
rect 110708 1426 110736 2382
rect 110892 2106 110920 3470
rect 111076 2774 111104 7142
rect 111168 4078 111196 9046
rect 111340 8832 111392 8838
rect 111340 8774 111392 8780
rect 111352 7410 111380 8774
rect 111524 8288 111576 8294
rect 111524 8230 111576 8236
rect 111536 7546 111564 8230
rect 111524 7540 111576 7546
rect 111524 7482 111576 7488
rect 111616 7540 111668 7546
rect 111616 7482 111668 7488
rect 111248 7404 111300 7410
rect 111248 7346 111300 7352
rect 111340 7404 111392 7410
rect 111340 7346 111392 7352
rect 111156 4072 111208 4078
rect 111260 4049 111288 7346
rect 111340 6656 111392 6662
rect 111340 6598 111392 6604
rect 111156 4014 111208 4020
rect 111246 4040 111302 4049
rect 111246 3975 111302 3984
rect 111248 3392 111300 3398
rect 111352 3380 111380 6598
rect 111432 5636 111484 5642
rect 111432 5578 111484 5584
rect 111444 5545 111472 5578
rect 111430 5536 111486 5545
rect 111430 5471 111486 5480
rect 111430 5264 111486 5273
rect 111430 5199 111486 5208
rect 111444 5098 111472 5199
rect 111432 5092 111484 5098
rect 111432 5034 111484 5040
rect 111628 4706 111656 7482
rect 111536 4678 111656 4706
rect 111536 3602 111564 4678
rect 111616 4616 111668 4622
rect 111616 4558 111668 4564
rect 111628 4282 111656 4558
rect 111800 4480 111852 4486
rect 111800 4422 111852 4428
rect 111616 4276 111668 4282
rect 111616 4218 111668 4224
rect 111812 4078 111840 4422
rect 111616 4072 111668 4078
rect 111616 4014 111668 4020
rect 111800 4072 111852 4078
rect 111800 4014 111852 4020
rect 111628 3738 111656 4014
rect 111708 3936 111760 3942
rect 111708 3878 111760 3884
rect 111720 3738 111748 3878
rect 111616 3732 111668 3738
rect 111616 3674 111668 3680
rect 111708 3732 111760 3738
rect 111708 3674 111760 3680
rect 111524 3596 111576 3602
rect 111524 3538 111576 3544
rect 111800 3596 111852 3602
rect 111800 3538 111852 3544
rect 111300 3352 111380 3380
rect 111248 3334 111300 3340
rect 110984 2746 111104 2774
rect 111260 2774 111288 3334
rect 111616 2984 111668 2990
rect 111616 2926 111668 2932
rect 111260 2746 111380 2774
rect 110880 2100 110932 2106
rect 110880 2042 110932 2048
rect 110880 1896 110932 1902
rect 110880 1838 110932 1844
rect 110696 1420 110748 1426
rect 110696 1362 110748 1368
rect 110788 1352 110840 1358
rect 110788 1294 110840 1300
rect 110328 1216 110380 1222
rect 110328 1158 110380 1164
rect 110800 1018 110828 1294
rect 110696 1012 110748 1018
rect 110696 954 110748 960
rect 110788 1012 110840 1018
rect 110788 954 110840 960
rect 110708 746 110736 954
rect 110892 814 110920 1838
rect 110880 808 110932 814
rect 110880 750 110932 756
rect 108486 711 108542 720
rect 109960 740 110012 746
rect 109960 682 110012 688
rect 110696 740 110748 746
rect 110696 682 110748 688
rect 108120 672 108172 678
rect 108120 614 108172 620
rect 107384 536 107436 542
rect 107384 478 107436 484
rect 110984 474 111012 2746
rect 111352 1834 111380 2746
rect 111340 1828 111392 1834
rect 111340 1770 111392 1776
rect 111352 1562 111380 1770
rect 111340 1556 111392 1562
rect 111340 1498 111392 1504
rect 111338 1456 111394 1465
rect 111338 1391 111340 1400
rect 111392 1391 111394 1400
rect 111340 1362 111392 1368
rect 111628 1358 111656 2926
rect 111708 2916 111760 2922
rect 111708 2858 111760 2864
rect 111720 2825 111748 2858
rect 111706 2816 111762 2825
rect 111706 2751 111762 2760
rect 111812 1952 111840 3538
rect 111904 2774 111932 9114
rect 111984 4684 112036 4690
rect 111984 4626 112036 4632
rect 111996 4078 112024 4626
rect 111984 4072 112036 4078
rect 111984 4014 112036 4020
rect 111904 2746 112024 2774
rect 111892 1964 111944 1970
rect 111812 1924 111892 1952
rect 111812 1426 111840 1924
rect 111892 1906 111944 1912
rect 111996 1766 112024 2746
rect 112088 2446 112116 9386
rect 112364 8974 112392 10231
rect 112916 9586 112944 10231
rect 113560 9586 113588 10231
rect 113824 9716 113876 9722
rect 113824 9658 113876 9664
rect 112904 9580 112956 9586
rect 112904 9522 112956 9528
rect 113548 9580 113600 9586
rect 113548 9522 113600 9528
rect 112628 9376 112680 9382
rect 112628 9318 112680 9324
rect 113180 9376 113232 9382
rect 113180 9318 113232 9324
rect 112352 8968 112404 8974
rect 112352 8910 112404 8916
rect 112168 8832 112220 8838
rect 112168 8774 112220 8780
rect 112180 6905 112208 8774
rect 112536 7268 112588 7274
rect 112536 7210 112588 7216
rect 112548 6934 112576 7210
rect 112536 6928 112588 6934
rect 112166 6896 112222 6905
rect 112536 6870 112588 6876
rect 112166 6831 112222 6840
rect 112352 6792 112404 6798
rect 112352 6734 112404 6740
rect 112260 6112 112312 6118
rect 112260 6054 112312 6060
rect 112168 5908 112220 5914
rect 112168 5850 112220 5856
rect 112180 5710 112208 5850
rect 112168 5704 112220 5710
rect 112168 5646 112220 5652
rect 112168 4004 112220 4010
rect 112168 3946 112220 3952
rect 112180 3466 112208 3946
rect 112168 3460 112220 3466
rect 112168 3402 112220 3408
rect 112272 2774 112300 6054
rect 112364 4049 112392 6734
rect 112548 6662 112576 6870
rect 112536 6656 112588 6662
rect 112536 6598 112588 6604
rect 112350 4040 112406 4049
rect 112350 3975 112406 3984
rect 112536 3596 112588 3602
rect 112536 3538 112588 3544
rect 112272 2746 112392 2774
rect 112076 2440 112128 2446
rect 112076 2382 112128 2388
rect 112168 2440 112220 2446
rect 112168 2382 112220 2388
rect 111984 1760 112036 1766
rect 111984 1702 112036 1708
rect 111800 1420 111852 1426
rect 111800 1362 111852 1368
rect 111616 1352 111668 1358
rect 111616 1294 111668 1300
rect 112180 1222 112208 2382
rect 112364 2378 112392 2746
rect 112352 2372 112404 2378
rect 112352 2314 112404 2320
rect 112548 2106 112576 3538
rect 112536 2100 112588 2106
rect 112536 2042 112588 2048
rect 112352 1352 112404 1358
rect 112352 1294 112404 1300
rect 112168 1216 112220 1222
rect 112364 1193 112392 1294
rect 112168 1158 112220 1164
rect 112350 1184 112406 1193
rect 112350 1119 112406 1128
rect 112640 678 112668 9318
rect 112812 7948 112864 7954
rect 112812 7890 112864 7896
rect 112824 7410 112852 7890
rect 113088 7540 113140 7546
rect 113088 7482 113140 7488
rect 113100 7410 113128 7482
rect 112812 7404 112864 7410
rect 112812 7346 112864 7352
rect 113088 7404 113140 7410
rect 113088 7346 113140 7352
rect 112996 6792 113048 6798
rect 112996 6734 113048 6740
rect 112812 6656 112864 6662
rect 112812 6598 112864 6604
rect 112720 6112 112772 6118
rect 112720 6054 112772 6060
rect 112732 5914 112760 6054
rect 112720 5908 112772 5914
rect 112720 5850 112772 5856
rect 112824 746 112852 6598
rect 112902 6216 112958 6225
rect 112902 6151 112958 6160
rect 112916 5846 112944 6151
rect 112904 5840 112956 5846
rect 112904 5782 112956 5788
rect 113008 4049 113036 6734
rect 113088 6724 113140 6730
rect 113088 6666 113140 6672
rect 113100 5817 113128 6666
rect 113086 5808 113142 5817
rect 113086 5743 113142 5752
rect 113086 5128 113142 5137
rect 113086 5063 113142 5072
rect 113100 4622 113128 5063
rect 113088 4616 113140 4622
rect 113088 4558 113140 4564
rect 112994 4040 113050 4049
rect 112994 3975 113050 3984
rect 113088 1352 113140 1358
rect 113192 1340 113220 9318
rect 113836 8362 113864 9658
rect 114204 9586 114232 10231
rect 115216 9586 115244 10231
rect 115768 9586 115796 10231
rect 116688 9586 116716 10231
rect 117044 9920 117096 9926
rect 117044 9862 117096 9868
rect 114192 9580 114244 9586
rect 114192 9522 114244 9528
rect 115204 9580 115256 9586
rect 115204 9522 115256 9528
rect 115756 9580 115808 9586
rect 115756 9522 115808 9528
rect 116676 9580 116728 9586
rect 116676 9522 116728 9528
rect 116032 9444 116084 9450
rect 116032 9386 116084 9392
rect 115020 9376 115072 9382
rect 115020 9318 115072 9324
rect 115756 9376 115808 9382
rect 115756 9318 115808 9324
rect 115848 9376 115900 9382
rect 115848 9318 115900 9324
rect 115032 9178 115060 9318
rect 115020 9172 115072 9178
rect 115020 9114 115072 9120
rect 115768 9110 115796 9318
rect 115756 9104 115808 9110
rect 115756 9046 115808 9052
rect 113824 8356 113876 8362
rect 113824 8298 113876 8304
rect 113822 8120 113878 8129
rect 113822 8055 113878 8064
rect 113272 7200 113324 7206
rect 113272 7142 113324 7148
rect 113732 7200 113784 7206
rect 113732 7142 113784 7148
rect 113284 6390 113312 7142
rect 113548 6928 113600 6934
rect 113548 6870 113600 6876
rect 113560 6390 113588 6870
rect 113744 6866 113772 7142
rect 113732 6860 113784 6866
rect 113732 6802 113784 6808
rect 113272 6384 113324 6390
rect 113548 6384 113600 6390
rect 113272 6326 113324 6332
rect 113454 6352 113510 6361
rect 113284 5930 113312 6326
rect 113548 6326 113600 6332
rect 113454 6287 113456 6296
rect 113508 6287 113510 6296
rect 113732 6316 113784 6322
rect 113456 6258 113508 6264
rect 113732 6258 113784 6264
rect 113468 6186 113496 6258
rect 113456 6180 113508 6186
rect 113456 6122 113508 6128
rect 113284 5902 113496 5930
rect 113364 5840 113416 5846
rect 113364 5782 113416 5788
rect 113376 5030 113404 5782
rect 113364 5024 113416 5030
rect 113364 4966 113416 4972
rect 113364 4752 113416 4758
rect 113364 4694 113416 4700
rect 113376 4554 113404 4694
rect 113364 4548 113416 4554
rect 113364 4490 113416 4496
rect 113362 3496 113418 3505
rect 113362 3431 113418 3440
rect 113376 3194 113404 3431
rect 113364 3188 113416 3194
rect 113364 3130 113416 3136
rect 113468 2990 113496 5902
rect 113744 5778 113772 6258
rect 113732 5772 113784 5778
rect 113732 5714 113784 5720
rect 113640 5568 113692 5574
rect 113640 5510 113692 5516
rect 113546 5400 113602 5409
rect 113546 5335 113602 5344
rect 113560 5302 113588 5335
rect 113548 5296 113600 5302
rect 113548 5238 113600 5244
rect 113548 4684 113600 4690
rect 113652 4672 113680 5510
rect 113744 5302 113772 5714
rect 113732 5296 113784 5302
rect 113732 5238 113784 5244
rect 113744 5166 113772 5238
rect 113732 5160 113784 5166
rect 113732 5102 113784 5108
rect 113836 5012 113864 8055
rect 115388 7880 115440 7886
rect 114006 7848 114062 7857
rect 115388 7822 115440 7828
rect 114006 7783 114062 7792
rect 115296 7812 115348 7818
rect 113916 6724 113968 6730
rect 113916 6666 113968 6672
rect 113928 6458 113956 6666
rect 113916 6452 113968 6458
rect 113916 6394 113968 6400
rect 114020 5574 114048 7783
rect 115296 7754 115348 7760
rect 114928 7744 114980 7750
rect 114928 7686 114980 7692
rect 115112 7744 115164 7750
rect 115112 7686 115164 7692
rect 115204 7744 115256 7750
rect 115204 7686 115256 7692
rect 114652 6928 114704 6934
rect 114652 6870 114704 6876
rect 114560 6860 114612 6866
rect 114560 6802 114612 6808
rect 114572 6633 114600 6802
rect 114558 6624 114614 6633
rect 114558 6559 114614 6568
rect 114192 5704 114244 5710
rect 114192 5646 114244 5652
rect 114008 5568 114060 5574
rect 114008 5510 114060 5516
rect 114204 5234 114232 5646
rect 114468 5636 114520 5642
rect 114468 5578 114520 5584
rect 114480 5545 114508 5578
rect 114466 5536 114522 5545
rect 114466 5471 114522 5480
rect 114572 5409 114600 6559
rect 114664 6118 114692 6870
rect 114742 6352 114798 6361
rect 114742 6287 114798 6296
rect 114652 6112 114704 6118
rect 114652 6054 114704 6060
rect 114756 5846 114784 6287
rect 114834 6216 114890 6225
rect 114834 6151 114890 6160
rect 114848 5914 114876 6151
rect 114836 5908 114888 5914
rect 114836 5850 114888 5856
rect 114652 5840 114704 5846
rect 114652 5782 114704 5788
rect 114744 5840 114796 5846
rect 114744 5782 114796 5788
rect 114558 5400 114614 5409
rect 114558 5335 114614 5344
rect 114284 5296 114336 5302
rect 114284 5238 114336 5244
rect 114192 5228 114244 5234
rect 114192 5170 114244 5176
rect 114204 5114 114232 5170
rect 114112 5086 114232 5114
rect 113600 4644 113680 4672
rect 113744 4984 113864 5012
rect 114008 5024 114060 5030
rect 113548 4626 113600 4632
rect 113744 4486 113772 4984
rect 114008 4966 114060 4972
rect 114020 4826 114048 4966
rect 113824 4820 113876 4826
rect 113824 4762 113876 4768
rect 114008 4820 114060 4826
rect 114008 4762 114060 4768
rect 113732 4480 113784 4486
rect 113732 4422 113784 4428
rect 113744 3602 113772 4422
rect 113732 3596 113784 3602
rect 113732 3538 113784 3544
rect 113456 2984 113508 2990
rect 113456 2926 113508 2932
rect 113836 2514 113864 4762
rect 114112 4622 114140 5086
rect 114192 5024 114244 5030
rect 114192 4966 114244 4972
rect 114100 4616 114152 4622
rect 114100 4558 114152 4564
rect 114204 4146 114232 4966
rect 114296 4622 114324 5238
rect 114664 5137 114692 5782
rect 114940 5302 114968 7686
rect 115124 7342 115152 7686
rect 115216 7410 115244 7686
rect 115308 7546 115336 7754
rect 115400 7546 115428 7822
rect 115756 7812 115808 7818
rect 115756 7754 115808 7760
rect 115480 7744 115532 7750
rect 115480 7686 115532 7692
rect 115296 7540 115348 7546
rect 115296 7482 115348 7488
rect 115388 7540 115440 7546
rect 115388 7482 115440 7488
rect 115204 7404 115256 7410
rect 115204 7346 115256 7352
rect 115112 7336 115164 7342
rect 115112 7278 115164 7284
rect 115400 6662 115428 7482
rect 115492 7449 115520 7686
rect 115478 7440 115534 7449
rect 115478 7375 115534 7384
rect 115572 7404 115624 7410
rect 115572 7346 115624 7352
rect 115480 7336 115532 7342
rect 115480 7278 115532 7284
rect 115112 6656 115164 6662
rect 115112 6598 115164 6604
rect 115388 6656 115440 6662
rect 115388 6598 115440 6604
rect 115018 6488 115074 6497
rect 115018 6423 115074 6432
rect 115032 6322 115060 6423
rect 115020 6316 115072 6322
rect 115020 6258 115072 6264
rect 115020 6180 115072 6186
rect 115020 6122 115072 6128
rect 114928 5296 114980 5302
rect 115032 5273 115060 6122
rect 115124 5710 115152 6598
rect 115492 6458 115520 7278
rect 115584 6780 115612 7346
rect 115662 7304 115718 7313
rect 115662 7239 115664 7248
rect 115716 7239 115718 7248
rect 115664 7210 115716 7216
rect 115664 6792 115716 6798
rect 115584 6752 115664 6780
rect 115664 6734 115716 6740
rect 115204 6452 115256 6458
rect 115204 6394 115256 6400
rect 115480 6452 115532 6458
rect 115480 6394 115532 6400
rect 115216 5778 115244 6394
rect 115204 5772 115256 5778
rect 115204 5714 115256 5720
rect 115676 5710 115704 6734
rect 115768 5778 115796 7754
rect 115756 5772 115808 5778
rect 115756 5714 115808 5720
rect 115112 5704 115164 5710
rect 115112 5646 115164 5652
rect 115664 5704 115716 5710
rect 115664 5646 115716 5652
rect 115204 5364 115256 5370
rect 115204 5306 115256 5312
rect 114928 5238 114980 5244
rect 115018 5264 115074 5273
rect 115018 5199 115074 5208
rect 114650 5128 114706 5137
rect 114468 5092 114520 5098
rect 114650 5063 114706 5072
rect 115112 5092 115164 5098
rect 114468 5034 114520 5040
rect 115112 5034 115164 5040
rect 114376 5024 114428 5030
rect 114376 4966 114428 4972
rect 114388 4826 114416 4966
rect 114480 4826 114508 5034
rect 114376 4820 114428 4826
rect 114376 4762 114428 4768
rect 114468 4820 114520 4826
rect 114468 4762 114520 4768
rect 114836 4752 114888 4758
rect 114836 4694 114888 4700
rect 114926 4720 114982 4729
rect 114284 4616 114336 4622
rect 114284 4558 114336 4564
rect 114558 4584 114614 4593
rect 114558 4519 114614 4528
rect 114192 4140 114244 4146
rect 114192 4082 114244 4088
rect 114572 4078 114600 4519
rect 114560 4072 114612 4078
rect 114560 4014 114612 4020
rect 114744 4072 114796 4078
rect 114744 4014 114796 4020
rect 114756 2650 114784 4014
rect 114848 3602 114876 4694
rect 115124 4690 115152 5034
rect 114926 4655 114982 4664
rect 115112 4684 115164 4690
rect 114940 4622 114968 4655
rect 115112 4626 115164 4632
rect 114928 4616 114980 4622
rect 114928 4558 114980 4564
rect 115018 3632 115074 3641
rect 114836 3596 114888 3602
rect 115018 3567 115074 3576
rect 114836 3538 114888 3544
rect 114928 3528 114980 3534
rect 114928 3470 114980 3476
rect 114940 2961 114968 3470
rect 115032 3058 115060 3567
rect 115020 3052 115072 3058
rect 115020 2994 115072 3000
rect 115216 2990 115244 5306
rect 115204 2984 115256 2990
rect 114926 2952 114982 2961
rect 115204 2926 115256 2932
rect 114926 2887 114982 2896
rect 114744 2644 114796 2650
rect 114744 2586 114796 2592
rect 114560 2576 114612 2582
rect 114560 2518 114612 2524
rect 113364 2508 113416 2514
rect 113364 2450 113416 2456
rect 113824 2508 113876 2514
rect 113824 2450 113876 2456
rect 113140 1312 113220 1340
rect 113272 1352 113324 1358
rect 113088 1294 113140 1300
rect 113272 1294 113324 1300
rect 113284 950 113312 1294
rect 113272 944 113324 950
rect 113272 886 113324 892
rect 112812 740 112864 746
rect 112812 682 112864 688
rect 113376 678 113404 2450
rect 114572 2281 114600 2518
rect 115020 2304 115072 2310
rect 114558 2272 114614 2281
rect 115020 2246 115072 2252
rect 114558 2207 114614 2216
rect 114560 2100 114612 2106
rect 114560 2042 114612 2048
rect 114572 1465 114600 2042
rect 115032 1902 115060 2246
rect 114836 1896 114888 1902
rect 114836 1838 114888 1844
rect 115020 1896 115072 1902
rect 115020 1838 115072 1844
rect 115204 1896 115256 1902
rect 115204 1838 115256 1844
rect 115572 1896 115624 1902
rect 115572 1838 115624 1844
rect 114848 1465 114876 1838
rect 114558 1456 114614 1465
rect 114558 1391 114614 1400
rect 114834 1456 114890 1465
rect 114834 1391 114890 1400
rect 114928 1352 114980 1358
rect 114928 1294 114980 1300
rect 115112 1352 115164 1358
rect 115112 1294 115164 1300
rect 114940 1222 114968 1294
rect 114928 1216 114980 1222
rect 114928 1158 114980 1164
rect 114940 921 114968 1158
rect 115124 1057 115152 1294
rect 115110 1048 115166 1057
rect 115110 983 115166 992
rect 114926 912 114982 921
rect 114926 847 114982 856
rect 112628 672 112680 678
rect 112628 614 112680 620
rect 113364 672 113416 678
rect 113364 614 113416 620
rect 115216 610 115244 1838
rect 115584 1465 115612 1838
rect 115664 1828 115716 1834
rect 115664 1770 115716 1776
rect 115676 1494 115704 1770
rect 115664 1488 115716 1494
rect 115570 1456 115626 1465
rect 115664 1430 115716 1436
rect 115570 1391 115626 1400
rect 115860 1358 115888 9318
rect 116044 6338 116072 9386
rect 116492 8832 116544 8838
rect 116492 8774 116544 8780
rect 116308 7404 116360 7410
rect 116308 7346 116360 7352
rect 116216 6792 116268 6798
rect 116214 6760 116216 6769
rect 116268 6760 116270 6769
rect 116214 6695 116270 6704
rect 115952 6322 116072 6338
rect 115940 6316 116072 6322
rect 115992 6310 116072 6316
rect 115940 6258 115992 6264
rect 116124 6248 116176 6254
rect 116124 6190 116176 6196
rect 115938 6080 115994 6089
rect 115938 6015 115994 6024
rect 115952 1970 115980 6015
rect 116032 5908 116084 5914
rect 116032 5850 116084 5856
rect 116044 5574 116072 5850
rect 116032 5568 116084 5574
rect 116032 5510 116084 5516
rect 116030 5264 116086 5273
rect 116030 5199 116086 5208
rect 116044 5166 116072 5199
rect 116032 5160 116084 5166
rect 116032 5102 116084 5108
rect 116032 5024 116084 5030
rect 116032 4966 116084 4972
rect 116044 4729 116072 4966
rect 116030 4720 116086 4729
rect 116030 4655 116086 4664
rect 116136 2854 116164 6190
rect 116216 6112 116268 6118
rect 116216 6054 116268 6060
rect 116228 5234 116256 6054
rect 116216 5228 116268 5234
rect 116216 5170 116268 5176
rect 116320 5030 116348 7346
rect 116400 7200 116452 7206
rect 116400 7142 116452 7148
rect 116412 6254 116440 7142
rect 116400 6248 116452 6254
rect 116400 6190 116452 6196
rect 116400 6112 116452 6118
rect 116504 6089 116532 8774
rect 116860 8084 116912 8090
rect 116860 8026 116912 8032
rect 116584 7472 116636 7478
rect 116584 7414 116636 7420
rect 116596 7206 116624 7414
rect 116768 7404 116820 7410
rect 116768 7346 116820 7352
rect 116584 7200 116636 7206
rect 116584 7142 116636 7148
rect 116584 6928 116636 6934
rect 116582 6896 116584 6905
rect 116636 6896 116638 6905
rect 116582 6831 116638 6840
rect 116676 6656 116728 6662
rect 116676 6598 116728 6604
rect 116584 6248 116636 6254
rect 116584 6190 116636 6196
rect 116400 6054 116452 6060
rect 116490 6080 116546 6089
rect 116412 5817 116440 6054
rect 116490 6015 116546 6024
rect 116490 5944 116546 5953
rect 116596 5914 116624 6190
rect 116490 5879 116546 5888
rect 116584 5908 116636 5914
rect 116398 5808 116454 5817
rect 116504 5778 116532 5879
rect 116584 5850 116636 5856
rect 116398 5743 116454 5752
rect 116492 5772 116544 5778
rect 116412 5710 116440 5743
rect 116492 5714 116544 5720
rect 116400 5704 116452 5710
rect 116400 5646 116452 5652
rect 116688 5166 116716 6598
rect 116780 5914 116808 7346
rect 116872 6934 116900 8026
rect 116950 7984 117006 7993
rect 116950 7919 117006 7928
rect 116860 6928 116912 6934
rect 116860 6870 116912 6876
rect 116860 6724 116912 6730
rect 116860 6666 116912 6672
rect 116872 6458 116900 6666
rect 116860 6452 116912 6458
rect 116860 6394 116912 6400
rect 116872 6254 116900 6394
rect 116860 6248 116912 6254
rect 116860 6190 116912 6196
rect 116768 5908 116820 5914
rect 116768 5850 116820 5856
rect 116964 5234 116992 7919
rect 116952 5228 117004 5234
rect 116952 5170 117004 5176
rect 116676 5160 116728 5166
rect 116676 5102 116728 5108
rect 116308 5024 116360 5030
rect 116308 4966 116360 4972
rect 116320 4758 116348 4966
rect 116308 4752 116360 4758
rect 116308 4694 116360 4700
rect 116124 2848 116176 2854
rect 116124 2790 116176 2796
rect 116032 2304 116084 2310
rect 116032 2246 116084 2252
rect 116044 1970 116072 2246
rect 115940 1964 115992 1970
rect 115940 1906 115992 1912
rect 116032 1964 116084 1970
rect 116032 1906 116084 1912
rect 116216 1964 116268 1970
rect 116320 1952 116348 4694
rect 116688 4214 116716 5102
rect 116676 4208 116728 4214
rect 116676 4150 116728 4156
rect 117056 4146 117084 9862
rect 117240 8974 117268 10231
rect 117320 9648 117372 9654
rect 117320 9590 117372 9596
rect 117228 8968 117280 8974
rect 117228 8910 117280 8916
rect 117136 7200 117188 7206
rect 117136 7142 117188 7148
rect 117148 5030 117176 7142
rect 117332 6202 117360 9590
rect 118068 9586 118096 10231
rect 118712 9586 118740 10231
rect 119356 9586 119384 10231
rect 120368 9586 120396 10231
rect 121104 9586 121132 10231
rect 121644 9920 121696 9926
rect 121644 9862 121696 9868
rect 121656 9722 121684 9862
rect 121748 9722 121776 10231
rect 121644 9716 121696 9722
rect 121644 9658 121696 9664
rect 121736 9716 121788 9722
rect 121736 9658 121788 9664
rect 118056 9580 118108 9586
rect 118056 9522 118108 9528
rect 118700 9580 118752 9586
rect 118700 9522 118752 9528
rect 119344 9580 119396 9586
rect 119344 9522 119396 9528
rect 120356 9580 120408 9586
rect 120356 9522 120408 9528
rect 121092 9580 121144 9586
rect 121092 9522 121144 9528
rect 121644 9580 121696 9586
rect 121644 9522 121696 9528
rect 121552 9444 121604 9450
rect 121552 9386 121604 9392
rect 117964 9376 118016 9382
rect 117964 9318 118016 9324
rect 118332 9376 118384 9382
rect 118332 9318 118384 9324
rect 119160 9376 119212 9382
rect 119160 9318 119212 9324
rect 120908 9376 120960 9382
rect 120908 9318 120960 9324
rect 117872 8016 117924 8022
rect 117872 7958 117924 7964
rect 117504 7880 117556 7886
rect 117504 7822 117556 7828
rect 117516 7546 117544 7822
rect 117504 7540 117556 7546
rect 117504 7482 117556 7488
rect 117516 6746 117544 7482
rect 117688 7336 117740 7342
rect 117688 7278 117740 7284
rect 117240 6174 117360 6202
rect 117424 6718 117544 6746
rect 117136 5024 117188 5030
rect 117136 4966 117188 4972
rect 117240 4434 117268 6174
rect 117320 6112 117372 6118
rect 117320 6054 117372 6060
rect 117332 5778 117360 6054
rect 117320 5772 117372 5778
rect 117320 5714 117372 5720
rect 117320 5364 117372 5370
rect 117320 5306 117372 5312
rect 117332 4622 117360 5306
rect 117424 5166 117452 6718
rect 117596 6656 117648 6662
rect 117516 6604 117596 6610
rect 117516 6598 117648 6604
rect 117516 6582 117636 6598
rect 117516 5642 117544 6582
rect 117700 6304 117728 7278
rect 117780 6724 117832 6730
rect 117780 6666 117832 6672
rect 117608 6276 117728 6304
rect 117608 5930 117636 6276
rect 117608 5902 117728 5930
rect 117596 5772 117648 5778
rect 117596 5714 117648 5720
rect 117504 5636 117556 5642
rect 117504 5578 117556 5584
rect 117516 5302 117544 5578
rect 117608 5574 117636 5714
rect 117596 5568 117648 5574
rect 117596 5510 117648 5516
rect 117504 5296 117556 5302
rect 117596 5296 117648 5302
rect 117504 5238 117556 5244
rect 117594 5264 117596 5273
rect 117648 5264 117650 5273
rect 117594 5199 117650 5208
rect 117412 5160 117464 5166
rect 117412 5102 117464 5108
rect 117424 4826 117452 5102
rect 117412 4820 117464 4826
rect 117412 4762 117464 4768
rect 117320 4616 117372 4622
rect 117320 4558 117372 4564
rect 117240 4406 117360 4434
rect 117044 4140 117096 4146
rect 117044 4082 117096 4088
rect 117228 4072 117280 4078
rect 117228 4014 117280 4020
rect 117240 3369 117268 4014
rect 117332 3534 117360 4406
rect 117412 3664 117464 3670
rect 117412 3606 117464 3612
rect 117320 3528 117372 3534
rect 117320 3470 117372 3476
rect 117226 3360 117282 3369
rect 117226 3295 117282 3304
rect 117226 2816 117282 2825
rect 117282 2774 117360 2802
rect 117226 2751 117282 2760
rect 117332 2582 117360 2774
rect 117320 2576 117372 2582
rect 117320 2518 117372 2524
rect 117228 2440 117280 2446
rect 117228 2382 117280 2388
rect 117320 2440 117372 2446
rect 117320 2382 117372 2388
rect 117240 2038 117268 2382
rect 117136 2032 117188 2038
rect 117136 1974 117188 1980
rect 117228 2032 117280 2038
rect 117228 1974 117280 1980
rect 116268 1924 116348 1952
rect 116216 1906 116268 1912
rect 115848 1352 115900 1358
rect 115848 1294 115900 1300
rect 116124 1352 116176 1358
rect 116228 1340 116256 1906
rect 117148 1494 117176 1974
rect 117136 1488 117188 1494
rect 117332 1465 117360 2382
rect 117424 1970 117452 3606
rect 117700 3602 117728 5902
rect 117792 4672 117820 6666
rect 117884 6458 117912 7958
rect 117872 6452 117924 6458
rect 117872 6394 117924 6400
rect 117870 6352 117926 6361
rect 117870 6287 117926 6296
rect 117884 6254 117912 6287
rect 117872 6248 117924 6254
rect 117872 6190 117924 6196
rect 117884 5953 117912 6190
rect 117870 5944 117926 5953
rect 117870 5879 117926 5888
rect 117872 4684 117924 4690
rect 117792 4644 117872 4672
rect 117872 4626 117924 4632
rect 117976 4078 118004 9318
rect 118056 7404 118108 7410
rect 118056 7346 118108 7352
rect 118068 6662 118096 7346
rect 118148 7200 118200 7206
rect 118148 7142 118200 7148
rect 118160 6882 118188 7142
rect 118160 6866 118280 6882
rect 118148 6860 118280 6866
rect 118200 6854 118280 6860
rect 118148 6802 118200 6808
rect 118148 6724 118200 6730
rect 118148 6666 118200 6672
rect 118056 6656 118108 6662
rect 118056 6598 118108 6604
rect 118160 6458 118188 6666
rect 118252 6458 118280 6854
rect 118056 6452 118108 6458
rect 118056 6394 118108 6400
rect 118148 6452 118200 6458
rect 118148 6394 118200 6400
rect 118240 6452 118292 6458
rect 118240 6394 118292 6400
rect 118068 4758 118096 6394
rect 118146 6216 118202 6225
rect 118146 6151 118202 6160
rect 118160 6118 118188 6151
rect 118148 6112 118200 6118
rect 118148 6054 118200 6060
rect 118252 5642 118280 6394
rect 118240 5636 118292 5642
rect 118240 5578 118292 5584
rect 118148 5024 118200 5030
rect 118148 4966 118200 4972
rect 118056 4752 118108 4758
rect 118056 4694 118108 4700
rect 118160 4128 118188 4966
rect 118240 4480 118292 4486
rect 118240 4422 118292 4428
rect 118252 4282 118280 4422
rect 118240 4276 118292 4282
rect 118240 4218 118292 4224
rect 118240 4140 118292 4146
rect 118160 4100 118240 4128
rect 118240 4082 118292 4088
rect 117964 4072 118016 4078
rect 117964 4014 118016 4020
rect 118056 4072 118108 4078
rect 118056 4014 118108 4020
rect 117688 3596 117740 3602
rect 117688 3538 117740 3544
rect 117872 3528 117924 3534
rect 117872 3470 117924 3476
rect 117504 2984 117556 2990
rect 117504 2926 117556 2932
rect 117412 1964 117464 1970
rect 117412 1906 117464 1912
rect 117424 1562 117452 1906
rect 117412 1556 117464 1562
rect 117412 1498 117464 1504
rect 117136 1430 117188 1436
rect 117318 1456 117374 1465
rect 117318 1391 117374 1400
rect 117516 1358 117544 2926
rect 117884 2774 117912 3470
rect 118068 2774 118096 4014
rect 118148 3664 118200 3670
rect 118148 3606 118200 3612
rect 117792 2746 117912 2774
rect 117976 2746 118096 2774
rect 117596 2304 117648 2310
rect 117596 2246 117648 2252
rect 116176 1312 116256 1340
rect 117504 1352 117556 1358
rect 116124 1294 116176 1300
rect 117504 1294 117556 1300
rect 117608 1290 117636 2246
rect 117686 2000 117742 2009
rect 117686 1935 117688 1944
rect 117740 1935 117742 1944
rect 117688 1906 117740 1912
rect 117596 1284 117648 1290
rect 117596 1226 117648 1232
rect 115204 604 115256 610
rect 115204 546 115256 552
rect 117792 513 117820 2746
rect 117976 1222 118004 2746
rect 118056 2304 118108 2310
rect 118056 2246 118108 2252
rect 118068 1442 118096 2246
rect 118160 1902 118188 3606
rect 118148 1896 118200 1902
rect 118148 1838 118200 1844
rect 118148 1760 118200 1766
rect 118344 1714 118372 9318
rect 118516 7472 118568 7478
rect 118516 7414 118568 7420
rect 118424 6792 118476 6798
rect 118424 6734 118476 6740
rect 118436 6254 118464 6734
rect 118424 6248 118476 6254
rect 118424 6190 118476 6196
rect 118424 4684 118476 4690
rect 118424 4626 118476 4632
rect 118436 3670 118464 4626
rect 118528 4622 118556 7414
rect 118608 7268 118660 7274
rect 118608 7210 118660 7216
rect 118620 7002 118648 7210
rect 118608 6996 118660 7002
rect 118608 6938 118660 6944
rect 118882 6760 118938 6769
rect 118882 6695 118938 6704
rect 118896 6322 118924 6695
rect 118884 6316 118936 6322
rect 118884 6258 118936 6264
rect 118700 6248 118752 6254
rect 118700 6190 118752 6196
rect 119068 6248 119120 6254
rect 119068 6190 119120 6196
rect 118712 5574 118740 6190
rect 119080 5778 119108 6190
rect 119068 5772 119120 5778
rect 119068 5714 119120 5720
rect 118700 5568 118752 5574
rect 118700 5510 118752 5516
rect 118976 4820 119028 4826
rect 118976 4762 119028 4768
rect 118700 4752 118752 4758
rect 118700 4694 118752 4700
rect 118516 4616 118568 4622
rect 118516 4558 118568 4564
rect 118424 3664 118476 3670
rect 118424 3606 118476 3612
rect 118516 3596 118568 3602
rect 118516 3538 118568 3544
rect 118528 1986 118556 3538
rect 118608 2984 118660 2990
rect 118608 2926 118660 2932
rect 118200 1708 118372 1714
rect 118148 1702 118372 1708
rect 118160 1686 118372 1702
rect 118436 1958 118556 1986
rect 118068 1414 118188 1442
rect 118056 1352 118108 1358
rect 118056 1294 118108 1300
rect 117964 1216 118016 1222
rect 117964 1158 118016 1164
rect 118068 513 118096 1294
rect 118160 1018 118188 1414
rect 118436 1290 118464 1958
rect 118516 1896 118568 1902
rect 118516 1838 118568 1844
rect 118528 1562 118556 1838
rect 118620 1766 118648 2926
rect 118712 2514 118740 4694
rect 118988 3534 119016 4762
rect 119172 3602 119200 9318
rect 120816 8424 120868 8430
rect 120816 8366 120868 8372
rect 120262 7848 120318 7857
rect 120262 7783 120318 7792
rect 120080 7404 120132 7410
rect 120080 7346 120132 7352
rect 119436 7200 119488 7206
rect 119250 7168 119306 7177
rect 119436 7142 119488 7148
rect 119250 7103 119306 7112
rect 119264 5710 119292 7103
rect 119252 5704 119304 5710
rect 119252 5646 119304 5652
rect 119264 5234 119292 5646
rect 119252 5228 119304 5234
rect 119252 5170 119304 5176
rect 119448 4622 119476 7142
rect 119986 6896 120042 6905
rect 119986 6831 120042 6840
rect 120000 6662 120028 6831
rect 119988 6656 120040 6662
rect 119988 6598 120040 6604
rect 119896 6112 119948 6118
rect 119896 6054 119948 6060
rect 119908 5642 119936 6054
rect 119896 5636 119948 5642
rect 119896 5578 119948 5584
rect 120000 5234 120028 6598
rect 120092 6458 120120 7346
rect 120080 6452 120132 6458
rect 120080 6394 120132 6400
rect 119988 5228 120040 5234
rect 119988 5170 120040 5176
rect 120172 5092 120224 5098
rect 120172 5034 120224 5040
rect 119436 4616 119488 4622
rect 119436 4558 119488 4564
rect 119160 3596 119212 3602
rect 119160 3538 119212 3544
rect 118884 3528 118936 3534
rect 118884 3470 118936 3476
rect 118976 3528 119028 3534
rect 118976 3470 119028 3476
rect 118700 2508 118752 2514
rect 118700 2450 118752 2456
rect 118608 1760 118660 1766
rect 118608 1702 118660 1708
rect 118516 1556 118568 1562
rect 118516 1498 118568 1504
rect 118700 1352 118752 1358
rect 118700 1294 118752 1300
rect 118424 1284 118476 1290
rect 118424 1226 118476 1232
rect 118148 1012 118200 1018
rect 118148 954 118200 960
rect 118712 513 118740 1294
rect 118896 1222 118924 3470
rect 118988 2990 119016 3470
rect 119252 3392 119304 3398
rect 119252 3334 119304 3340
rect 119264 3058 119292 3334
rect 119252 3052 119304 3058
rect 119252 2994 119304 3000
rect 118976 2984 119028 2990
rect 119028 2944 119108 2972
rect 118976 2926 119028 2932
rect 118976 2440 119028 2446
rect 118976 2382 119028 2388
rect 118988 2106 119016 2382
rect 118976 2100 119028 2106
rect 118976 2042 119028 2048
rect 119080 1902 119108 2944
rect 119448 2553 119476 4558
rect 120080 4548 120132 4554
rect 120080 4490 120132 4496
rect 119988 4480 120040 4486
rect 119988 4422 120040 4428
rect 120000 3058 120028 4422
rect 120092 4214 120120 4490
rect 120080 4208 120132 4214
rect 120080 4150 120132 4156
rect 120080 3936 120132 3942
rect 120080 3878 120132 3884
rect 120092 3602 120120 3878
rect 120080 3596 120132 3602
rect 120080 3538 120132 3544
rect 119988 3052 120040 3058
rect 119988 2994 120040 3000
rect 120080 2848 120132 2854
rect 120080 2790 120132 2796
rect 119434 2544 119490 2553
rect 119434 2479 119490 2488
rect 119068 1896 119120 1902
rect 119068 1838 119120 1844
rect 120092 1562 120120 2790
rect 120184 1970 120212 5034
rect 120276 4010 120304 7783
rect 120540 6180 120592 6186
rect 120540 6122 120592 6128
rect 120552 5642 120580 6122
rect 120540 5636 120592 5642
rect 120724 5636 120776 5642
rect 120592 5596 120724 5624
rect 120540 5578 120592 5584
rect 120724 5578 120776 5584
rect 120448 4548 120500 4554
rect 120448 4490 120500 4496
rect 120460 4146 120488 4490
rect 120448 4140 120500 4146
rect 120448 4082 120500 4088
rect 120264 4004 120316 4010
rect 120264 3946 120316 3952
rect 120276 2514 120304 3946
rect 120724 2984 120776 2990
rect 120724 2926 120776 2932
rect 120264 2508 120316 2514
rect 120264 2450 120316 2456
rect 120736 2106 120764 2926
rect 120828 2689 120856 8366
rect 120920 7954 120948 9318
rect 121000 9172 121052 9178
rect 121000 9114 121052 9120
rect 121012 8974 121040 9114
rect 121000 8968 121052 8974
rect 121000 8910 121052 8916
rect 120908 7948 120960 7954
rect 120908 7890 120960 7896
rect 121012 7546 121040 8910
rect 121564 8634 121592 9386
rect 121656 8634 121684 9522
rect 121828 9104 121880 9110
rect 121828 9046 121880 9052
rect 121840 8906 121868 9046
rect 121828 8900 121880 8906
rect 121828 8842 121880 8848
rect 121736 8832 121788 8838
rect 121736 8774 121788 8780
rect 121552 8628 121604 8634
rect 121552 8570 121604 8576
rect 121644 8628 121696 8634
rect 121644 8570 121696 8576
rect 121000 7540 121052 7546
rect 121000 7482 121052 7488
rect 121644 5840 121696 5846
rect 121472 5788 121644 5794
rect 121472 5782 121696 5788
rect 121472 5778 121684 5782
rect 121460 5772 121684 5778
rect 121512 5766 121684 5772
rect 121460 5714 121512 5720
rect 121184 5568 121236 5574
rect 121184 5510 121236 5516
rect 121000 5228 121052 5234
rect 121000 5170 121052 5176
rect 120908 5024 120960 5030
rect 120908 4966 120960 4972
rect 120920 4826 120948 4966
rect 120908 4820 120960 4826
rect 120908 4762 120960 4768
rect 120920 3942 120948 4762
rect 121012 4690 121040 5170
rect 121000 4684 121052 4690
rect 121000 4626 121052 4632
rect 121012 4146 121040 4626
rect 121000 4140 121052 4146
rect 121000 4082 121052 4088
rect 120908 3936 120960 3942
rect 120908 3878 120960 3884
rect 120920 3670 120948 3878
rect 120908 3664 120960 3670
rect 120908 3606 120960 3612
rect 120814 2680 120870 2689
rect 120814 2615 120870 2624
rect 121090 2680 121146 2689
rect 121090 2615 121146 2624
rect 121104 2106 121132 2615
rect 121196 2446 121224 5510
rect 121276 5160 121328 5166
rect 121276 5102 121328 5108
rect 121288 4622 121316 5102
rect 121644 5024 121696 5030
rect 121644 4966 121696 4972
rect 121366 4720 121422 4729
rect 121366 4655 121422 4664
rect 121276 4616 121328 4622
rect 121276 4558 121328 4564
rect 121380 4554 121408 4655
rect 121368 4548 121420 4554
rect 121368 4490 121420 4496
rect 121460 4072 121512 4078
rect 121460 4014 121512 4020
rect 121472 3738 121500 4014
rect 121460 3732 121512 3738
rect 121460 3674 121512 3680
rect 121656 2990 121684 4966
rect 121748 4706 121776 8774
rect 121840 8498 121868 8842
rect 122196 8832 122248 8838
rect 122196 8774 122248 8780
rect 122208 8498 122236 8774
rect 122392 8634 122420 10231
rect 122656 8968 122708 8974
rect 122852 8922 122880 10406
rect 123206 10296 123262 10305
rect 123206 10231 123262 10240
rect 124034 10296 124090 10305
rect 124034 10231 124090 10240
rect 122708 8916 122880 8922
rect 122656 8910 122880 8916
rect 122668 8906 122880 8910
rect 122668 8900 122892 8906
rect 122668 8894 122840 8900
rect 122840 8842 122892 8848
rect 122380 8628 122432 8634
rect 122380 8570 122432 8576
rect 121828 8492 121880 8498
rect 121828 8434 121880 8440
rect 122196 8492 122248 8498
rect 122196 8434 122248 8440
rect 122102 7440 122158 7449
rect 122102 7375 122158 7384
rect 121918 6080 121974 6089
rect 121918 6015 121974 6024
rect 121932 5710 121960 6015
rect 121920 5704 121972 5710
rect 121918 5672 121920 5681
rect 121972 5672 121974 5681
rect 121918 5607 121974 5616
rect 121828 5228 121880 5234
rect 121828 5170 121880 5176
rect 121920 5228 121972 5234
rect 121920 5170 121972 5176
rect 121840 4826 121868 5170
rect 121828 4820 121880 4826
rect 121828 4762 121880 4768
rect 121748 4678 121868 4706
rect 121644 2984 121696 2990
rect 121644 2926 121696 2932
rect 121736 2916 121788 2922
rect 121736 2858 121788 2864
rect 121184 2440 121236 2446
rect 121184 2382 121236 2388
rect 120724 2100 120776 2106
rect 120724 2042 120776 2048
rect 121092 2100 121144 2106
rect 121092 2042 121144 2048
rect 121748 2038 121776 2858
rect 121736 2032 121788 2038
rect 121736 1974 121788 1980
rect 120172 1964 120224 1970
rect 120172 1906 120224 1912
rect 120724 1964 120776 1970
rect 120724 1906 120776 1912
rect 121460 1964 121512 1970
rect 121460 1906 121512 1912
rect 120540 1760 120592 1766
rect 120540 1702 120592 1708
rect 120080 1556 120132 1562
rect 120080 1498 120132 1504
rect 119344 1352 119396 1358
rect 119344 1294 119396 1300
rect 120356 1352 120408 1358
rect 120356 1294 120408 1300
rect 118884 1216 118936 1222
rect 118884 1158 118936 1164
rect 119356 513 119384 1294
rect 120368 513 120396 1294
rect 120552 1018 120580 1702
rect 120736 1494 120764 1906
rect 120724 1488 120776 1494
rect 120724 1430 120776 1436
rect 121092 1352 121144 1358
rect 121092 1294 121144 1300
rect 120540 1012 120592 1018
rect 120540 954 120592 960
rect 121104 513 121132 1294
rect 121472 882 121500 1906
rect 121840 1873 121868 4678
rect 121932 4010 121960 5170
rect 122116 4214 122144 7375
rect 122472 5364 122524 5370
rect 122472 5306 122524 5312
rect 122380 5092 122432 5098
rect 122380 5034 122432 5040
rect 122288 5024 122340 5030
rect 122288 4966 122340 4972
rect 122104 4208 122156 4214
rect 122104 4150 122156 4156
rect 121920 4004 121972 4010
rect 121920 3946 121972 3952
rect 122012 4004 122064 4010
rect 122012 3946 122064 3952
rect 122024 2774 122052 3946
rect 122116 3534 122144 4150
rect 122300 3602 122328 4966
rect 122392 4486 122420 5034
rect 122484 4622 122512 5306
rect 122748 5160 122800 5166
rect 122748 5102 122800 5108
rect 122760 4690 122788 5102
rect 122748 4684 122800 4690
rect 122748 4626 122800 4632
rect 122472 4616 122524 4622
rect 122472 4558 122524 4564
rect 122380 4480 122432 4486
rect 122380 4422 122432 4428
rect 122472 4072 122524 4078
rect 122472 4014 122524 4020
rect 122484 3738 122512 4014
rect 122472 3732 122524 3738
rect 122472 3674 122524 3680
rect 122288 3596 122340 3602
rect 122288 3538 122340 3544
rect 122104 3528 122156 3534
rect 122104 3470 122156 3476
rect 121932 2746 122052 2774
rect 121932 2514 121960 2746
rect 121920 2508 121972 2514
rect 121920 2450 121972 2456
rect 122656 2304 122708 2310
rect 122656 2246 122708 2252
rect 122668 1970 122696 2246
rect 122656 1964 122708 1970
rect 122656 1906 122708 1912
rect 122852 1902 122880 8842
rect 123024 8832 123076 8838
rect 123024 8774 123076 8780
rect 123036 8498 123064 8774
rect 123220 8634 123248 10231
rect 123300 9648 123352 9654
rect 123300 9590 123352 9596
rect 123312 9042 123340 9590
rect 123300 9036 123352 9042
rect 123300 8978 123352 8984
rect 123484 9036 123536 9042
rect 123484 8978 123536 8984
rect 123392 8900 123444 8906
rect 123392 8842 123444 8848
rect 123208 8628 123260 8634
rect 123208 8570 123260 8576
rect 123404 8566 123432 8842
rect 123392 8560 123444 8566
rect 123392 8502 123444 8508
rect 123024 8492 123076 8498
rect 123024 8434 123076 8440
rect 123024 4480 123076 4486
rect 123024 4422 123076 4428
rect 123036 3534 123064 4422
rect 123024 3528 123076 3534
rect 123024 3470 123076 3476
rect 123496 2145 123524 8978
rect 123852 8832 123904 8838
rect 123852 8774 123904 8780
rect 123864 8498 123892 8774
rect 124048 8634 124076 10231
rect 124128 8968 124180 8974
rect 124232 8922 124260 10474
rect 124692 10130 124720 10474
rect 125598 10432 125654 10441
rect 125598 10367 125654 10376
rect 125230 10296 125286 10305
rect 125230 10231 125286 10240
rect 124680 10124 124732 10130
rect 124680 10066 124732 10072
rect 124404 9580 124456 9586
rect 124404 9522 124456 9528
rect 124416 9178 124444 9522
rect 124692 9178 124720 10066
rect 125244 9722 125272 10231
rect 125232 9716 125284 9722
rect 125232 9658 125284 9664
rect 124404 9172 124456 9178
rect 124404 9114 124456 9120
rect 124680 9172 124732 9178
rect 124680 9114 124732 9120
rect 124692 8974 124720 9114
rect 124180 8916 124260 8922
rect 124128 8910 124260 8916
rect 124680 8968 124732 8974
rect 124680 8910 124732 8916
rect 125048 8968 125100 8974
rect 125048 8910 125100 8916
rect 124140 8894 124260 8910
rect 124036 8628 124088 8634
rect 124036 8570 124088 8576
rect 123852 8492 123904 8498
rect 123852 8434 123904 8440
rect 124232 7410 124260 8894
rect 124220 7404 124272 7410
rect 124220 7346 124272 7352
rect 124772 7404 124824 7410
rect 124772 7346 124824 7352
rect 124126 2816 124182 2825
rect 124182 2774 124260 2802
rect 124126 2751 124182 2760
rect 124126 2680 124182 2689
rect 124232 2650 124260 2774
rect 124126 2615 124182 2624
rect 124220 2644 124272 2650
rect 124140 2145 124168 2615
rect 124220 2586 124272 2592
rect 124784 2514 124812 7346
rect 124772 2508 124824 2514
rect 124772 2450 124824 2456
rect 124312 2440 124364 2446
rect 124312 2382 124364 2388
rect 124956 2440 125008 2446
rect 124956 2382 125008 2388
rect 123482 2136 123538 2145
rect 124126 2136 124182 2145
rect 123482 2071 123538 2080
rect 124048 2094 124126 2122
rect 124048 1902 124076 2094
rect 124324 2106 124352 2382
rect 124126 2071 124182 2080
rect 124312 2100 124364 2106
rect 124312 2042 124364 2048
rect 124968 1970 124996 2382
rect 125060 1970 125088 8910
rect 125416 8832 125468 8838
rect 125416 8774 125468 8780
rect 125428 8498 125456 8774
rect 125612 8634 125640 10367
rect 125888 10130 125916 10678
rect 127624 10668 127676 10674
rect 127624 10610 127676 10616
rect 131120 10668 131172 10674
rect 131120 10610 131172 10616
rect 131856 10668 131908 10674
rect 131856 10610 131908 10616
rect 126704 10396 126756 10402
rect 126704 10338 126756 10344
rect 126334 10296 126390 10305
rect 126334 10231 126390 10240
rect 125876 10124 125928 10130
rect 125876 10066 125928 10072
rect 125888 8974 125916 10066
rect 126348 9722 126376 10231
rect 126716 10198 126744 10338
rect 126978 10296 127034 10305
rect 126978 10231 127034 10240
rect 126704 10192 126756 10198
rect 126704 10134 126756 10140
rect 126336 9716 126388 9722
rect 126336 9658 126388 9664
rect 126244 9580 126296 9586
rect 126244 9522 126296 9528
rect 126256 9178 126284 9522
rect 126244 9172 126296 9178
rect 126244 9114 126296 9120
rect 126716 8974 126744 10134
rect 125876 8968 125928 8974
rect 125876 8910 125928 8916
rect 126336 8968 126388 8974
rect 126336 8910 126388 8916
rect 126704 8968 126756 8974
rect 126704 8910 126756 8916
rect 125600 8628 125652 8634
rect 125600 8570 125652 8576
rect 125416 8492 125468 8498
rect 125416 8434 125468 8440
rect 125888 2774 125916 8910
rect 125888 2746 126192 2774
rect 126060 2440 126112 2446
rect 126060 2382 126112 2388
rect 125140 2304 125192 2310
rect 125140 2246 125192 2252
rect 124956 1964 125008 1970
rect 124956 1906 125008 1912
rect 125048 1964 125100 1970
rect 125048 1906 125100 1912
rect 122104 1896 122156 1902
rect 121826 1864 121882 1873
rect 121826 1799 121882 1808
rect 122102 1864 122104 1873
rect 122840 1896 122892 1902
rect 122156 1864 122158 1873
rect 122840 1838 122892 1844
rect 123116 1896 123168 1902
rect 123116 1838 123168 1844
rect 124036 1896 124088 1902
rect 124036 1838 124088 1844
rect 122102 1799 122158 1808
rect 121644 1760 121696 1766
rect 121644 1702 121696 1708
rect 122472 1760 122524 1766
rect 122472 1702 122524 1708
rect 121656 1358 121684 1702
rect 122484 1358 122512 1702
rect 123128 1494 123156 1838
rect 123208 1760 123260 1766
rect 123208 1702 123260 1708
rect 123116 1488 123168 1494
rect 123116 1430 123168 1436
rect 123220 1358 123248 1702
rect 125152 1358 125180 2246
rect 125784 1760 125836 1766
rect 125784 1702 125836 1708
rect 125796 1358 125824 1702
rect 126072 1562 126100 2382
rect 126060 1556 126112 1562
rect 126060 1498 126112 1504
rect 126164 1426 126192 2746
rect 126244 2304 126296 2310
rect 126244 2246 126296 2252
rect 126152 1420 126204 1426
rect 126152 1362 126204 1368
rect 121644 1352 121696 1358
rect 121644 1294 121696 1300
rect 122472 1352 122524 1358
rect 122472 1294 122524 1300
rect 123208 1352 123260 1358
rect 123208 1294 123260 1300
rect 125140 1352 125192 1358
rect 125140 1294 125192 1300
rect 125784 1352 125836 1358
rect 125784 1294 125836 1300
rect 121828 1216 121880 1222
rect 121828 1158 121880 1164
rect 122656 1216 122708 1222
rect 122656 1158 122708 1164
rect 123392 1216 123444 1222
rect 123392 1158 123444 1164
rect 124404 1216 124456 1222
rect 124404 1158 124456 1164
rect 125324 1216 125376 1222
rect 125324 1158 125376 1164
rect 121460 876 121512 882
rect 121460 818 121512 824
rect 121840 513 121868 1158
rect 122668 513 122696 1158
rect 123404 513 123432 1158
rect 124416 649 124444 1158
rect 125336 649 125364 1158
rect 126256 649 126284 2246
rect 126348 1970 126376 8910
rect 126796 8832 126848 8838
rect 126796 8774 126848 8780
rect 126808 8498 126836 8774
rect 126992 8634 127020 10231
rect 127636 9178 127664 10610
rect 127714 10296 127770 10305
rect 127714 10231 127770 10240
rect 128266 10296 128322 10305
rect 128266 10231 128322 10240
rect 129278 10296 129334 10305
rect 129278 10231 129334 10240
rect 129646 10296 129702 10305
rect 129646 10231 129702 10240
rect 130750 10296 130806 10305
rect 131132 10266 131160 10610
rect 131486 10296 131542 10305
rect 130750 10231 130806 10240
rect 131120 10260 131172 10266
rect 127624 9172 127676 9178
rect 127624 9114 127676 9120
rect 127636 8974 127664 9114
rect 127624 8968 127676 8974
rect 127624 8910 127676 8916
rect 127532 8832 127584 8838
rect 127532 8774 127584 8780
rect 126980 8628 127032 8634
rect 126980 8570 127032 8576
rect 127544 8498 127572 8774
rect 126796 8492 126848 8498
rect 126796 8434 126848 8440
rect 127532 8492 127584 8498
rect 127532 8434 127584 8440
rect 127636 2774 127664 8910
rect 127728 8634 127756 10231
rect 127992 9512 128044 9518
rect 127992 9454 128044 9460
rect 127808 8968 127860 8974
rect 127808 8910 127860 8916
rect 127716 8628 127768 8634
rect 127716 8570 127768 8576
rect 127820 8566 127848 8910
rect 127808 8560 127860 8566
rect 127808 8502 127860 8508
rect 127714 6216 127770 6225
rect 127714 6151 127770 6160
rect 127728 5710 127756 6151
rect 127716 5704 127768 5710
rect 127716 5646 127768 5652
rect 127452 2746 127664 2774
rect 126704 2440 126756 2446
rect 126704 2382 126756 2388
rect 126716 2106 126744 2382
rect 126980 2304 127032 2310
rect 126980 2246 127032 2252
rect 126704 2100 126756 2106
rect 126704 2042 126756 2048
rect 126336 1964 126388 1970
rect 126336 1906 126388 1912
rect 126428 1896 126480 1902
rect 126428 1838 126480 1844
rect 126440 1358 126468 1838
rect 126992 1465 127020 2246
rect 127452 1902 127480 2746
rect 128004 1970 128032 9454
rect 128084 9376 128136 9382
rect 128084 9318 128136 9324
rect 128096 8498 128124 9318
rect 128280 8634 128308 10231
rect 128820 9580 128872 9586
rect 128820 9522 128872 9528
rect 128728 9376 128780 9382
rect 128728 9318 128780 9324
rect 128740 9178 128768 9318
rect 128728 9172 128780 9178
rect 128728 9114 128780 9120
rect 128832 9042 128860 9522
rect 128820 9036 128872 9042
rect 128820 8978 128872 8984
rect 128268 8628 128320 8634
rect 128268 8570 128320 8576
rect 128832 8498 128860 8978
rect 128084 8492 128136 8498
rect 128084 8434 128136 8440
rect 128820 8492 128872 8498
rect 128820 8434 128872 8440
rect 128912 8424 128964 8430
rect 128912 8366 128964 8372
rect 128084 6656 128136 6662
rect 128084 6598 128136 6604
rect 128096 5710 128124 6598
rect 128084 5704 128136 5710
rect 128084 5646 128136 5652
rect 128360 2440 128412 2446
rect 128360 2382 128412 2388
rect 128372 2106 128400 2382
rect 128820 2372 128872 2378
rect 128820 2314 128872 2320
rect 128452 2304 128504 2310
rect 128452 2246 128504 2252
rect 128360 2100 128412 2106
rect 128360 2042 128412 2048
rect 127992 1964 128044 1970
rect 127992 1906 128044 1912
rect 127440 1896 127492 1902
rect 127440 1838 127492 1844
rect 127624 1760 127676 1766
rect 127624 1702 127676 1708
rect 126978 1456 127034 1465
rect 126978 1391 127034 1400
rect 127636 1358 127664 1702
rect 128464 1465 128492 2246
rect 128832 1970 128860 2314
rect 128820 1964 128872 1970
rect 128820 1906 128872 1912
rect 128450 1456 128506 1465
rect 128924 1426 128952 8366
rect 129096 8288 129148 8294
rect 129096 8230 129148 8236
rect 129108 7886 129136 8230
rect 129292 8090 129320 10231
rect 129660 9722 129688 10231
rect 130108 10056 130160 10062
rect 130108 9998 130160 10004
rect 129648 9716 129700 9722
rect 129648 9658 129700 9664
rect 129372 9580 129424 9586
rect 129372 9522 129424 9528
rect 129384 8634 129412 9522
rect 130120 8974 130148 9998
rect 130200 9920 130252 9926
rect 130200 9862 130252 9868
rect 130108 8968 130160 8974
rect 130108 8910 130160 8916
rect 129372 8628 129424 8634
rect 129372 8570 129424 8576
rect 129280 8084 129332 8090
rect 129280 8026 129332 8032
rect 129096 7880 129148 7886
rect 129096 7822 129148 7828
rect 129004 2440 129056 2446
rect 129004 2382 129056 2388
rect 129648 2440 129700 2446
rect 129648 2382 129700 2388
rect 129016 1562 129044 2382
rect 129188 2304 129240 2310
rect 129188 2246 129240 2252
rect 129096 1896 129148 1902
rect 129096 1838 129148 1844
rect 129004 1556 129056 1562
rect 129004 1498 129056 1504
rect 128450 1391 128506 1400
rect 128912 1420 128964 1426
rect 128912 1362 128964 1368
rect 129108 1358 129136 1838
rect 126428 1352 126480 1358
rect 126428 1294 126480 1300
rect 127624 1352 127676 1358
rect 127624 1294 127676 1300
rect 129096 1352 129148 1358
rect 129096 1294 129148 1300
rect 127808 1216 127860 1222
rect 127808 1158 127860 1164
rect 124402 640 124458 649
rect 124402 575 124458 584
rect 125322 640 125378 649
rect 125322 575 125378 584
rect 126242 640 126298 649
rect 126242 575 126298 584
rect 127820 513 127848 1158
rect 129200 649 129228 2246
rect 129660 1902 129688 2382
rect 130120 1970 130148 8910
rect 130212 8430 130240 9862
rect 130764 9722 130792 10231
rect 131486 10231 131542 10240
rect 131120 10202 131172 10208
rect 131500 9722 131528 10231
rect 130752 9716 130804 9722
rect 130752 9658 130804 9664
rect 131488 9716 131540 9722
rect 131488 9658 131540 9664
rect 131120 9648 131172 9654
rect 131120 9590 131172 9596
rect 130568 9580 130620 9586
rect 130568 9522 130620 9528
rect 130580 9178 130608 9522
rect 130568 9172 130620 9178
rect 130568 9114 130620 9120
rect 131132 8974 131160 9590
rect 131396 9580 131448 9586
rect 131396 9522 131448 9528
rect 131408 9178 131436 9522
rect 131396 9172 131448 9178
rect 131396 9114 131448 9120
rect 131868 8974 131896 10610
rect 132130 10296 132186 10305
rect 132130 10231 132186 10240
rect 131120 8968 131172 8974
rect 131120 8910 131172 8916
rect 131856 8968 131908 8974
rect 131856 8910 131908 8916
rect 130844 8900 130896 8906
rect 130844 8842 130896 8848
rect 130856 8430 130884 8842
rect 130200 8424 130252 8430
rect 130200 8366 130252 8372
rect 130844 8424 130896 8430
rect 130844 8366 130896 8372
rect 130212 2514 130240 8366
rect 130384 6452 130436 6458
rect 130384 6394 130436 6400
rect 130396 6254 130424 6394
rect 130384 6248 130436 6254
rect 130384 6190 130436 6196
rect 130200 2508 130252 2514
rect 130200 2450 130252 2456
rect 130752 2304 130804 2310
rect 130752 2246 130804 2252
rect 130108 1964 130160 1970
rect 130108 1906 130160 1912
rect 129648 1896 129700 1902
rect 129648 1838 129700 1844
rect 130660 1760 130712 1766
rect 130660 1702 130712 1708
rect 130672 1358 130700 1702
rect 130660 1352 130712 1358
rect 130660 1294 130712 1300
rect 129186 640 129242 649
rect 129186 575 129242 584
rect 117778 504 117834 513
rect 105728 468 105780 474
rect 105728 410 105780 416
rect 110972 468 111024 474
rect 117778 439 117834 448
rect 118054 504 118110 513
rect 118054 439 118110 448
rect 118698 504 118754 513
rect 118698 439 118754 448
rect 119342 504 119398 513
rect 119342 439 119398 448
rect 120354 504 120410 513
rect 120354 439 120410 448
rect 121090 504 121146 513
rect 121090 439 121146 448
rect 121826 504 121882 513
rect 121826 439 121882 448
rect 122654 504 122710 513
rect 122654 439 122710 448
rect 123390 504 123446 513
rect 123390 439 123446 448
rect 127806 504 127862 513
rect 127806 439 127862 448
rect 110972 410 111024 416
rect 130764 377 130792 2246
rect 131132 1970 131160 8910
rect 131764 2440 131816 2446
rect 131764 2382 131816 2388
rect 131672 2304 131724 2310
rect 131672 2246 131724 2252
rect 131120 1964 131172 1970
rect 131120 1906 131172 1912
rect 130844 1216 130896 1222
rect 130844 1158 130896 1164
rect 130856 649 130884 1158
rect 131684 649 131712 2246
rect 131776 2038 131804 2382
rect 131764 2032 131816 2038
rect 131764 1974 131816 1980
rect 131868 1970 131896 8910
rect 131948 8832 132000 8838
rect 131948 8774 132000 8780
rect 131960 8498 131988 8774
rect 132144 8634 132172 10231
rect 132684 9444 132736 9450
rect 132684 9386 132736 9392
rect 132592 8968 132644 8974
rect 132592 8910 132644 8916
rect 132132 8628 132184 8634
rect 132132 8570 132184 8576
rect 131948 8492 132000 8498
rect 131948 8434 132000 8440
rect 132604 1970 132632 8910
rect 132696 8430 132724 9386
rect 132788 8974 132816 10746
rect 132958 10296 133014 10305
rect 132958 10231 133014 10240
rect 133418 10296 133474 10305
rect 133800 10266 133828 10746
rect 145380 10464 145432 10470
rect 145380 10406 145432 10412
rect 140228 10328 140280 10334
rect 134154 10296 134210 10305
rect 133418 10231 133474 10240
rect 133788 10260 133840 10266
rect 132776 8968 132828 8974
rect 132776 8910 132828 8916
rect 132868 8968 132920 8974
rect 132868 8910 132920 8916
rect 132880 8498 132908 8910
rect 132868 8492 132920 8498
rect 132868 8434 132920 8440
rect 132684 8424 132736 8430
rect 132684 8366 132736 8372
rect 132696 6914 132724 8366
rect 132776 8288 132828 8294
rect 132776 8230 132828 8236
rect 132788 7886 132816 8230
rect 132972 8090 133000 10231
rect 133432 9722 133460 10231
rect 134154 10231 134210 10240
rect 134706 10296 134762 10305
rect 134706 10231 134762 10240
rect 138754 10296 138810 10305
rect 140228 10270 140280 10276
rect 143262 10296 143318 10305
rect 138754 10231 138810 10240
rect 133788 10202 133840 10208
rect 134168 9722 134196 10231
rect 133420 9716 133472 9722
rect 133420 9658 133472 9664
rect 134156 9716 134208 9722
rect 134156 9658 134208 9664
rect 133052 9580 133104 9586
rect 133052 9522 133104 9528
rect 134064 9580 134116 9586
rect 134064 9522 134116 9528
rect 133064 9178 133092 9522
rect 134076 9178 134104 9522
rect 134720 9178 134748 10231
rect 136143 9820 136451 9829
rect 136143 9818 136149 9820
rect 136205 9818 136229 9820
rect 136285 9818 136309 9820
rect 136365 9818 136389 9820
rect 136445 9818 136451 9820
rect 136205 9766 136207 9818
rect 136387 9766 136389 9818
rect 136143 9764 136149 9766
rect 136205 9764 136229 9766
rect 136285 9764 136309 9766
rect 136365 9764 136389 9766
rect 136445 9764 136451 9766
rect 136143 9755 136451 9764
rect 138018 9616 138074 9625
rect 138768 9586 138796 10231
rect 139398 10160 139454 10169
rect 139398 10095 139454 10104
rect 139412 9586 139440 10095
rect 139766 9888 139822 9897
rect 139766 9823 139822 9832
rect 138018 9551 138020 9560
rect 138072 9551 138074 9560
rect 138756 9580 138808 9586
rect 138020 9522 138072 9528
rect 138756 9522 138808 9528
rect 139400 9580 139452 9586
rect 139400 9522 139452 9528
rect 138572 9376 138624 9382
rect 138572 9318 138624 9324
rect 133052 9172 133104 9178
rect 133052 9114 133104 9120
rect 134064 9172 134116 9178
rect 134064 9114 134116 9120
rect 134708 9172 134760 9178
rect 134708 9114 134760 9120
rect 133880 9104 133932 9110
rect 133880 9046 133932 9052
rect 133788 8968 133840 8974
rect 133892 8922 133920 9046
rect 133840 8916 133920 8922
rect 133788 8910 133920 8916
rect 134524 8968 134576 8974
rect 134524 8910 134576 8916
rect 133800 8894 133920 8910
rect 133892 8838 133920 8894
rect 133880 8832 133932 8838
rect 133880 8774 133932 8780
rect 134156 8832 134208 8838
rect 134156 8774 134208 8780
rect 132960 8084 133012 8090
rect 132960 8026 133012 8032
rect 132776 7880 132828 7886
rect 132776 7822 132828 7828
rect 132696 6886 132816 6914
rect 131856 1964 131908 1970
rect 131856 1906 131908 1912
rect 132592 1964 132644 1970
rect 132592 1906 132644 1912
rect 132684 1760 132736 1766
rect 132684 1702 132736 1708
rect 132696 1358 132724 1702
rect 132788 1426 132816 6886
rect 133236 6860 133288 6866
rect 133236 6802 133288 6808
rect 132868 6384 132920 6390
rect 132868 6326 132920 6332
rect 132880 5642 132908 6326
rect 133248 5642 133276 6802
rect 132868 5636 132920 5642
rect 132868 5578 132920 5584
rect 133236 5636 133288 5642
rect 133236 5578 133288 5584
rect 133786 2816 133842 2825
rect 133842 2774 133920 2802
rect 133786 2751 133842 2760
rect 133892 2650 133920 2774
rect 133880 2644 133932 2650
rect 133880 2586 133932 2592
rect 134168 2553 134196 8774
rect 134536 8634 134564 8910
rect 136143 8732 136451 8741
rect 136143 8730 136149 8732
rect 136205 8730 136229 8732
rect 136285 8730 136309 8732
rect 136365 8730 136389 8732
rect 136445 8730 136451 8732
rect 136205 8678 136207 8730
rect 136387 8678 136389 8730
rect 136143 8676 136149 8678
rect 136205 8676 136229 8678
rect 136285 8676 136309 8678
rect 136365 8676 136389 8678
rect 136445 8676 136451 8678
rect 136143 8667 136451 8676
rect 134524 8628 134576 8634
rect 134524 8570 134576 8576
rect 137192 8628 137244 8634
rect 137192 8570 137244 8576
rect 135536 8560 135588 8566
rect 135536 8502 135588 8508
rect 134248 8492 134300 8498
rect 134248 8434 134300 8440
rect 134260 7954 134288 8434
rect 134248 7948 134300 7954
rect 134248 7890 134300 7896
rect 135548 6254 135576 8502
rect 136143 7644 136451 7653
rect 136143 7642 136149 7644
rect 136205 7642 136229 7644
rect 136285 7642 136309 7644
rect 136365 7642 136389 7644
rect 136445 7642 136451 7644
rect 136205 7590 136207 7642
rect 136387 7590 136389 7642
rect 136143 7588 136149 7590
rect 136205 7588 136229 7590
rect 136285 7588 136309 7590
rect 136365 7588 136389 7590
rect 136445 7588 136451 7590
rect 136143 7579 136451 7588
rect 136143 6556 136451 6565
rect 136143 6554 136149 6556
rect 136205 6554 136229 6556
rect 136285 6554 136309 6556
rect 136365 6554 136389 6556
rect 136445 6554 136451 6556
rect 136205 6502 136207 6554
rect 136387 6502 136389 6554
rect 136143 6500 136149 6502
rect 136205 6500 136229 6502
rect 136285 6500 136309 6502
rect 136365 6500 136389 6502
rect 136445 6500 136451 6502
rect 136143 6491 136451 6500
rect 137008 6316 137060 6322
rect 137008 6258 137060 6264
rect 135536 6248 135588 6254
rect 135536 6190 135588 6196
rect 135548 5846 135576 6190
rect 137020 6118 137048 6258
rect 137204 6254 137232 8570
rect 137192 6248 137244 6254
rect 137192 6190 137244 6196
rect 137008 6112 137060 6118
rect 137008 6054 137060 6060
rect 135536 5840 135588 5846
rect 135536 5782 135588 5788
rect 137204 5778 137232 6190
rect 137282 5808 137338 5817
rect 137192 5772 137244 5778
rect 137282 5743 137338 5752
rect 137192 5714 137244 5720
rect 136088 5704 136140 5710
rect 136086 5672 136088 5681
rect 136140 5672 136142 5681
rect 136086 5607 136142 5616
rect 135904 5568 135956 5574
rect 135904 5510 135956 5516
rect 135916 5030 135944 5510
rect 136143 5468 136451 5477
rect 136143 5466 136149 5468
rect 136205 5466 136229 5468
rect 136285 5466 136309 5468
rect 136365 5466 136389 5468
rect 136445 5466 136451 5468
rect 136205 5414 136207 5466
rect 136387 5414 136389 5466
rect 136143 5412 136149 5414
rect 136205 5412 136229 5414
rect 136285 5412 136309 5414
rect 136365 5412 136389 5414
rect 136445 5412 136451 5414
rect 136143 5403 136451 5412
rect 137296 5098 137324 5743
rect 138112 5704 138164 5710
rect 138112 5646 138164 5652
rect 137468 5228 137520 5234
rect 137468 5170 137520 5176
rect 137284 5092 137336 5098
rect 137284 5034 137336 5040
rect 135904 5024 135956 5030
rect 135904 4966 135956 4972
rect 135916 4486 135944 4966
rect 137480 4826 137508 5170
rect 138124 5098 138152 5646
rect 138112 5092 138164 5098
rect 138112 5034 138164 5040
rect 137468 4820 137520 4826
rect 137468 4762 137520 4768
rect 138584 4690 138612 9318
rect 139780 8974 139808 9823
rect 139768 8968 139820 8974
rect 139768 8910 139820 8916
rect 139308 8832 139360 8838
rect 139308 8774 139360 8780
rect 138846 7576 138902 7585
rect 138846 7511 138902 7520
rect 138664 6316 138716 6322
rect 138664 6258 138716 6264
rect 138676 4706 138704 6258
rect 138756 5772 138808 5778
rect 138756 5714 138808 5720
rect 138768 5234 138796 5714
rect 138756 5228 138808 5234
rect 138756 5170 138808 5176
rect 138860 4826 138888 7511
rect 139216 7336 139268 7342
rect 139216 7278 139268 7284
rect 139032 5092 139084 5098
rect 139032 5034 139084 5040
rect 138848 4820 138900 4826
rect 138848 4762 138900 4768
rect 138676 4690 138888 4706
rect 138572 4684 138624 4690
rect 138676 4684 138900 4690
rect 138676 4678 138848 4684
rect 138572 4626 138624 4632
rect 138848 4626 138900 4632
rect 138388 4616 138440 4622
rect 138388 4558 138440 4564
rect 135904 4480 135956 4486
rect 135904 4422 135956 4428
rect 136143 4380 136451 4389
rect 136143 4378 136149 4380
rect 136205 4378 136229 4380
rect 136285 4378 136309 4380
rect 136365 4378 136389 4380
rect 136445 4378 136451 4380
rect 136205 4326 136207 4378
rect 136387 4326 136389 4378
rect 136143 4324 136149 4326
rect 136205 4324 136229 4326
rect 136285 4324 136309 4326
rect 136365 4324 136389 4326
rect 136445 4324 136451 4326
rect 136143 4315 136451 4324
rect 138296 3392 138348 3398
rect 138296 3334 138348 3340
rect 136143 3292 136451 3301
rect 136143 3290 136149 3292
rect 136205 3290 136229 3292
rect 136285 3290 136309 3292
rect 136365 3290 136389 3292
rect 136445 3290 136451 3292
rect 136205 3238 136207 3290
rect 136387 3238 136389 3290
rect 136143 3236 136149 3238
rect 136205 3236 136229 3238
rect 136285 3236 136309 3238
rect 136365 3236 136389 3238
rect 136445 3236 136451 3238
rect 136143 3227 136451 3236
rect 138308 3126 138336 3334
rect 138296 3120 138348 3126
rect 138296 3062 138348 3068
rect 135352 2984 135404 2990
rect 135352 2926 135404 2932
rect 134154 2544 134210 2553
rect 135364 2514 135392 2926
rect 138204 2848 138256 2854
rect 138204 2790 138256 2796
rect 138216 2530 138244 2790
rect 134154 2479 134210 2488
rect 135352 2508 135404 2514
rect 133512 2440 133564 2446
rect 133512 2382 133564 2388
rect 133696 2440 133748 2446
rect 133696 2382 133748 2388
rect 133236 2304 133288 2310
rect 133236 2246 133288 2252
rect 132776 1420 132828 1426
rect 132776 1362 132828 1368
rect 132684 1352 132736 1358
rect 132684 1294 132736 1300
rect 132132 1216 132184 1222
rect 132132 1158 132184 1164
rect 130842 640 130898 649
rect 130842 575 130898 584
rect 131670 640 131726 649
rect 131670 575 131726 584
rect 132144 377 132172 1158
rect 133248 377 133276 2246
rect 133420 1964 133472 1970
rect 133420 1906 133472 1912
rect 133432 1358 133460 1906
rect 133524 1494 133552 2382
rect 133708 2106 133736 2382
rect 133696 2100 133748 2106
rect 133696 2042 133748 2048
rect 134168 1902 134196 2479
rect 138216 2502 138336 2530
rect 135352 2450 135404 2456
rect 134340 2440 134392 2446
rect 134340 2382 134392 2388
rect 134352 1970 134380 2382
rect 135352 2304 135404 2310
rect 135352 2246 135404 2252
rect 135364 1970 135392 2246
rect 136143 2204 136451 2213
rect 136143 2202 136149 2204
rect 136205 2202 136229 2204
rect 136285 2202 136309 2204
rect 136365 2202 136389 2204
rect 136445 2202 136451 2204
rect 136205 2150 136207 2202
rect 136387 2150 136389 2202
rect 136143 2148 136149 2150
rect 136205 2148 136229 2150
rect 136285 2148 136309 2150
rect 136365 2148 136389 2150
rect 136445 2148 136451 2150
rect 136143 2139 136451 2148
rect 134340 1964 134392 1970
rect 134340 1906 134392 1912
rect 135352 1964 135404 1970
rect 135352 1906 135404 1912
rect 134156 1896 134208 1902
rect 134156 1838 134208 1844
rect 134340 1760 134392 1766
rect 134340 1702 134392 1708
rect 135260 1760 135312 1766
rect 135260 1702 135312 1708
rect 133512 1488 133564 1494
rect 133512 1430 133564 1436
rect 134352 1358 134380 1702
rect 135272 1465 135300 1702
rect 138308 1562 138336 2502
rect 138296 1556 138348 1562
rect 138296 1498 138348 1504
rect 138020 1488 138072 1494
rect 135258 1456 135314 1465
rect 135258 1391 135314 1400
rect 138018 1456 138020 1465
rect 138072 1456 138074 1465
rect 138018 1391 138074 1400
rect 133420 1352 133472 1358
rect 133420 1294 133472 1300
rect 134340 1352 134392 1358
rect 134340 1294 134392 1300
rect 138400 1222 138428 4558
rect 138860 4214 138888 4626
rect 138848 4208 138900 4214
rect 138848 4150 138900 4156
rect 139044 4078 139072 5034
rect 139124 4820 139176 4826
rect 139124 4762 139176 4768
rect 139032 4072 139084 4078
rect 139032 4014 139084 4020
rect 138940 3936 138992 3942
rect 138940 3878 138992 3884
rect 138952 3534 138980 3878
rect 139136 3534 139164 4762
rect 139228 4690 139256 7278
rect 139216 4684 139268 4690
rect 139216 4626 139268 4632
rect 139214 4448 139270 4457
rect 139214 4383 139270 4392
rect 138940 3528 138992 3534
rect 138940 3470 138992 3476
rect 139124 3528 139176 3534
rect 139124 3470 139176 3476
rect 139032 3392 139084 3398
rect 139032 3334 139084 3340
rect 139044 3058 139072 3334
rect 138940 3052 138992 3058
rect 138940 2994 138992 3000
rect 139032 3052 139084 3058
rect 139032 2994 139084 3000
rect 138952 2582 138980 2994
rect 138940 2576 138992 2582
rect 138940 2518 138992 2524
rect 138940 2032 138992 2038
rect 138940 1974 138992 1980
rect 138756 1352 138808 1358
rect 138756 1294 138808 1300
rect 138848 1352 138900 1358
rect 138848 1294 138900 1300
rect 134524 1216 134576 1222
rect 134524 1158 134576 1164
rect 138388 1216 138440 1222
rect 138388 1158 138440 1164
rect 134536 649 134564 1158
rect 136143 1116 136451 1125
rect 136143 1114 136149 1116
rect 136205 1114 136229 1116
rect 136285 1114 136309 1116
rect 136365 1114 136389 1116
rect 136445 1114 136451 1116
rect 136205 1062 136207 1114
rect 136387 1062 136389 1114
rect 136143 1060 136149 1062
rect 136205 1060 136229 1062
rect 136285 1060 136309 1062
rect 136365 1060 136389 1062
rect 136445 1060 136451 1062
rect 136143 1051 136451 1060
rect 138768 649 138796 1294
rect 138860 785 138888 1294
rect 138952 950 138980 1974
rect 139032 1964 139084 1970
rect 139032 1906 139084 1912
rect 139044 1834 139072 1906
rect 139032 1828 139084 1834
rect 139032 1770 139084 1776
rect 139228 1222 139256 4383
rect 139320 2514 139348 8774
rect 139766 6352 139822 6361
rect 139766 6287 139822 6296
rect 140044 6316 140096 6322
rect 139584 6248 139636 6254
rect 139584 6190 139636 6196
rect 139400 5228 139452 5234
rect 139400 5170 139452 5176
rect 139412 4146 139440 5170
rect 139596 5166 139624 6190
rect 139780 5953 139808 6287
rect 140044 6258 140096 6264
rect 139952 6112 140004 6118
rect 139952 6054 140004 6060
rect 139766 5944 139822 5953
rect 139766 5879 139822 5888
rect 139780 5710 139808 5879
rect 139768 5704 139820 5710
rect 139768 5646 139820 5652
rect 139584 5160 139636 5166
rect 139584 5102 139636 5108
rect 139768 5160 139820 5166
rect 139768 5102 139820 5108
rect 139492 5024 139544 5030
rect 139492 4966 139544 4972
rect 139400 4140 139452 4146
rect 139400 4082 139452 4088
rect 139504 4010 139532 4966
rect 139676 4480 139728 4486
rect 139676 4422 139728 4428
rect 139688 4026 139716 4422
rect 139780 4078 139808 5102
rect 139860 4752 139912 4758
rect 139860 4694 139912 4700
rect 139872 4457 139900 4694
rect 139964 4690 139992 6054
rect 140056 5778 140084 6258
rect 140044 5772 140096 5778
rect 140044 5714 140096 5720
rect 140044 5092 140096 5098
rect 140044 5034 140096 5040
rect 140056 4826 140084 5034
rect 140044 4820 140096 4826
rect 140044 4762 140096 4768
rect 139952 4684 140004 4690
rect 139952 4626 140004 4632
rect 139858 4448 139914 4457
rect 139858 4383 139914 4392
rect 139492 4004 139544 4010
rect 139492 3946 139544 3952
rect 139596 3998 139716 4026
rect 139768 4072 139820 4078
rect 139768 4014 139820 4020
rect 139504 3670 139532 3946
rect 139492 3664 139544 3670
rect 139492 3606 139544 3612
rect 139596 3534 139624 3998
rect 139676 3936 139728 3942
rect 139676 3878 139728 3884
rect 139584 3528 139636 3534
rect 139584 3470 139636 3476
rect 139492 3460 139544 3466
rect 139492 3402 139544 3408
rect 139504 2922 139532 3402
rect 139688 3058 139716 3878
rect 139950 3496 140006 3505
rect 139950 3431 140006 3440
rect 139676 3052 139728 3058
rect 139676 2994 139728 3000
rect 139964 2990 139992 3431
rect 139952 2984 140004 2990
rect 139952 2926 140004 2932
rect 139492 2916 139544 2922
rect 139492 2858 139544 2864
rect 140042 2816 140098 2825
rect 140042 2751 140098 2760
rect 140056 2666 140084 2751
rect 139964 2650 140084 2666
rect 139952 2644 140084 2650
rect 140004 2638 140084 2644
rect 139952 2586 140004 2592
rect 139308 2508 139360 2514
rect 139308 2450 139360 2456
rect 139952 2508 140004 2514
rect 139952 2450 140004 2456
rect 139492 2440 139544 2446
rect 139492 2382 139544 2388
rect 139504 2106 139532 2382
rect 139964 2106 139992 2450
rect 140240 2446 140268 10270
rect 143262 10231 143318 10240
rect 141424 10192 141476 10198
rect 140686 10160 140742 10169
rect 140686 10095 140742 10104
rect 141330 10160 141386 10169
rect 141424 10134 141476 10140
rect 141974 10160 142030 10169
rect 141330 10095 141386 10104
rect 140700 9586 140728 10095
rect 141344 9586 141372 10095
rect 140688 9580 140740 9586
rect 140688 9522 140740 9528
rect 141332 9580 141384 9586
rect 141332 9522 141384 9528
rect 140412 9376 140464 9382
rect 140412 9318 140464 9324
rect 140504 9376 140556 9382
rect 140504 9318 140556 9324
rect 140596 9376 140648 9382
rect 140596 9318 140648 9324
rect 140320 6656 140372 6662
rect 140320 6598 140372 6604
rect 140332 5574 140360 6598
rect 140320 5568 140372 5574
rect 140320 5510 140372 5516
rect 140332 5234 140360 5510
rect 140320 5228 140372 5234
rect 140320 5170 140372 5176
rect 140424 4690 140452 9318
rect 140412 4684 140464 4690
rect 140412 4626 140464 4632
rect 140228 2440 140280 2446
rect 140228 2382 140280 2388
rect 140320 2440 140372 2446
rect 140320 2382 140372 2388
rect 139492 2100 139544 2106
rect 139492 2042 139544 2048
rect 139952 2100 140004 2106
rect 139952 2042 140004 2048
rect 140228 2032 140280 2038
rect 140228 1974 140280 1980
rect 139768 1964 139820 1970
rect 139768 1906 139820 1912
rect 139216 1216 139268 1222
rect 139216 1158 139268 1164
rect 139780 1057 139808 1906
rect 140240 1873 140268 1974
rect 140226 1864 140282 1873
rect 140226 1799 140282 1808
rect 140228 1760 140280 1766
rect 140228 1702 140280 1708
rect 140240 1426 140268 1702
rect 140228 1420 140280 1426
rect 140228 1362 140280 1368
rect 139766 1048 139822 1057
rect 139766 983 139822 992
rect 138940 944 138992 950
rect 138940 886 138992 892
rect 138846 776 138902 785
rect 138846 711 138902 720
rect 134522 640 134578 649
rect 134522 575 134578 584
rect 138754 640 138810 649
rect 138754 575 138810 584
rect 130750 368 130806 377
rect 130750 303 130806 312
rect 132130 368 132186 377
rect 132130 303 132186 312
rect 133234 368 133290 377
rect 133234 303 133290 312
rect 140332 241 140360 2382
rect 140516 1970 140544 9318
rect 140504 1964 140556 1970
rect 140504 1906 140556 1912
rect 140412 1352 140464 1358
rect 140608 1340 140636 9318
rect 141436 9194 141464 10134
rect 141974 10095 142030 10104
rect 142436 10124 142488 10130
rect 141988 9586 142016 10095
rect 142436 10066 142488 10072
rect 141976 9580 142028 9586
rect 141976 9522 142028 9528
rect 141344 9166 141464 9194
rect 140688 5840 140740 5846
rect 140688 5782 140740 5788
rect 140700 5681 140728 5782
rect 140686 5672 140742 5681
rect 140686 5607 140742 5616
rect 141148 4752 141200 4758
rect 141148 4694 141200 4700
rect 141160 4214 141188 4694
rect 141148 4208 141200 4214
rect 141068 4156 141148 4162
rect 141068 4150 141200 4156
rect 141068 4134 141188 4150
rect 140688 4072 140740 4078
rect 140964 4072 141016 4078
rect 140688 4014 140740 4020
rect 140962 4040 140964 4049
rect 141016 4040 141018 4049
rect 140700 3738 140728 4014
rect 140962 3975 141018 3984
rect 140780 3936 140832 3942
rect 140780 3878 140832 3884
rect 140688 3732 140740 3738
rect 140688 3674 140740 3680
rect 140688 2508 140740 2514
rect 140688 2450 140740 2456
rect 140700 2122 140728 2450
rect 140792 2310 140820 3878
rect 140872 3120 140924 3126
rect 140872 3062 140924 3068
rect 140884 2825 140912 3062
rect 140870 2816 140926 2825
rect 140870 2751 140926 2760
rect 140964 2644 141016 2650
rect 140964 2586 141016 2592
rect 140976 2310 141004 2586
rect 140780 2304 140832 2310
rect 140780 2246 140832 2252
rect 140964 2304 141016 2310
rect 140964 2246 141016 2252
rect 140700 2106 140912 2122
rect 140700 2100 140924 2106
rect 140700 2094 140872 2100
rect 140872 2042 140924 2048
rect 141068 1902 141096 4134
rect 141148 2984 141200 2990
rect 141148 2926 141200 2932
rect 141160 2650 141188 2926
rect 141344 2774 141372 9166
rect 141424 9104 141476 9110
rect 141424 9046 141476 9052
rect 141436 4690 141464 9046
rect 142448 6769 142476 10066
rect 143276 9586 143304 10231
rect 143538 10160 143594 10169
rect 143538 10095 143594 10104
rect 144550 10160 144606 10169
rect 144550 10095 144606 10104
rect 143552 9586 143580 10095
rect 144564 9586 144592 10095
rect 144918 9888 144974 9897
rect 144918 9823 144974 9832
rect 143264 9580 143316 9586
rect 143264 9522 143316 9528
rect 143540 9580 143592 9586
rect 143540 9522 143592 9528
rect 144552 9580 144604 9586
rect 144552 9522 144604 9528
rect 142804 9444 142856 9450
rect 142804 9386 142856 9392
rect 142712 9376 142764 9382
rect 142712 9318 142764 9324
rect 142434 6760 142490 6769
rect 142434 6695 142490 6704
rect 142252 6112 142304 6118
rect 142252 6054 142304 6060
rect 141884 5228 141936 5234
rect 141884 5170 141936 5176
rect 141514 4992 141570 5001
rect 141514 4927 141570 4936
rect 141424 4684 141476 4690
rect 141424 4626 141476 4632
rect 141528 4185 141556 4927
rect 141700 4684 141752 4690
rect 141700 4626 141752 4632
rect 141608 4616 141660 4622
rect 141608 4558 141660 4564
rect 141620 4457 141648 4558
rect 141712 4486 141740 4626
rect 141700 4480 141752 4486
rect 141606 4448 141662 4457
rect 141700 4422 141752 4428
rect 141606 4383 141662 4392
rect 141514 4176 141570 4185
rect 141514 4111 141570 4120
rect 141528 3534 141556 4111
rect 141516 3528 141568 3534
rect 141516 3470 141568 3476
rect 141608 3528 141660 3534
rect 141608 3470 141660 3476
rect 141344 2746 141464 2774
rect 141148 2644 141200 2650
rect 141148 2586 141200 2592
rect 141240 2372 141292 2378
rect 141240 2314 141292 2320
rect 141056 1896 141108 1902
rect 141056 1838 141108 1844
rect 140688 1760 140740 1766
rect 140688 1702 140740 1708
rect 140872 1760 140924 1766
rect 140872 1702 140924 1708
rect 140700 1465 140728 1702
rect 140884 1494 140912 1702
rect 141068 1494 141096 1838
rect 141252 1562 141280 2314
rect 141436 1970 141464 2746
rect 141620 2446 141648 3470
rect 141608 2440 141660 2446
rect 141608 2382 141660 2388
rect 141712 2106 141740 4422
rect 141896 4146 141924 5170
rect 142264 5030 142292 6054
rect 142448 5710 142476 6695
rect 142724 6066 142752 9318
rect 142816 9178 142844 9386
rect 143080 9376 143132 9382
rect 143080 9318 143132 9324
rect 144368 9376 144420 9382
rect 144368 9318 144420 9324
rect 142804 9172 142856 9178
rect 142804 9114 142856 9120
rect 142804 8900 142856 8906
rect 142804 8842 142856 8848
rect 142816 8430 142844 8842
rect 142804 8424 142856 8430
rect 142804 8366 142856 8372
rect 142804 6724 142856 6730
rect 142804 6666 142856 6672
rect 142816 6186 142844 6666
rect 142804 6180 142856 6186
rect 142804 6122 142856 6128
rect 142724 6038 142844 6066
rect 142436 5704 142488 5710
rect 142436 5646 142488 5652
rect 142528 5092 142580 5098
rect 142528 5034 142580 5040
rect 142252 5024 142304 5030
rect 142252 4966 142304 4972
rect 142264 4826 142292 4966
rect 142252 4820 142304 4826
rect 142252 4762 142304 4768
rect 142160 4480 142212 4486
rect 142160 4422 142212 4428
rect 141884 4140 141936 4146
rect 141884 4082 141936 4088
rect 141790 4040 141846 4049
rect 141790 3975 141846 3984
rect 141804 2582 141832 3975
rect 141896 3534 141924 4082
rect 142172 4010 142200 4422
rect 142160 4004 142212 4010
rect 142160 3946 142212 3952
rect 142264 3924 142292 4762
rect 142540 4078 142568 5034
rect 142712 5024 142764 5030
rect 142712 4966 142764 4972
rect 142724 4214 142752 4966
rect 142712 4208 142764 4214
rect 142712 4150 142764 4156
rect 142528 4072 142580 4078
rect 142528 4014 142580 4020
rect 142344 3936 142396 3942
rect 142264 3896 142344 3924
rect 142264 3738 142292 3896
rect 142344 3878 142396 3884
rect 142252 3732 142304 3738
rect 142252 3674 142304 3680
rect 141884 3528 141936 3534
rect 141884 3470 141936 3476
rect 141976 3460 142028 3466
rect 141976 3402 142028 3408
rect 141792 2576 141844 2582
rect 141792 2518 141844 2524
rect 141988 2446 142016 3402
rect 142066 3088 142122 3097
rect 142066 3023 142122 3032
rect 142080 2990 142108 3023
rect 142068 2984 142120 2990
rect 142068 2926 142120 2932
rect 142264 2650 142292 3674
rect 142344 3528 142396 3534
rect 142344 3470 142396 3476
rect 142252 2644 142304 2650
rect 142252 2586 142304 2592
rect 141976 2440 142028 2446
rect 141976 2382 142028 2388
rect 142160 2440 142212 2446
rect 142160 2382 142212 2388
rect 141700 2100 141752 2106
rect 141700 2042 141752 2048
rect 141712 1970 141740 2042
rect 141424 1964 141476 1970
rect 141424 1906 141476 1912
rect 141700 1964 141752 1970
rect 141700 1906 141752 1912
rect 141608 1896 141660 1902
rect 141606 1864 141608 1873
rect 141660 1864 141662 1873
rect 141606 1799 141662 1808
rect 141240 1556 141292 1562
rect 141240 1498 141292 1504
rect 140872 1488 140924 1494
rect 140686 1456 140742 1465
rect 140872 1430 140924 1436
rect 141056 1488 141108 1494
rect 141056 1430 141108 1436
rect 141712 1426 141740 1906
rect 142172 1562 142200 2382
rect 142356 2106 142384 3470
rect 142540 3466 142568 4014
rect 142528 3460 142580 3466
rect 142528 3402 142580 3408
rect 142436 2644 142488 2650
rect 142436 2586 142488 2592
rect 142344 2100 142396 2106
rect 142344 2042 142396 2048
rect 142448 1766 142476 2586
rect 142816 1970 142844 6038
rect 142988 4616 143040 4622
rect 142988 4558 143040 4564
rect 143000 4146 143028 4558
rect 142988 4140 143040 4146
rect 142988 4082 143040 4088
rect 142804 1964 142856 1970
rect 142804 1906 142856 1912
rect 142436 1760 142488 1766
rect 142436 1702 142488 1708
rect 142160 1556 142212 1562
rect 142160 1498 142212 1504
rect 140686 1391 140742 1400
rect 141700 1420 141752 1426
rect 141700 1362 141752 1368
rect 143092 1358 143120 9318
rect 143724 8560 143776 8566
rect 143724 8502 143776 8508
rect 143172 6112 143224 6118
rect 143172 6054 143224 6060
rect 143184 4690 143212 6054
rect 143264 5704 143316 5710
rect 143264 5646 143316 5652
rect 143540 5704 143592 5710
rect 143540 5646 143592 5652
rect 143172 4684 143224 4690
rect 143172 4626 143224 4632
rect 143276 4010 143304 5646
rect 143356 5568 143408 5574
rect 143356 5510 143408 5516
rect 143264 4004 143316 4010
rect 143264 3946 143316 3952
rect 143264 3460 143316 3466
rect 143264 3402 143316 3408
rect 143276 2854 143304 3402
rect 143264 2848 143316 2854
rect 143264 2790 143316 2796
rect 143368 2514 143396 5510
rect 143552 5386 143580 5646
rect 143460 5358 143580 5386
rect 143460 5302 143488 5358
rect 143448 5296 143500 5302
rect 143448 5238 143500 5244
rect 143632 5228 143684 5234
rect 143632 5170 143684 5176
rect 143448 5024 143500 5030
rect 143448 4966 143500 4972
rect 143460 4826 143488 4966
rect 143644 4826 143672 5170
rect 143448 4820 143500 4826
rect 143448 4762 143500 4768
rect 143632 4820 143684 4826
rect 143632 4762 143684 4768
rect 143460 3942 143488 4762
rect 143448 3936 143500 3942
rect 143448 3878 143500 3884
rect 143538 3904 143594 3913
rect 143538 3839 143594 3848
rect 143552 2990 143580 3839
rect 143632 3460 143684 3466
rect 143632 3402 143684 3408
rect 143540 2984 143592 2990
rect 143540 2926 143592 2932
rect 143356 2508 143408 2514
rect 143356 2450 143408 2456
rect 143448 1828 143500 1834
rect 143448 1770 143500 1776
rect 143460 1562 143488 1770
rect 143448 1556 143500 1562
rect 143448 1498 143500 1504
rect 143460 1426 143488 1498
rect 143448 1420 143500 1426
rect 143448 1362 143500 1368
rect 140464 1312 140636 1340
rect 141240 1352 141292 1358
rect 140412 1294 140464 1300
rect 141240 1294 141292 1300
rect 141424 1352 141476 1358
rect 141424 1294 141476 1300
rect 143080 1352 143132 1358
rect 143080 1294 143132 1300
rect 100484 206 100536 212
rect 104162 232 104218 241
rect 104162 167 104218 176
rect 140318 232 140374 241
rect 140318 167 140374 176
rect 141252 105 141280 1294
rect 141436 377 141464 1294
rect 141700 1012 141752 1018
rect 141700 954 141752 960
rect 141792 1012 141844 1018
rect 141792 954 141844 960
rect 141712 814 141740 954
rect 141700 808 141752 814
rect 141804 785 141832 954
rect 143644 921 143672 3402
rect 143736 1970 143764 8502
rect 144000 7948 144052 7954
rect 144000 7890 144052 7896
rect 143906 2952 143962 2961
rect 143906 2887 143962 2896
rect 143920 1970 143948 2887
rect 143724 1964 143776 1970
rect 143724 1906 143776 1912
rect 143908 1964 143960 1970
rect 143908 1906 143960 1912
rect 144012 1358 144040 7890
rect 144380 4690 144408 9318
rect 144932 8974 144960 9823
rect 145196 9444 145248 9450
rect 145196 9386 145248 9392
rect 145012 9036 145064 9042
rect 145012 8978 145064 8984
rect 144920 8968 144972 8974
rect 144920 8910 144972 8916
rect 144736 8832 144788 8838
rect 144736 8774 144788 8780
rect 144368 4684 144420 4690
rect 144368 4626 144420 4632
rect 144748 4078 144776 8774
rect 144920 6996 144972 7002
rect 144920 6938 144972 6944
rect 144932 6497 144960 6938
rect 145024 6934 145052 8978
rect 145102 8528 145158 8537
rect 145102 8463 145158 8472
rect 145012 6928 145064 6934
rect 145012 6870 145064 6876
rect 144918 6488 144974 6497
rect 144918 6423 144974 6432
rect 145116 5778 145144 8463
rect 145104 5772 145156 5778
rect 145104 5714 145156 5720
rect 144828 5704 144880 5710
rect 144826 5672 144828 5681
rect 144880 5672 144882 5681
rect 144826 5607 144882 5616
rect 145012 4684 145064 4690
rect 145012 4626 145064 4632
rect 145104 4684 145156 4690
rect 145104 4626 145156 4632
rect 144736 4072 144788 4078
rect 144736 4014 144788 4020
rect 144736 3664 144788 3670
rect 144736 3606 144788 3612
rect 144748 3233 144776 3606
rect 144828 3460 144880 3466
rect 144828 3402 144880 3408
rect 144840 3369 144868 3402
rect 144826 3360 144882 3369
rect 144826 3295 144882 3304
rect 144734 3224 144790 3233
rect 144734 3159 144790 3168
rect 144552 2984 144604 2990
rect 144552 2926 144604 2932
rect 144276 2304 144328 2310
rect 144276 2246 144328 2252
rect 144184 1896 144236 1902
rect 144288 1884 144316 2246
rect 144236 1856 144316 1884
rect 144184 1838 144236 1844
rect 144288 1426 144316 1856
rect 144276 1420 144328 1426
rect 144276 1362 144328 1368
rect 144000 1352 144052 1358
rect 144000 1294 144052 1300
rect 144092 1352 144144 1358
rect 144564 1329 144592 2926
rect 144644 2916 144696 2922
rect 144644 2858 144696 2864
rect 144656 2106 144684 2858
rect 144736 2372 144788 2378
rect 144736 2314 144788 2320
rect 144644 2100 144696 2106
rect 144644 2042 144696 2048
rect 144092 1294 144144 1300
rect 144550 1320 144606 1329
rect 143630 912 143686 921
rect 143630 847 143686 856
rect 144000 808 144052 814
rect 141700 750 141752 756
rect 141790 776 141846 785
rect 144000 750 144052 756
rect 141790 711 141846 720
rect 144012 513 144040 750
rect 144104 610 144132 1294
rect 144550 1255 144606 1264
rect 144748 921 144776 2314
rect 144828 1760 144880 1766
rect 144828 1702 144880 1708
rect 144840 1222 144868 1702
rect 144920 1352 144972 1358
rect 144920 1294 144972 1300
rect 144828 1216 144880 1222
rect 144828 1158 144880 1164
rect 144734 912 144790 921
rect 144734 847 144790 856
rect 144092 604 144144 610
rect 144092 546 144144 552
rect 143998 504 144054 513
rect 143998 439 144054 448
rect 141422 368 141478 377
rect 141422 303 141478 312
rect 144748 270 144776 847
rect 144932 785 144960 1294
rect 144918 776 144974 785
rect 144918 711 144974 720
rect 144920 672 144972 678
rect 144918 640 144920 649
rect 144972 640 144974 649
rect 144918 575 144974 584
rect 145024 406 145052 4626
rect 145116 4214 145144 4626
rect 145104 4208 145156 4214
rect 145104 4150 145156 4156
rect 145208 1970 145236 9386
rect 145392 4690 145420 10406
rect 145838 10160 145894 10169
rect 145838 10095 145894 10104
rect 146298 10160 146354 10169
rect 146298 10095 146354 10104
rect 145852 9586 145880 10095
rect 146312 9586 146340 10095
rect 145840 9580 145892 9586
rect 145840 9522 145892 9528
rect 146300 9580 146352 9586
rect 146300 9522 146352 9528
rect 145748 9376 145800 9382
rect 145748 9318 145800 9324
rect 145564 5636 145616 5642
rect 145564 5578 145616 5584
rect 145576 5370 145604 5578
rect 145564 5364 145616 5370
rect 145564 5306 145616 5312
rect 145576 5166 145604 5306
rect 145564 5160 145616 5166
rect 145564 5102 145616 5108
rect 145656 5024 145708 5030
rect 145656 4966 145708 4972
rect 145380 4684 145432 4690
rect 145380 4626 145432 4632
rect 145564 4616 145616 4622
rect 145564 4558 145616 4564
rect 145576 4185 145604 4558
rect 145562 4176 145618 4185
rect 145562 4111 145618 4120
rect 145564 3936 145616 3942
rect 145564 3878 145616 3884
rect 145576 3466 145604 3878
rect 145564 3460 145616 3466
rect 145564 3402 145616 3408
rect 145668 3126 145696 4966
rect 145656 3120 145708 3126
rect 145656 3062 145708 3068
rect 145472 2848 145524 2854
rect 145470 2816 145472 2825
rect 145524 2816 145526 2825
rect 145470 2751 145526 2760
rect 145380 2440 145432 2446
rect 145380 2382 145432 2388
rect 145196 1964 145248 1970
rect 145196 1906 145248 1912
rect 145392 1562 145420 2382
rect 145760 2106 145788 9318
rect 146484 7880 146536 7886
rect 146484 7822 146536 7828
rect 146300 7200 146352 7206
rect 146300 7142 146352 7148
rect 146392 7200 146444 7206
rect 146392 7142 146444 7148
rect 146312 6361 146340 7142
rect 146298 6352 146354 6361
rect 146298 6287 146354 6296
rect 146404 5166 146432 7142
rect 146392 5160 146444 5166
rect 146392 5102 146444 5108
rect 146300 4480 146352 4486
rect 146300 4422 146352 4428
rect 145840 4072 145892 4078
rect 145840 4014 145892 4020
rect 146208 4072 146260 4078
rect 146208 4014 146260 4020
rect 145852 3738 145880 4014
rect 145840 3732 145892 3738
rect 145840 3674 145892 3680
rect 145932 3664 145984 3670
rect 145932 3606 145984 3612
rect 145944 3466 145972 3606
rect 145932 3460 145984 3466
rect 145932 3402 145984 3408
rect 146220 3210 146248 4014
rect 146312 3398 146340 4422
rect 146404 3641 146432 5102
rect 146390 3632 146446 3641
rect 146390 3567 146446 3576
rect 146496 3505 146524 7822
rect 146482 3496 146538 3505
rect 146482 3431 146538 3440
rect 146300 3392 146352 3398
rect 146300 3334 146352 3340
rect 146220 3182 146432 3210
rect 146300 2508 146352 2514
rect 146300 2450 146352 2456
rect 146312 2417 146340 2450
rect 146298 2408 146354 2417
rect 146404 2378 146432 3182
rect 146496 2990 146524 3431
rect 146484 2984 146536 2990
rect 146484 2926 146536 2932
rect 146298 2343 146354 2352
rect 146392 2372 146444 2378
rect 146392 2314 146444 2320
rect 145748 2100 145800 2106
rect 145748 2042 145800 2048
rect 146404 1986 146432 2314
rect 146312 1958 146432 1986
rect 146588 1970 146616 10746
rect 151728 10736 151780 10742
rect 151728 10678 151780 10684
rect 148692 10600 148744 10606
rect 148414 10568 148470 10577
rect 148692 10542 148744 10548
rect 148414 10503 148470 10512
rect 147126 10160 147182 10169
rect 147126 10095 147182 10104
rect 147140 9586 147168 10095
rect 147864 9648 147916 9654
rect 147864 9590 147916 9596
rect 147128 9580 147180 9586
rect 147128 9522 147180 9528
rect 147128 5772 147180 5778
rect 147128 5714 147180 5720
rect 146852 4684 146904 4690
rect 146852 4626 146904 4632
rect 146864 4146 146892 4626
rect 147140 4622 147168 5714
rect 147496 5296 147548 5302
rect 147496 5238 147548 5244
rect 147128 4616 147180 4622
rect 147128 4558 147180 4564
rect 147312 4548 147364 4554
rect 147312 4490 147364 4496
rect 146852 4140 146904 4146
rect 146852 4082 146904 4088
rect 146666 3768 146722 3777
rect 146666 3703 146722 3712
rect 146680 2650 146708 3703
rect 146668 2644 146720 2650
rect 146668 2586 146720 2592
rect 146864 2310 146892 4082
rect 147324 3942 147352 4490
rect 147508 4146 147536 5238
rect 147496 4140 147548 4146
rect 147496 4082 147548 4088
rect 147876 4010 147904 9590
rect 148428 9586 148456 10503
rect 148416 9580 148468 9586
rect 148416 9522 148468 9528
rect 148048 9444 148100 9450
rect 148048 9386 148100 9392
rect 147956 5704 148008 5710
rect 147956 5646 148008 5652
rect 147968 4146 147996 5646
rect 147956 4140 148008 4146
rect 147956 4082 148008 4088
rect 147864 4004 147916 4010
rect 147864 3946 147916 3952
rect 147312 3936 147364 3942
rect 147312 3878 147364 3884
rect 147218 3496 147274 3505
rect 147218 3431 147220 3440
rect 147272 3431 147274 3440
rect 147220 3402 147272 3408
rect 147232 3194 147260 3402
rect 147220 3188 147272 3194
rect 147220 3130 147272 3136
rect 147404 2916 147456 2922
rect 147404 2858 147456 2864
rect 146852 2304 146904 2310
rect 146852 2246 146904 2252
rect 146576 1964 146628 1970
rect 146312 1834 146340 1958
rect 146576 1906 146628 1912
rect 146864 1902 146892 2246
rect 147416 2106 147444 2858
rect 147586 2136 147642 2145
rect 147404 2100 147456 2106
rect 147586 2071 147642 2080
rect 147404 2042 147456 2048
rect 146392 1896 146444 1902
rect 146392 1838 146444 1844
rect 146668 1896 146720 1902
rect 146668 1838 146720 1844
rect 146852 1896 146904 1902
rect 146852 1838 146904 1844
rect 146300 1828 146352 1834
rect 146300 1770 146352 1776
rect 145380 1556 145432 1562
rect 145380 1498 145432 1504
rect 146312 1494 146340 1770
rect 146404 1494 146432 1838
rect 146680 1562 146708 1838
rect 146864 1737 146892 1838
rect 146850 1728 146906 1737
rect 146850 1663 146906 1672
rect 146668 1556 146720 1562
rect 146668 1498 146720 1504
rect 146300 1488 146352 1494
rect 146300 1430 146352 1436
rect 146392 1488 146444 1494
rect 146392 1430 146444 1436
rect 146208 1420 146260 1426
rect 146208 1362 146260 1368
rect 145840 1352 145892 1358
rect 145840 1294 145892 1300
rect 145852 1018 145880 1294
rect 145840 1012 145892 1018
rect 145840 954 145892 960
rect 146220 678 146248 1362
rect 146208 672 146260 678
rect 146208 614 146260 620
rect 147600 542 147628 2071
rect 148060 1358 148088 9386
rect 148232 9376 148284 9382
rect 148232 9318 148284 9324
rect 148140 6452 148192 6458
rect 148140 6394 148192 6400
rect 148152 5710 148180 6394
rect 148140 5704 148192 5710
rect 148140 5646 148192 5652
rect 148152 5234 148180 5646
rect 148140 5228 148192 5234
rect 148140 5170 148192 5176
rect 148140 5092 148192 5098
rect 148140 5034 148192 5040
rect 148152 4622 148180 5034
rect 148140 4616 148192 4622
rect 148140 4558 148192 4564
rect 148244 3058 148272 9318
rect 148600 9172 148652 9178
rect 148600 9114 148652 9120
rect 148612 8090 148640 9114
rect 148600 8084 148652 8090
rect 148600 8026 148652 8032
rect 148506 6080 148562 6089
rect 148506 6015 148562 6024
rect 148324 5908 148376 5914
rect 148324 5850 148376 5856
rect 148336 5030 148364 5850
rect 148520 5778 148548 6015
rect 148508 5772 148560 5778
rect 148508 5714 148560 5720
rect 148520 5234 148548 5714
rect 148508 5228 148560 5234
rect 148508 5170 148560 5176
rect 148324 5024 148376 5030
rect 148324 4966 148376 4972
rect 148416 4616 148468 4622
rect 148416 4558 148468 4564
rect 148324 4548 148376 4554
rect 148324 4490 148376 4496
rect 148232 3052 148284 3058
rect 148232 2994 148284 3000
rect 148336 2310 148364 4490
rect 148428 4282 148456 4558
rect 148416 4276 148468 4282
rect 148416 4218 148468 4224
rect 148704 3754 148732 10542
rect 149058 10296 149114 10305
rect 149058 10231 149114 10240
rect 149072 9586 149100 10231
rect 149702 10160 149758 10169
rect 149702 10095 149758 10104
rect 150990 10160 151046 10169
rect 150990 10095 151046 10104
rect 151634 10160 151690 10169
rect 151634 10095 151690 10104
rect 149716 9586 149744 10095
rect 150070 9888 150126 9897
rect 150070 9823 150126 9832
rect 149060 9580 149112 9586
rect 149060 9522 149112 9528
rect 149704 9580 149756 9586
rect 149704 9522 149756 9528
rect 148876 9376 148928 9382
rect 148876 9318 148928 9324
rect 148784 8424 148836 8430
rect 148784 8366 148836 8372
rect 148796 5098 148824 8366
rect 148784 5092 148836 5098
rect 148784 5034 148836 5040
rect 148888 4690 148916 9318
rect 149612 9036 149664 9042
rect 149612 8978 149664 8984
rect 149336 7268 149388 7274
rect 149336 7210 149388 7216
rect 148968 6928 149020 6934
rect 148968 6870 149020 6876
rect 148980 6662 149008 6870
rect 148968 6656 149020 6662
rect 148968 6598 149020 6604
rect 149060 6452 149112 6458
rect 149060 6394 149112 6400
rect 149072 6118 149100 6394
rect 149060 6112 149112 6118
rect 149060 6054 149112 6060
rect 148876 4684 148928 4690
rect 148876 4626 148928 4632
rect 148784 4480 148836 4486
rect 148784 4422 148836 4428
rect 148612 3726 148732 3754
rect 148508 3664 148560 3670
rect 148508 3606 148560 3612
rect 148520 2922 148548 3606
rect 148508 2916 148560 2922
rect 148508 2858 148560 2864
rect 148520 2378 148548 2858
rect 148612 2802 148640 3726
rect 148612 2774 148732 2802
rect 148600 2508 148652 2514
rect 148600 2450 148652 2456
rect 148508 2372 148560 2378
rect 148508 2314 148560 2320
rect 148324 2304 148376 2310
rect 148324 2246 148376 2252
rect 148336 1494 148364 2246
rect 148520 1902 148548 2314
rect 148612 2106 148640 2450
rect 148600 2100 148652 2106
rect 148600 2042 148652 2048
rect 148704 1902 148732 2774
rect 148796 2514 148824 4422
rect 149072 4078 149100 6054
rect 149244 5024 149296 5030
rect 149244 4966 149296 4972
rect 149152 4140 149204 4146
rect 149152 4082 149204 4088
rect 149060 4072 149112 4078
rect 149060 4014 149112 4020
rect 149164 3534 149192 4082
rect 149256 3942 149284 4966
rect 149244 3936 149296 3942
rect 149244 3878 149296 3884
rect 149256 3738 149284 3878
rect 149244 3732 149296 3738
rect 149244 3674 149296 3680
rect 149152 3528 149204 3534
rect 149152 3470 149204 3476
rect 149244 3460 149296 3466
rect 149244 3402 149296 3408
rect 149152 2984 149204 2990
rect 149072 2932 149152 2938
rect 149072 2926 149204 2932
rect 149072 2910 149192 2926
rect 149072 2582 149100 2910
rect 149256 2774 149284 3402
rect 149348 3058 149376 7210
rect 149428 4072 149480 4078
rect 149428 4014 149480 4020
rect 149440 3534 149468 4014
rect 149520 3596 149572 3602
rect 149520 3538 149572 3544
rect 149428 3528 149480 3534
rect 149428 3470 149480 3476
rect 149336 3052 149388 3058
rect 149336 2994 149388 3000
rect 149164 2746 149284 2774
rect 149060 2576 149112 2582
rect 149060 2518 149112 2524
rect 148784 2508 148836 2514
rect 148784 2450 148836 2456
rect 148508 1896 148560 1902
rect 148508 1838 148560 1844
rect 148692 1896 148744 1902
rect 148692 1838 148744 1844
rect 148968 1896 149020 1902
rect 148968 1838 149020 1844
rect 148324 1488 148376 1494
rect 148324 1430 148376 1436
rect 148048 1352 148100 1358
rect 148048 1294 148100 1300
rect 148322 1048 148378 1057
rect 147680 1012 147732 1018
rect 148322 983 148378 992
rect 147680 954 147732 960
rect 147692 785 147720 954
rect 148336 882 148364 983
rect 148324 876 148376 882
rect 148324 818 148376 824
rect 148416 876 148468 882
rect 148416 818 148468 824
rect 148428 785 148456 818
rect 147678 776 147734 785
rect 148414 776 148470 785
rect 147678 711 147734 720
rect 147864 740 147916 746
rect 148414 711 148470 720
rect 147864 682 147916 688
rect 147680 672 147732 678
rect 147876 649 147904 682
rect 147680 614 147732 620
rect 147862 640 147918 649
rect 147588 536 147640 542
rect 147588 478 147640 484
rect 146944 468 146996 474
rect 146944 410 146996 416
rect 145012 400 145064 406
rect 146956 377 146984 410
rect 145012 342 145064 348
rect 146942 368 146998 377
rect 147692 338 147720 614
rect 147862 575 147918 584
rect 148980 474 149008 1838
rect 149164 1358 149192 2746
rect 149336 1896 149388 1902
rect 149336 1838 149388 1844
rect 149348 1737 149376 1838
rect 149334 1728 149390 1737
rect 149334 1663 149390 1672
rect 149152 1352 149204 1358
rect 149152 1294 149204 1300
rect 149336 1352 149388 1358
rect 149336 1294 149388 1300
rect 148968 468 149020 474
rect 148968 410 149020 416
rect 146942 303 146998 312
rect 147680 332 147732 338
rect 147680 274 147732 280
rect 144736 264 144788 270
rect 144736 206 144788 212
rect 29000 70 29052 76
rect 92202 96 92258 105
rect 92202 31 92258 40
rect 98274 96 98330 105
rect 98274 31 98330 40
rect 141238 96 141294 105
rect 149348 66 149376 1294
rect 149532 1193 149560 3538
rect 149624 3466 149652 8978
rect 150084 8974 150112 9823
rect 151004 9586 151032 10095
rect 151648 9586 151676 10095
rect 150992 9580 151044 9586
rect 150992 9522 151044 9528
rect 151636 9580 151688 9586
rect 151636 9522 151688 9528
rect 150716 9444 150768 9450
rect 150716 9386 150768 9392
rect 150532 9376 150584 9382
rect 150532 9318 150584 9324
rect 150072 8968 150124 8974
rect 150072 8910 150124 8916
rect 150348 8832 150400 8838
rect 150348 8774 150400 8780
rect 149978 7984 150034 7993
rect 149978 7919 150034 7928
rect 149796 5908 149848 5914
rect 149796 5850 149848 5856
rect 149808 5642 149836 5850
rect 149704 5636 149756 5642
rect 149704 5578 149756 5584
rect 149796 5636 149848 5642
rect 149796 5578 149848 5584
rect 149716 5234 149744 5578
rect 149704 5228 149756 5234
rect 149704 5170 149756 5176
rect 149808 5030 149836 5578
rect 149992 5273 150020 7919
rect 150256 6452 150308 6458
rect 150256 6394 150308 6400
rect 150164 6248 150216 6254
rect 150164 6190 150216 6196
rect 150072 6112 150124 6118
rect 150072 6054 150124 6060
rect 150084 5545 150112 6054
rect 150070 5536 150126 5545
rect 150070 5471 150126 5480
rect 149978 5264 150034 5273
rect 149978 5199 150034 5208
rect 149796 5024 149848 5030
rect 149796 4966 149848 4972
rect 149992 4865 150020 5199
rect 150176 4865 150204 6190
rect 150268 5710 150296 6394
rect 150360 5710 150388 8774
rect 150440 6928 150492 6934
rect 150440 6870 150492 6876
rect 150256 5704 150308 5710
rect 150256 5646 150308 5652
rect 150348 5704 150400 5710
rect 150348 5646 150400 5652
rect 150254 5264 150310 5273
rect 150254 5199 150310 5208
rect 149978 4856 150034 4865
rect 149978 4791 150034 4800
rect 150162 4856 150218 4865
rect 150162 4791 150218 4800
rect 149886 4720 149942 4729
rect 149886 4655 149888 4664
rect 149940 4655 149942 4664
rect 150164 4684 150216 4690
rect 149888 4626 149940 4632
rect 150164 4626 150216 4632
rect 150072 4616 150124 4622
rect 150072 4558 150124 4564
rect 150084 4321 150112 4558
rect 150070 4312 150126 4321
rect 150070 4247 150126 4256
rect 149980 4004 150032 4010
rect 149980 3946 150032 3952
rect 149612 3460 149664 3466
rect 149612 3402 149664 3408
rect 149610 3224 149666 3233
rect 149610 3159 149666 3168
rect 149624 3058 149652 3159
rect 149612 3052 149664 3058
rect 149664 3012 149744 3040
rect 149612 2994 149664 3000
rect 149610 2000 149666 2009
rect 149610 1935 149666 1944
rect 149624 1737 149652 1935
rect 149716 1902 149744 3012
rect 149992 2009 150020 3946
rect 149978 2000 150034 2009
rect 149978 1935 150034 1944
rect 149704 1896 149756 1902
rect 149704 1838 149756 1844
rect 149610 1728 149666 1737
rect 149610 1663 149666 1672
rect 150176 1426 150204 4626
rect 150268 2514 150296 5199
rect 150452 5098 150480 6870
rect 150544 5234 150572 9318
rect 150624 6792 150676 6798
rect 150624 6734 150676 6740
rect 150636 6322 150664 6734
rect 150624 6316 150676 6322
rect 150624 6258 150676 6264
rect 150636 5302 150664 6258
rect 150624 5296 150676 5302
rect 150624 5238 150676 5244
rect 150532 5228 150584 5234
rect 150532 5170 150584 5176
rect 150636 5098 150664 5238
rect 150440 5092 150492 5098
rect 150440 5034 150492 5040
rect 150624 5092 150676 5098
rect 150624 5034 150676 5040
rect 150348 5024 150400 5030
rect 150728 4978 150756 9386
rect 150808 9376 150860 9382
rect 150808 9318 150860 9324
rect 150820 9042 150848 9318
rect 150808 9036 150860 9042
rect 150808 8978 150860 8984
rect 151452 8356 151504 8362
rect 151452 8298 151504 8304
rect 151464 7206 151492 8298
rect 151740 8294 151768 10678
rect 158548 10674 158576 10814
rect 162768 10736 162820 10742
rect 162768 10678 162820 10684
rect 165068 10736 165120 10742
rect 165068 10678 165120 10684
rect 158536 10668 158588 10674
rect 158536 10610 158588 10616
rect 158628 10668 158680 10674
rect 158628 10610 158680 10616
rect 154302 10432 154358 10441
rect 154302 10367 154358 10376
rect 152278 10160 152334 10169
rect 152830 10160 152886 10169
rect 152278 10095 152334 10104
rect 152556 10124 152608 10130
rect 152292 9586 152320 10095
rect 152830 10095 152886 10104
rect 154210 10160 154266 10169
rect 154210 10095 154266 10104
rect 152556 10066 152608 10072
rect 152464 9988 152516 9994
rect 152464 9930 152516 9936
rect 152280 9580 152332 9586
rect 152280 9522 152332 9528
rect 152476 9518 152504 9930
rect 152464 9512 152516 9518
rect 152464 9454 152516 9460
rect 152464 9172 152516 9178
rect 152464 9114 152516 9120
rect 152476 8566 152504 9114
rect 152464 8560 152516 8566
rect 152464 8502 152516 8508
rect 151728 8288 151780 8294
rect 151728 8230 151780 8236
rect 152004 7812 152056 7818
rect 152004 7754 152056 7760
rect 151820 7744 151872 7750
rect 151820 7686 151872 7692
rect 151832 7562 151860 7686
rect 151544 7540 151596 7546
rect 151544 7482 151596 7488
rect 151740 7534 151860 7562
rect 151452 7200 151504 7206
rect 151452 7142 151504 7148
rect 151556 7002 151584 7482
rect 151740 7410 151768 7534
rect 151728 7404 151780 7410
rect 151728 7346 151780 7352
rect 151820 7404 151872 7410
rect 151820 7346 151872 7352
rect 151636 7336 151688 7342
rect 151636 7278 151688 7284
rect 150900 6996 150952 7002
rect 150900 6938 150952 6944
rect 151544 6996 151596 7002
rect 151544 6938 151596 6944
rect 150912 6118 150940 6938
rect 151084 6860 151136 6866
rect 151084 6802 151136 6808
rect 150992 6452 151044 6458
rect 150992 6394 151044 6400
rect 151004 6254 151032 6394
rect 150992 6248 151044 6254
rect 150992 6190 151044 6196
rect 150900 6112 150952 6118
rect 150900 6054 150952 6060
rect 150912 5642 150940 6054
rect 150900 5636 150952 5642
rect 150900 5578 150952 5584
rect 150348 4966 150400 4972
rect 150360 4690 150388 4966
rect 150636 4950 150756 4978
rect 150348 4684 150400 4690
rect 150348 4626 150400 4632
rect 150348 4208 150400 4214
rect 150348 4150 150400 4156
rect 150360 3641 150388 4150
rect 150346 3632 150402 3641
rect 150346 3567 150402 3576
rect 150440 3460 150492 3466
rect 150440 3402 150492 3408
rect 150452 3194 150480 3402
rect 150440 3188 150492 3194
rect 150440 3130 150492 3136
rect 150346 2952 150402 2961
rect 150402 2910 150480 2938
rect 150346 2887 150402 2896
rect 150348 2848 150400 2854
rect 150348 2790 150400 2796
rect 150256 2508 150308 2514
rect 150256 2450 150308 2456
rect 150254 1592 150310 1601
rect 150254 1527 150310 1536
rect 150164 1420 150216 1426
rect 150164 1362 150216 1368
rect 149518 1184 149574 1193
rect 149518 1119 149574 1128
rect 150268 950 150296 1527
rect 150360 1426 150388 2790
rect 150452 2378 150480 2910
rect 150440 2372 150492 2378
rect 150440 2314 150492 2320
rect 150636 1970 150664 4950
rect 150912 4826 150940 5578
rect 150992 5160 151044 5166
rect 150992 5102 151044 5108
rect 150900 4820 150952 4826
rect 150900 4762 150952 4768
rect 150808 4480 150860 4486
rect 150808 4422 150860 4428
rect 150820 4146 150848 4422
rect 151004 4282 151032 5102
rect 150992 4276 151044 4282
rect 150992 4218 151044 4224
rect 150808 4140 150860 4146
rect 150808 4082 150860 4088
rect 150808 3664 150860 3670
rect 150808 3606 150860 3612
rect 150820 2514 150848 3606
rect 150808 2508 150860 2514
rect 150808 2450 150860 2456
rect 150900 2440 150952 2446
rect 150900 2382 150952 2388
rect 150624 1964 150676 1970
rect 150624 1906 150676 1912
rect 150624 1828 150676 1834
rect 150624 1770 150676 1776
rect 150636 1465 150664 1770
rect 150622 1456 150678 1465
rect 150348 1420 150400 1426
rect 150622 1391 150678 1400
rect 150348 1362 150400 1368
rect 150912 1358 150940 2382
rect 151096 2310 151124 6802
rect 151544 6792 151596 6798
rect 151544 6734 151596 6740
rect 151452 6656 151504 6662
rect 151452 6598 151504 6604
rect 151464 6458 151492 6598
rect 151268 6452 151320 6458
rect 151268 6394 151320 6400
rect 151452 6452 151504 6458
rect 151452 6394 151504 6400
rect 151280 5778 151308 6394
rect 151556 6254 151584 6734
rect 151544 6248 151596 6254
rect 151544 6190 151596 6196
rect 151268 5772 151320 5778
rect 151268 5714 151320 5720
rect 151360 5772 151412 5778
rect 151360 5714 151412 5720
rect 151176 5704 151228 5710
rect 151176 5646 151228 5652
rect 151372 5658 151400 5714
rect 151084 2304 151136 2310
rect 151084 2246 151136 2252
rect 150900 1352 150952 1358
rect 150900 1294 150952 1300
rect 150992 1352 151044 1358
rect 150992 1294 151044 1300
rect 150808 1216 150860 1222
rect 150808 1158 150860 1164
rect 150256 944 150308 950
rect 150256 886 150308 892
rect 150440 944 150492 950
rect 150440 886 150492 892
rect 150452 785 150480 886
rect 150438 776 150494 785
rect 150438 711 150494 720
rect 150820 406 150848 1158
rect 151004 814 151032 1294
rect 151188 814 151216 5646
rect 151372 5630 151492 5658
rect 151464 5098 151492 5630
rect 151268 5092 151320 5098
rect 151268 5034 151320 5040
rect 151452 5092 151504 5098
rect 151452 5034 151504 5040
rect 151280 4622 151308 5034
rect 151360 4684 151412 4690
rect 151360 4626 151412 4632
rect 151268 4616 151320 4622
rect 151268 4558 151320 4564
rect 151268 2984 151320 2990
rect 151268 2926 151320 2932
rect 151280 2145 151308 2926
rect 151372 2774 151400 4626
rect 151464 3738 151492 5034
rect 151556 4622 151584 6190
rect 151648 5778 151676 7278
rect 151832 6866 151860 7346
rect 151820 6860 151872 6866
rect 151820 6802 151872 6808
rect 151728 6656 151780 6662
rect 152016 6610 152044 7754
rect 152568 7546 152596 10066
rect 152844 9586 152872 10095
rect 154224 9586 154252 10095
rect 154316 9586 154344 10367
rect 158640 9926 158668 10610
rect 158812 10532 158864 10538
rect 158812 10474 158864 10480
rect 160468 10532 160520 10538
rect 160468 10474 160520 10480
rect 158628 9920 158680 9926
rect 155222 9888 155278 9897
rect 158628 9862 158680 9868
rect 158720 9920 158772 9926
rect 158720 9862 158772 9868
rect 155222 9823 155278 9832
rect 152832 9580 152884 9586
rect 152832 9522 152884 9528
rect 154212 9580 154264 9586
rect 154212 9522 154264 9528
rect 154304 9580 154356 9586
rect 154304 9522 154356 9528
rect 153200 9444 153252 9450
rect 153200 9386 153252 9392
rect 152556 7540 152608 7546
rect 152556 7482 152608 7488
rect 152740 7404 152792 7410
rect 152740 7346 152792 7352
rect 152188 7200 152240 7206
rect 152188 7142 152240 7148
rect 152096 6996 152148 7002
rect 152096 6938 152148 6944
rect 152108 6798 152136 6938
rect 152096 6792 152148 6798
rect 152096 6734 152148 6740
rect 151780 6604 151860 6610
rect 151728 6598 151860 6604
rect 151740 6582 151860 6598
rect 151636 5772 151688 5778
rect 151636 5714 151688 5720
rect 151726 5400 151782 5409
rect 151726 5335 151782 5344
rect 151740 5232 151768 5335
rect 151728 5226 151780 5232
rect 151728 5168 151780 5174
rect 151726 5128 151782 5137
rect 151726 5063 151782 5072
rect 151544 4616 151596 4622
rect 151544 4558 151596 4564
rect 151452 3732 151504 3738
rect 151452 3674 151504 3680
rect 151740 3466 151768 5063
rect 151728 3460 151780 3466
rect 151728 3402 151780 3408
rect 151372 2746 151676 2774
rect 151360 2508 151412 2514
rect 151360 2450 151412 2456
rect 151266 2136 151322 2145
rect 151266 2071 151322 2080
rect 151268 1760 151320 1766
rect 151268 1702 151320 1708
rect 151280 1562 151308 1702
rect 151268 1556 151320 1562
rect 151268 1498 151320 1504
rect 151372 1057 151400 2450
rect 151452 2304 151504 2310
rect 151452 2246 151504 2252
rect 151464 1834 151492 2246
rect 151544 1896 151596 1902
rect 151544 1838 151596 1844
rect 151452 1828 151504 1834
rect 151452 1770 151504 1776
rect 151556 1426 151584 1838
rect 151544 1420 151596 1426
rect 151544 1362 151596 1368
rect 151358 1048 151414 1057
rect 151358 983 151414 992
rect 150992 808 151044 814
rect 150992 750 151044 756
rect 151176 808 151228 814
rect 151176 750 151228 756
rect 151648 542 151676 2746
rect 151832 2514 151860 6582
rect 151924 6582 152044 6610
rect 151924 5710 151952 6582
rect 152002 6488 152058 6497
rect 152002 6423 152058 6432
rect 151912 5704 151964 5710
rect 151912 5646 151964 5652
rect 151912 5160 151964 5166
rect 151910 5128 151912 5137
rect 151964 5128 151966 5137
rect 151910 5063 151966 5072
rect 152016 4078 152044 6423
rect 152200 5710 152228 7142
rect 152280 6860 152332 6866
rect 152280 6802 152332 6808
rect 152292 6254 152320 6802
rect 152462 6760 152518 6769
rect 152462 6695 152464 6704
rect 152516 6695 152518 6704
rect 152464 6666 152516 6672
rect 152372 6452 152424 6458
rect 152372 6394 152424 6400
rect 152280 6248 152332 6254
rect 152280 6190 152332 6196
rect 152096 5704 152148 5710
rect 152094 5672 152096 5681
rect 152188 5704 152240 5710
rect 152148 5672 152150 5681
rect 152188 5646 152240 5652
rect 152094 5607 152150 5616
rect 152004 4072 152056 4078
rect 152002 4040 152004 4049
rect 152056 4040 152058 4049
rect 152200 4010 152228 5646
rect 152188 4004 152240 4010
rect 152002 3975 152058 3984
rect 152108 3964 152188 3992
rect 152108 3652 152136 3964
rect 152188 3946 152240 3952
rect 152384 3913 152412 6394
rect 152556 6316 152608 6322
rect 152556 6258 152608 6264
rect 152568 4690 152596 6258
rect 152752 6118 152780 7346
rect 152740 6112 152792 6118
rect 152740 6054 152792 6060
rect 152648 5568 152700 5574
rect 152648 5510 152700 5516
rect 152660 5302 152688 5510
rect 152648 5296 152700 5302
rect 152648 5238 152700 5244
rect 152752 5234 152780 6054
rect 152832 5568 152884 5574
rect 152832 5510 152884 5516
rect 152740 5228 152792 5234
rect 152740 5170 152792 5176
rect 152844 4690 152872 5510
rect 153106 5128 153162 5137
rect 152924 5092 152976 5098
rect 153106 5063 153162 5072
rect 152924 5034 152976 5040
rect 152936 5001 152964 5034
rect 152922 4992 152978 5001
rect 152922 4927 152978 4936
rect 153120 4826 153148 5063
rect 153108 4820 153160 4826
rect 153108 4762 153160 4768
rect 152556 4684 152608 4690
rect 152556 4626 152608 4632
rect 152832 4684 152884 4690
rect 152832 4626 152884 4632
rect 152556 4480 152608 4486
rect 152556 4422 152608 4428
rect 152832 4480 152884 4486
rect 152832 4422 152884 4428
rect 152924 4480 152976 4486
rect 152924 4422 152976 4428
rect 152370 3904 152426 3913
rect 152370 3839 152426 3848
rect 152016 3624 152136 3652
rect 152016 3233 152044 3624
rect 152464 3392 152516 3398
rect 152464 3334 152516 3340
rect 152002 3224 152058 3233
rect 152002 3159 152058 3168
rect 151820 2508 151872 2514
rect 151820 2450 151872 2456
rect 151726 2408 151782 2417
rect 151726 2343 151782 2352
rect 151740 1970 151768 2343
rect 152016 1970 152044 3159
rect 152476 3126 152504 3334
rect 152464 3120 152516 3126
rect 152464 3062 152516 3068
rect 152568 3058 152596 4422
rect 152844 4214 152872 4422
rect 152832 4208 152884 4214
rect 152832 4150 152884 4156
rect 152740 3936 152792 3942
rect 152740 3878 152792 3884
rect 152648 3596 152700 3602
rect 152648 3538 152700 3544
rect 152556 3052 152608 3058
rect 152556 2994 152608 3000
rect 152660 2774 152688 3538
rect 152752 3534 152780 3878
rect 152832 3664 152884 3670
rect 152832 3606 152884 3612
rect 152740 3528 152792 3534
rect 152740 3470 152792 3476
rect 152844 2990 152872 3606
rect 152936 3369 152964 4422
rect 153212 4146 153240 9386
rect 153292 9376 153344 9382
rect 153292 9318 153344 9324
rect 154028 9376 154080 9382
rect 154028 9318 154080 9324
rect 153304 5778 153332 9318
rect 153476 9036 153528 9042
rect 153476 8978 153528 8984
rect 153384 6860 153436 6866
rect 153384 6802 153436 6808
rect 153292 5772 153344 5778
rect 153292 5714 153344 5720
rect 153396 5302 153424 6802
rect 153384 5296 153436 5302
rect 153384 5238 153436 5244
rect 153488 5148 153516 8978
rect 153844 8628 153896 8634
rect 153844 8570 153896 8576
rect 153752 8492 153804 8498
rect 153752 8434 153804 8440
rect 153568 8084 153620 8090
rect 153568 8026 153620 8032
rect 153580 6458 153608 8026
rect 153660 7268 153712 7274
rect 153660 7210 153712 7216
rect 153568 6452 153620 6458
rect 153568 6394 153620 6400
rect 153566 5536 153622 5545
rect 153566 5471 153622 5480
rect 153396 5120 153516 5148
rect 153292 5024 153344 5030
rect 153292 4966 153344 4972
rect 153200 4140 153252 4146
rect 153200 4082 153252 4088
rect 153304 3534 153332 4966
rect 153396 3602 153424 5120
rect 153580 4690 153608 5471
rect 153568 4684 153620 4690
rect 153568 4626 153620 4632
rect 153476 4072 153528 4078
rect 153476 4014 153528 4020
rect 153384 3596 153436 3602
rect 153384 3538 153436 3544
rect 153292 3528 153344 3534
rect 153292 3470 153344 3476
rect 153292 3392 153344 3398
rect 152922 3360 152978 3369
rect 153292 3334 153344 3340
rect 152922 3295 152978 3304
rect 152832 2984 152884 2990
rect 152832 2926 152884 2932
rect 152924 2848 152976 2854
rect 152924 2790 152976 2796
rect 153016 2848 153068 2854
rect 153016 2790 153068 2796
rect 152568 2746 152688 2774
rect 152568 2106 152596 2746
rect 152936 2582 152964 2790
rect 153028 2650 153056 2790
rect 153016 2644 153068 2650
rect 153016 2586 153068 2592
rect 152740 2576 152792 2582
rect 152740 2518 152792 2524
rect 152924 2576 152976 2582
rect 152924 2518 152976 2524
rect 152752 2106 152780 2518
rect 152096 2100 152148 2106
rect 152096 2042 152148 2048
rect 152556 2100 152608 2106
rect 152556 2042 152608 2048
rect 152740 2100 152792 2106
rect 153304 2088 153332 3334
rect 153384 2440 153436 2446
rect 153384 2382 153436 2388
rect 152740 2042 152792 2048
rect 153120 2060 153332 2088
rect 151728 1964 151780 1970
rect 151728 1906 151780 1912
rect 152004 1964 152056 1970
rect 152004 1906 152056 1912
rect 151728 1556 151780 1562
rect 151728 1498 151780 1504
rect 151740 746 151768 1498
rect 152108 1465 152136 2042
rect 153120 1601 153148 2060
rect 153396 1970 153424 2382
rect 153488 2310 153516 4014
rect 153672 3670 153700 7210
rect 153764 6798 153792 8434
rect 153856 6866 153884 8570
rect 154040 8566 154068 9318
rect 155236 8974 155264 9823
rect 158732 9722 158760 9862
rect 158720 9716 158772 9722
rect 158720 9658 158772 9664
rect 155684 9648 155736 9654
rect 155684 9590 155736 9596
rect 155696 9382 155724 9590
rect 157340 9580 157392 9586
rect 157340 9522 157392 9528
rect 157524 9580 157576 9586
rect 157524 9522 157576 9528
rect 156972 9512 157024 9518
rect 156694 9480 156750 9489
rect 156972 9454 157024 9460
rect 156694 9415 156696 9424
rect 156748 9415 156750 9424
rect 156696 9386 156748 9392
rect 155592 9376 155644 9382
rect 155592 9318 155644 9324
rect 155684 9376 155736 9382
rect 155684 9318 155736 9324
rect 155224 8968 155276 8974
rect 155224 8910 155276 8916
rect 155040 8832 155092 8838
rect 155040 8774 155092 8780
rect 154028 8560 154080 8566
rect 154028 8502 154080 8508
rect 154028 8356 154080 8362
rect 154028 8298 154080 8304
rect 154672 8356 154724 8362
rect 154672 8298 154724 8304
rect 153934 7032 153990 7041
rect 153934 6967 153990 6976
rect 153844 6860 153896 6866
rect 153844 6802 153896 6808
rect 153752 6792 153804 6798
rect 153752 6734 153804 6740
rect 153842 6760 153898 6769
rect 153842 6695 153844 6704
rect 153896 6695 153898 6704
rect 153844 6666 153896 6672
rect 153752 6316 153804 6322
rect 153752 6258 153804 6264
rect 153764 6186 153792 6258
rect 153752 6180 153804 6186
rect 153752 6122 153804 6128
rect 153764 5794 153792 6122
rect 153764 5778 153884 5794
rect 153764 5772 153896 5778
rect 153764 5766 153844 5772
rect 153844 5714 153896 5720
rect 153752 4752 153804 4758
rect 153752 4694 153804 4700
rect 153660 3664 153712 3670
rect 153660 3606 153712 3612
rect 153660 2984 153712 2990
rect 153658 2952 153660 2961
rect 153712 2952 153714 2961
rect 153658 2887 153714 2896
rect 153764 2650 153792 4694
rect 153856 4434 153884 5714
rect 153948 5030 153976 6967
rect 154040 5030 154068 8298
rect 154580 7880 154632 7886
rect 154580 7822 154632 7828
rect 154592 7721 154620 7822
rect 154578 7712 154634 7721
rect 154578 7647 154634 7656
rect 154684 7478 154712 8298
rect 154762 8120 154818 8129
rect 154762 8055 154818 8064
rect 154672 7472 154724 7478
rect 154672 7414 154724 7420
rect 154672 7336 154724 7342
rect 154672 7278 154724 7284
rect 154488 5840 154540 5846
rect 154540 5788 154620 5794
rect 154488 5782 154620 5788
rect 154500 5766 154620 5782
rect 154684 5778 154712 7278
rect 153936 5024 153988 5030
rect 153936 4966 153988 4972
rect 154028 5024 154080 5030
rect 154028 4966 154080 4972
rect 154592 4842 154620 5766
rect 154672 5772 154724 5778
rect 154672 5714 154724 5720
rect 154776 5273 154804 8055
rect 155052 6866 155080 8774
rect 155040 6860 155092 6866
rect 155040 6802 155092 6808
rect 154856 6316 154908 6322
rect 154856 6258 154908 6264
rect 154868 5914 154896 6258
rect 154948 6248 155000 6254
rect 154948 6190 155000 6196
rect 154856 5908 154908 5914
rect 154856 5850 154908 5856
rect 154960 5710 154988 6190
rect 154948 5704 155000 5710
rect 154948 5646 155000 5652
rect 154856 5568 154908 5574
rect 154856 5510 154908 5516
rect 154762 5264 154818 5273
rect 154762 5199 154818 5208
rect 154776 5166 154804 5199
rect 154764 5160 154816 5166
rect 154764 5102 154816 5108
rect 154592 4814 154712 4842
rect 154580 4684 154632 4690
rect 154580 4626 154632 4632
rect 154592 4593 154620 4626
rect 154578 4584 154634 4593
rect 154578 4519 154634 4528
rect 153856 4406 153976 4434
rect 153844 4276 153896 4282
rect 153844 4218 153896 4224
rect 153752 2644 153804 2650
rect 153752 2586 153804 2592
rect 153476 2304 153528 2310
rect 153476 2246 153528 2252
rect 153856 2106 153884 4218
rect 153948 4078 153976 4406
rect 154026 4176 154082 4185
rect 154026 4111 154082 4120
rect 153936 4072 153988 4078
rect 153936 4014 153988 4020
rect 153936 3596 153988 3602
rect 153936 3538 153988 3544
rect 153948 2106 153976 3538
rect 153844 2100 153896 2106
rect 153844 2042 153896 2048
rect 153936 2100 153988 2106
rect 153936 2042 153988 2048
rect 153292 1964 153344 1970
rect 153292 1906 153344 1912
rect 153384 1964 153436 1970
rect 153384 1906 153436 1912
rect 153106 1592 153162 1601
rect 153304 1562 153332 1906
rect 153106 1527 153162 1536
rect 153292 1556 153344 1562
rect 153292 1498 153344 1504
rect 152094 1456 152150 1465
rect 152094 1391 152150 1400
rect 152280 1352 152332 1358
rect 153568 1352 153620 1358
rect 152280 1294 152332 1300
rect 152462 1320 152518 1329
rect 152292 1018 152320 1294
rect 152372 1284 152424 1290
rect 153568 1294 153620 1300
rect 152462 1255 152518 1264
rect 152372 1226 152424 1232
rect 152384 1057 152412 1226
rect 152370 1048 152426 1057
rect 152280 1012 152332 1018
rect 152370 983 152426 992
rect 152280 954 152332 960
rect 151728 740 151780 746
rect 151728 682 151780 688
rect 152476 678 152504 1255
rect 152464 672 152516 678
rect 152464 614 152516 620
rect 153580 610 153608 1294
rect 153936 1216 153988 1222
rect 153936 1158 153988 1164
rect 153568 604 153620 610
rect 153568 546 153620 552
rect 153948 542 153976 1158
rect 154040 1018 154068 4111
rect 154120 4072 154172 4078
rect 154120 4014 154172 4020
rect 154212 4072 154264 4078
rect 154212 4014 154264 4020
rect 154132 3233 154160 4014
rect 154118 3224 154174 3233
rect 154118 3159 154174 3168
rect 154120 2440 154172 2446
rect 154120 2382 154172 2388
rect 154028 1012 154080 1018
rect 154028 954 154080 960
rect 154132 649 154160 2382
rect 154224 1714 154252 4014
rect 154580 3936 154632 3942
rect 154580 3878 154632 3884
rect 154304 3732 154356 3738
rect 154304 3674 154356 3680
rect 154316 3369 154344 3674
rect 154592 3534 154620 3878
rect 154488 3528 154540 3534
rect 154488 3470 154540 3476
rect 154580 3528 154632 3534
rect 154580 3470 154632 3476
rect 154302 3360 154358 3369
rect 154302 3295 154358 3304
rect 154394 2816 154450 2825
rect 154394 2751 154450 2760
rect 154408 2281 154436 2751
rect 154500 2582 154528 3470
rect 154684 3058 154712 4814
rect 154764 4820 154816 4826
rect 154764 4762 154816 4768
rect 154672 3052 154724 3058
rect 154672 2994 154724 3000
rect 154488 2576 154540 2582
rect 154488 2518 154540 2524
rect 154488 2440 154540 2446
rect 154488 2382 154540 2388
rect 154394 2272 154450 2281
rect 154394 2207 154450 2216
rect 154224 1686 154344 1714
rect 154212 1352 154264 1358
rect 154212 1294 154264 1300
rect 154224 882 154252 1294
rect 154212 876 154264 882
rect 154212 818 154264 824
rect 154118 640 154174 649
rect 154118 575 154174 584
rect 154316 542 154344 1686
rect 154500 1329 154528 2382
rect 154580 1964 154632 1970
rect 154580 1906 154632 1912
rect 154592 1766 154620 1906
rect 154580 1760 154632 1766
rect 154580 1702 154632 1708
rect 154580 1420 154632 1426
rect 154580 1362 154632 1368
rect 154486 1320 154542 1329
rect 154486 1255 154542 1264
rect 151636 536 151688 542
rect 151636 478 151688 484
rect 153936 536 153988 542
rect 153936 478 153988 484
rect 154304 536 154356 542
rect 154304 478 154356 484
rect 150808 400 150860 406
rect 150808 342 150860 348
rect 154592 338 154620 1362
rect 154672 1216 154724 1222
rect 154672 1158 154724 1164
rect 154684 814 154712 1158
rect 154672 808 154724 814
rect 154672 750 154724 756
rect 154776 338 154804 4762
rect 154868 2774 154896 5510
rect 154960 5166 154988 5646
rect 154948 5160 155000 5166
rect 154948 5102 155000 5108
rect 154960 4214 154988 5102
rect 155316 5024 155368 5030
rect 155316 4966 155368 4972
rect 155132 4480 155184 4486
rect 155132 4422 155184 4428
rect 154948 4208 155000 4214
rect 154948 4150 155000 4156
rect 154948 4004 155000 4010
rect 154948 3946 155000 3952
rect 154960 3602 154988 3946
rect 154948 3596 155000 3602
rect 154948 3538 155000 3544
rect 155040 3120 155092 3126
rect 155040 3062 155092 3068
rect 155052 2961 155080 3062
rect 155038 2952 155094 2961
rect 155038 2887 155094 2896
rect 155144 2854 155172 4422
rect 155224 4072 155276 4078
rect 155224 4014 155276 4020
rect 155236 3738 155264 4014
rect 155224 3732 155276 3738
rect 155224 3674 155276 3680
rect 155224 3596 155276 3602
rect 155224 3538 155276 3544
rect 155132 2848 155184 2854
rect 155132 2790 155184 2796
rect 154868 2746 154988 2774
rect 154960 2106 154988 2746
rect 155236 2650 155264 3538
rect 155224 2644 155276 2650
rect 155224 2586 155276 2592
rect 154948 2100 155000 2106
rect 154948 2042 155000 2048
rect 154856 1352 154908 1358
rect 154856 1294 154908 1300
rect 154868 950 154896 1294
rect 154948 1284 155000 1290
rect 154948 1226 155000 1232
rect 154960 950 154988 1226
rect 154856 944 154908 950
rect 154856 886 154908 892
rect 154948 944 155000 950
rect 154948 886 155000 892
rect 154580 332 154632 338
rect 154580 274 154632 280
rect 154764 332 154816 338
rect 154764 274 154816 280
rect 155328 270 155356 4966
rect 155604 3534 155632 9318
rect 156050 9072 156106 9081
rect 156050 9007 156052 9016
rect 156104 9007 156106 9016
rect 156696 9036 156748 9042
rect 156052 8978 156104 8984
rect 156696 8978 156748 8984
rect 156236 8900 156288 8906
rect 156236 8842 156288 8848
rect 155960 8832 156012 8838
rect 155960 8774 156012 8780
rect 155972 8498 156000 8774
rect 156050 8664 156106 8673
rect 156248 8634 156276 8842
rect 156050 8599 156052 8608
rect 156104 8599 156106 8608
rect 156236 8628 156288 8634
rect 156052 8570 156104 8576
rect 156236 8570 156288 8576
rect 156512 8560 156564 8566
rect 156512 8502 156564 8508
rect 155960 8492 156012 8498
rect 155960 8434 156012 8440
rect 156144 8424 156196 8430
rect 156144 8366 156196 8372
rect 156236 8424 156288 8430
rect 156236 8366 156288 8372
rect 156050 7848 156106 7857
rect 156050 7783 156106 7792
rect 155868 6248 155920 6254
rect 155868 6190 155920 6196
rect 155776 6112 155828 6118
rect 155776 6054 155828 6060
rect 155684 4616 155736 4622
rect 155684 4558 155736 4564
rect 155696 4282 155724 4558
rect 155684 4276 155736 4282
rect 155684 4218 155736 4224
rect 155592 3528 155644 3534
rect 155592 3470 155644 3476
rect 155788 2990 155816 6054
rect 155880 5778 155908 6190
rect 155868 5772 155920 5778
rect 155868 5714 155920 5720
rect 155960 5636 156012 5642
rect 155960 5578 156012 5584
rect 155972 5234 156000 5578
rect 155960 5228 156012 5234
rect 155960 5170 156012 5176
rect 155868 4820 155920 4826
rect 155868 4762 155920 4768
rect 155880 4554 155908 4762
rect 156064 4690 156092 7783
rect 156156 6322 156184 8366
rect 156144 6316 156196 6322
rect 156144 6258 156196 6264
rect 156248 6202 156276 8366
rect 156328 6452 156380 6458
rect 156328 6394 156380 6400
rect 156340 6254 156368 6394
rect 156156 6174 156276 6202
rect 156328 6248 156380 6254
rect 156328 6190 156380 6196
rect 156052 4684 156104 4690
rect 156052 4626 156104 4632
rect 155868 4548 155920 4554
rect 155868 4490 155920 4496
rect 156156 3777 156184 6174
rect 156328 6112 156380 6118
rect 156328 6054 156380 6060
rect 156420 6112 156472 6118
rect 156420 6054 156472 6060
rect 156236 5636 156288 5642
rect 156236 5578 156288 5584
rect 156248 4214 156276 5578
rect 156340 4758 156368 6054
rect 156432 5914 156460 6054
rect 156420 5908 156472 5914
rect 156420 5850 156472 5856
rect 156420 5296 156472 5302
rect 156420 5238 156472 5244
rect 156328 4752 156380 4758
rect 156328 4694 156380 4700
rect 156236 4208 156288 4214
rect 156236 4150 156288 4156
rect 156236 4072 156288 4078
rect 156236 4014 156288 4020
rect 156142 3768 156198 3777
rect 156142 3703 156198 3712
rect 155868 3392 155920 3398
rect 155868 3334 155920 3340
rect 156144 3392 156196 3398
rect 156144 3334 156196 3340
rect 155880 3074 155908 3334
rect 155880 3046 156092 3074
rect 156156 3058 156184 3334
rect 156248 3194 156276 4014
rect 156340 3670 156368 4694
rect 156432 4690 156460 5238
rect 156524 4690 156552 8502
rect 156604 8016 156656 8022
rect 156604 7958 156656 7964
rect 156420 4684 156472 4690
rect 156420 4626 156472 4632
rect 156512 4684 156564 4690
rect 156512 4626 156564 4632
rect 156328 3664 156380 3670
rect 156328 3606 156380 3612
rect 156616 3602 156644 7958
rect 156604 3596 156656 3602
rect 156604 3538 156656 3544
rect 156236 3188 156288 3194
rect 156236 3130 156288 3136
rect 155776 2984 155828 2990
rect 155776 2926 155828 2932
rect 155866 2952 155922 2961
rect 156064 2938 156092 3046
rect 156144 3052 156196 3058
rect 156144 2994 156196 3000
rect 156420 2984 156472 2990
rect 156064 2932 156420 2938
rect 156064 2926 156472 2932
rect 156064 2910 156460 2926
rect 155866 2887 155922 2896
rect 155880 2774 155908 2887
rect 156236 2848 156288 2854
rect 156236 2790 156288 2796
rect 156418 2816 156474 2825
rect 155788 2746 155908 2774
rect 155592 2440 155644 2446
rect 155592 2382 155644 2388
rect 155604 1290 155632 2382
rect 155592 1284 155644 1290
rect 155592 1226 155644 1232
rect 155788 1193 155816 2746
rect 156248 2553 156276 2790
rect 156418 2751 156474 2760
rect 156432 2650 156460 2751
rect 156420 2644 156472 2650
rect 156420 2586 156472 2592
rect 156234 2544 156290 2553
rect 156234 2479 156290 2488
rect 156602 2544 156658 2553
rect 156602 2479 156658 2488
rect 156616 2446 156644 2479
rect 156604 2440 156656 2446
rect 156604 2382 156656 2388
rect 156708 2378 156736 8978
rect 156788 6112 156840 6118
rect 156788 6054 156840 6060
rect 156800 5574 156828 6054
rect 156880 5670 156932 5676
rect 156880 5612 156932 5618
rect 156788 5568 156840 5574
rect 156788 5510 156840 5516
rect 156892 5166 156920 5612
rect 156880 5160 156932 5166
rect 156880 5102 156932 5108
rect 156892 3534 156920 5102
rect 156880 3528 156932 3534
rect 156880 3470 156932 3476
rect 156984 2689 157012 9454
rect 157352 9042 157380 9522
rect 157430 9072 157486 9081
rect 157340 9036 157392 9042
rect 157430 9007 157432 9016
rect 157340 8978 157392 8984
rect 157484 9007 157486 9016
rect 157432 8978 157484 8984
rect 157536 8974 157564 9522
rect 158824 9518 158852 10474
rect 159640 10124 159692 10130
rect 159640 10066 159692 10072
rect 158812 9512 158864 9518
rect 158812 9454 158864 9460
rect 159548 9512 159600 9518
rect 159548 9454 159600 9460
rect 158536 9376 158588 9382
rect 158536 9318 158588 9324
rect 157064 8968 157116 8974
rect 157064 8910 157116 8916
rect 157524 8968 157576 8974
rect 157524 8910 157576 8916
rect 157076 8378 157104 8910
rect 157800 8900 157852 8906
rect 157800 8842 157852 8848
rect 157706 8528 157762 8537
rect 157706 8463 157762 8472
rect 157246 8392 157302 8401
rect 157076 8350 157196 8378
rect 157064 8288 157116 8294
rect 157064 8230 157116 8236
rect 157076 7886 157104 8230
rect 157064 7880 157116 7886
rect 157064 7822 157116 7828
rect 157064 4072 157116 4078
rect 157064 4014 157116 4020
rect 157076 2961 157104 4014
rect 157062 2952 157118 2961
rect 157062 2887 157118 2896
rect 156970 2680 157026 2689
rect 156970 2615 157026 2624
rect 156984 2446 157012 2615
rect 156972 2440 157024 2446
rect 156972 2382 157024 2388
rect 156420 2372 156472 2378
rect 156420 2314 156472 2320
rect 156696 2372 156748 2378
rect 156696 2314 156748 2320
rect 156328 1964 156380 1970
rect 156328 1906 156380 1912
rect 155960 1760 156012 1766
rect 155960 1702 156012 1708
rect 155972 1465 156000 1702
rect 156340 1562 156368 1906
rect 156328 1556 156380 1562
rect 156328 1498 156380 1504
rect 155958 1456 156014 1465
rect 155958 1391 156014 1400
rect 156432 1358 156460 2314
rect 156788 1964 156840 1970
rect 156788 1906 156840 1912
rect 156604 1896 156656 1902
rect 156604 1838 156656 1844
rect 156616 1737 156644 1838
rect 156800 1737 156828 1906
rect 157168 1902 157196 8350
rect 157246 8327 157302 8336
rect 157260 8090 157288 8327
rect 157248 8084 157300 8090
rect 157248 8026 157300 8032
rect 157248 6860 157300 6866
rect 157248 6802 157300 6808
rect 157260 5642 157288 6802
rect 157720 5914 157748 8463
rect 157812 8430 157840 8842
rect 157800 8424 157852 8430
rect 157800 8366 157852 8372
rect 158548 7886 158576 9318
rect 159180 8900 159232 8906
rect 159180 8842 159232 8848
rect 158718 8120 158774 8129
rect 158718 8055 158720 8064
rect 158772 8055 158774 8064
rect 158720 8026 158772 8032
rect 158536 7880 158588 7886
rect 158536 7822 158588 7828
rect 158076 7744 158128 7750
rect 158076 7686 158128 7692
rect 157798 7440 157854 7449
rect 157798 7375 157854 7384
rect 157708 5908 157760 5914
rect 157708 5850 157760 5856
rect 157248 5636 157300 5642
rect 157248 5578 157300 5584
rect 157812 5166 157840 7375
rect 157800 5160 157852 5166
rect 157800 5102 157852 5108
rect 157246 3768 157302 3777
rect 157246 3703 157302 3712
rect 157260 2394 157288 3703
rect 157708 2440 157760 2446
rect 157260 2366 157380 2394
rect 157708 2382 157760 2388
rect 157248 2304 157300 2310
rect 157248 2246 157300 2252
rect 157156 1896 157208 1902
rect 157156 1838 157208 1844
rect 156602 1728 156658 1737
rect 156602 1663 156658 1672
rect 156786 1728 156842 1737
rect 156786 1663 156842 1672
rect 156880 1488 156932 1494
rect 157064 1488 157116 1494
rect 156932 1436 157064 1442
rect 156880 1430 157116 1436
rect 156892 1414 157104 1430
rect 156420 1352 156472 1358
rect 156420 1294 156472 1300
rect 157168 1306 157196 1838
rect 157260 1465 157288 2246
rect 157352 2038 157380 2366
rect 157340 2032 157392 2038
rect 157340 1974 157392 1980
rect 157246 1456 157302 1465
rect 157246 1391 157302 1400
rect 157248 1352 157300 1358
rect 157168 1300 157248 1306
rect 157168 1294 157300 1300
rect 155774 1184 155830 1193
rect 155774 1119 155830 1128
rect 156432 746 156460 1294
rect 157168 1278 157288 1294
rect 157720 1290 157748 2382
rect 157708 1284 157760 1290
rect 157708 1226 157760 1232
rect 156420 740 156472 746
rect 156420 682 156472 688
rect 158088 406 158116 7686
rect 158166 6488 158222 6497
rect 158166 6423 158222 6432
rect 158180 4010 158208 6423
rect 158444 6180 158496 6186
rect 158444 6122 158496 6128
rect 158456 4078 158484 6122
rect 158812 5772 158864 5778
rect 158812 5714 158864 5720
rect 158628 5636 158680 5642
rect 158628 5578 158680 5584
rect 158534 4856 158590 4865
rect 158534 4791 158590 4800
rect 158548 4078 158576 4791
rect 158444 4072 158496 4078
rect 158444 4014 158496 4020
rect 158536 4072 158588 4078
rect 158536 4014 158588 4020
rect 158168 4004 158220 4010
rect 158168 3946 158220 3952
rect 158536 3936 158588 3942
rect 158536 3878 158588 3884
rect 158548 3398 158576 3878
rect 158640 3398 158668 5578
rect 158824 4690 158852 5714
rect 158812 4684 158864 4690
rect 158812 4626 158864 4632
rect 158536 3392 158588 3398
rect 158536 3334 158588 3340
rect 158628 3392 158680 3398
rect 158628 3334 158680 3340
rect 159088 3052 159140 3058
rect 159088 2994 159140 3000
rect 158444 2848 158496 2854
rect 158444 2790 158496 2796
rect 158628 2848 158680 2854
rect 158628 2790 158680 2796
rect 158456 2582 158484 2790
rect 158444 2576 158496 2582
rect 158444 2518 158496 2524
rect 158444 2440 158496 2446
rect 158444 2382 158496 2388
rect 158456 1057 158484 2382
rect 158536 2032 158588 2038
rect 158536 1974 158588 1980
rect 158548 1426 158576 1974
rect 158536 1420 158588 1426
rect 158536 1362 158588 1368
rect 158640 1329 158668 2790
rect 158996 2372 159048 2378
rect 158996 2314 159048 2320
rect 159008 1970 159036 2314
rect 159100 2106 159128 2994
rect 159088 2100 159140 2106
rect 159088 2042 159140 2048
rect 158996 1964 159048 1970
rect 158996 1906 159048 1912
rect 159192 1902 159220 8842
rect 159560 8430 159588 9454
rect 159652 8974 159680 10066
rect 159916 10056 159968 10062
rect 159916 9998 159968 10004
rect 159928 9518 159956 9998
rect 159916 9512 159968 9518
rect 159916 9454 159968 9460
rect 159640 8968 159692 8974
rect 159640 8910 159692 8916
rect 159928 8430 159956 9454
rect 160008 9376 160060 9382
rect 160008 9318 160060 9324
rect 159548 8424 159600 8430
rect 159362 8392 159418 8401
rect 159272 8356 159324 8362
rect 159548 8366 159600 8372
rect 159916 8424 159968 8430
rect 159916 8366 159968 8372
rect 159362 8327 159418 8336
rect 159272 8298 159324 8304
rect 159284 7886 159312 8298
rect 159272 7880 159324 7886
rect 159272 7822 159324 7828
rect 159376 7750 159404 8327
rect 159454 8120 159510 8129
rect 159454 8055 159456 8064
rect 159508 8055 159510 8064
rect 159456 8026 159508 8032
rect 159364 7744 159416 7750
rect 159364 7686 159416 7692
rect 159456 6452 159508 6458
rect 159456 6394 159508 6400
rect 159468 4622 159496 6394
rect 159456 4616 159508 4622
rect 159456 4558 159508 4564
rect 159364 3528 159416 3534
rect 159364 3470 159416 3476
rect 159376 3126 159404 3470
rect 159364 3120 159416 3126
rect 159364 3062 159416 3068
rect 159364 2848 159416 2854
rect 159364 2790 159416 2796
rect 159272 1964 159324 1970
rect 159272 1906 159324 1912
rect 159180 1896 159232 1902
rect 159180 1838 159232 1844
rect 159284 1358 159312 1906
rect 159272 1352 159324 1358
rect 158626 1320 158682 1329
rect 159272 1294 159324 1300
rect 158626 1255 158682 1264
rect 159376 1193 159404 2790
rect 159456 1420 159508 1426
rect 159560 1408 159588 8366
rect 159824 6112 159876 6118
rect 159824 6054 159876 6060
rect 159836 5710 159864 6054
rect 159732 5704 159784 5710
rect 159732 5646 159784 5652
rect 159824 5704 159876 5710
rect 159824 5646 159876 5652
rect 159744 5234 159772 5646
rect 159732 5228 159784 5234
rect 159732 5170 159784 5176
rect 159744 4622 159772 5170
rect 159640 4616 159692 4622
rect 159640 4558 159692 4564
rect 159732 4616 159784 4622
rect 159732 4558 159784 4564
rect 159652 3670 159680 4558
rect 159640 3664 159692 3670
rect 159640 3606 159692 3612
rect 159928 2446 159956 8366
rect 160020 7886 160048 9318
rect 160008 7880 160060 7886
rect 160008 7822 160060 7828
rect 160480 7410 160508 10474
rect 161112 10396 161164 10402
rect 161112 10338 161164 10344
rect 162124 10396 162176 10402
rect 162124 10338 162176 10344
rect 161124 8906 161152 10338
rect 161940 9988 161992 9994
rect 161940 9930 161992 9936
rect 161204 9580 161256 9586
rect 161204 9522 161256 9528
rect 161296 9580 161348 9586
rect 161296 9522 161348 9528
rect 161112 8900 161164 8906
rect 161112 8842 161164 8848
rect 161124 8430 161152 8842
rect 161112 8424 161164 8430
rect 160926 8392 160982 8401
rect 161112 8366 161164 8372
rect 160926 8327 160982 8336
rect 160744 8288 160796 8294
rect 160744 8230 160796 8236
rect 160756 7886 160784 8230
rect 160940 8090 160968 8327
rect 161018 8120 161074 8129
rect 160928 8084 160980 8090
rect 161018 8055 161020 8064
rect 160928 8026 160980 8032
rect 161072 8055 161074 8064
rect 161020 8026 161072 8032
rect 160744 7880 160796 7886
rect 160744 7822 160796 7828
rect 160468 7404 160520 7410
rect 160468 7346 160520 7352
rect 160376 4480 160428 4486
rect 160376 4422 160428 4428
rect 160284 4208 160336 4214
rect 160284 4150 160336 4156
rect 160008 4072 160060 4078
rect 160008 4014 160060 4020
rect 160020 3641 160048 4014
rect 160100 3732 160152 3738
rect 160100 3674 160152 3680
rect 160006 3632 160062 3641
rect 160006 3567 160062 3576
rect 159916 2440 159968 2446
rect 159916 2382 159968 2388
rect 160008 2440 160060 2446
rect 160008 2382 160060 2388
rect 160020 1970 160048 2382
rect 160008 1964 160060 1970
rect 160008 1906 160060 1912
rect 160112 1408 160140 3674
rect 160296 3194 160324 4150
rect 160388 4010 160416 4422
rect 160376 4004 160428 4010
rect 160376 3946 160428 3952
rect 160284 3188 160336 3194
rect 160284 3130 160336 3136
rect 160284 3052 160336 3058
rect 160284 2994 160336 3000
rect 160296 2106 160324 2994
rect 160836 2304 160888 2310
rect 160836 2246 160888 2252
rect 160192 2100 160244 2106
rect 160192 2042 160244 2048
rect 160284 2100 160336 2106
rect 160284 2042 160336 2048
rect 159508 1380 159588 1408
rect 160020 1380 160140 1408
rect 159456 1362 159508 1368
rect 159362 1184 159418 1193
rect 159362 1119 159418 1128
rect 158442 1048 158498 1057
rect 158442 983 158498 992
rect 158076 400 158128 406
rect 158076 342 158128 348
rect 155316 264 155368 270
rect 155316 206 155368 212
rect 160020 105 160048 1380
rect 160100 1216 160152 1222
rect 160100 1158 160152 1164
rect 160112 649 160140 1158
rect 160204 746 160232 2042
rect 160374 1320 160430 1329
rect 160374 1255 160430 1264
rect 160388 785 160416 1255
rect 160848 1193 160876 2246
rect 161124 1970 161152 8366
rect 161216 8129 161244 9522
rect 161308 8498 161336 9522
rect 161952 9518 161980 9930
rect 161664 9512 161716 9518
rect 161664 9454 161716 9460
rect 161940 9512 161992 9518
rect 161940 9454 161992 9460
rect 161296 8492 161348 8498
rect 161296 8434 161348 8440
rect 161202 8120 161258 8129
rect 161202 8055 161258 8064
rect 161308 7410 161336 8434
rect 161676 8430 161704 9454
rect 161940 8968 161992 8974
rect 161940 8910 161992 8916
rect 161848 8832 161900 8838
rect 161848 8774 161900 8780
rect 161860 8634 161888 8774
rect 161952 8634 161980 8910
rect 161848 8628 161900 8634
rect 161848 8570 161900 8576
rect 161940 8628 161992 8634
rect 161940 8570 161992 8576
rect 162136 8498 162164 10338
rect 162780 9586 162808 10678
rect 164516 10668 164568 10674
rect 164516 10610 164568 10616
rect 163872 9988 163924 9994
rect 163872 9930 163924 9936
rect 162768 9580 162820 9586
rect 162768 9522 162820 9528
rect 162676 9512 162728 9518
rect 162676 9454 162728 9460
rect 162216 9376 162268 9382
rect 162216 9318 162268 9324
rect 162124 8492 162176 8498
rect 162124 8434 162176 8440
rect 161664 8424 161716 8430
rect 161664 8366 161716 8372
rect 161480 8356 161532 8362
rect 161480 8298 161532 8304
rect 161492 7886 161520 8298
rect 161480 7880 161532 7886
rect 161480 7822 161532 7828
rect 161296 7404 161348 7410
rect 161296 7346 161348 7352
rect 161386 7032 161442 7041
rect 161386 6967 161442 6976
rect 161400 6934 161428 6967
rect 161296 6928 161348 6934
rect 161296 6870 161348 6876
rect 161388 6928 161440 6934
rect 161388 6870 161440 6876
rect 161308 6322 161336 6870
rect 161204 6316 161256 6322
rect 161204 6258 161256 6264
rect 161296 6316 161348 6322
rect 161296 6258 161348 6264
rect 161216 3466 161244 6258
rect 161676 6254 161704 8366
rect 161940 8288 161992 8294
rect 161940 8230 161992 8236
rect 161952 7954 161980 8230
rect 161940 7948 161992 7954
rect 161940 7890 161992 7896
rect 162228 7886 162256 9318
rect 162308 8900 162360 8906
rect 162308 8842 162360 8848
rect 162584 8900 162636 8906
rect 162584 8842 162636 8848
rect 162320 8430 162348 8842
rect 162308 8424 162360 8430
rect 162308 8366 162360 8372
rect 162398 8392 162454 8401
rect 162398 8327 162454 8336
rect 162412 8090 162440 8327
rect 162400 8084 162452 8090
rect 162400 8026 162452 8032
rect 162216 7880 162268 7886
rect 162216 7822 162268 7828
rect 162398 7848 162454 7857
rect 162124 7812 162176 7818
rect 162398 7783 162454 7792
rect 162124 7754 162176 7760
rect 162136 7546 162164 7754
rect 162412 7546 162440 7783
rect 162124 7540 162176 7546
rect 162124 7482 162176 7488
rect 162400 7540 162452 7546
rect 162400 7482 162452 7488
rect 162124 6384 162176 6390
rect 162124 6326 162176 6332
rect 161664 6248 161716 6254
rect 161664 6190 161716 6196
rect 161388 4820 161440 4826
rect 161388 4762 161440 4768
rect 161296 4208 161348 4214
rect 161296 4150 161348 4156
rect 161308 3913 161336 4150
rect 161400 4010 161428 4762
rect 161388 4004 161440 4010
rect 161388 3946 161440 3952
rect 161294 3904 161350 3913
rect 161294 3839 161350 3848
rect 161204 3460 161256 3466
rect 161204 3402 161256 3408
rect 161676 2774 161704 6190
rect 162136 5914 162164 6326
rect 162124 5908 162176 5914
rect 162124 5850 162176 5856
rect 161584 2746 161704 2774
rect 161480 2440 161532 2446
rect 161480 2382 161532 2388
rect 161492 2106 161520 2382
rect 161480 2100 161532 2106
rect 161480 2042 161532 2048
rect 161584 1970 161612 2746
rect 161664 2304 161716 2310
rect 161664 2246 161716 2252
rect 162400 2304 162452 2310
rect 162400 2246 162452 2252
rect 161112 1964 161164 1970
rect 161112 1906 161164 1912
rect 161572 1964 161624 1970
rect 161572 1906 161624 1912
rect 161480 1760 161532 1766
rect 161480 1702 161532 1708
rect 161492 1358 161520 1702
rect 161480 1352 161532 1358
rect 161480 1294 161532 1300
rect 161296 1216 161348 1222
rect 160834 1184 160890 1193
rect 161676 1193 161704 2246
rect 162412 2038 162440 2246
rect 162400 2032 162452 2038
rect 162400 1974 162452 1980
rect 162596 1426 162624 8842
rect 162688 8430 162716 9454
rect 162780 8906 162808 9522
rect 163596 9512 163648 9518
rect 163596 9454 163648 9460
rect 162952 9376 163004 9382
rect 162952 9318 163004 9324
rect 162860 8968 162912 8974
rect 162860 8910 162912 8916
rect 162768 8900 162820 8906
rect 162768 8842 162820 8848
rect 162676 8424 162728 8430
rect 162676 8366 162728 8372
rect 162688 1970 162716 8366
rect 162872 6254 162900 8910
rect 162964 7410 162992 9318
rect 163608 8430 163636 9454
rect 163688 9376 163740 9382
rect 163688 9318 163740 9324
rect 163596 8424 163648 8430
rect 163596 8366 163648 8372
rect 163318 8120 163374 8129
rect 163318 8055 163374 8064
rect 163332 7857 163360 8055
rect 163318 7848 163374 7857
rect 163318 7783 163374 7792
rect 162952 7404 163004 7410
rect 162952 7346 163004 7352
rect 162860 6248 162912 6254
rect 162860 6190 162912 6196
rect 163608 4214 163636 8366
rect 163700 7886 163728 9318
rect 163778 9072 163834 9081
rect 163778 9007 163834 9016
rect 163792 8974 163820 9007
rect 163780 8968 163832 8974
rect 163780 8910 163832 8916
rect 163884 8498 163912 9930
rect 164240 9920 164292 9926
rect 164240 9862 164292 9868
rect 163872 8492 163924 8498
rect 163872 8434 163924 8440
rect 163870 8392 163926 8401
rect 163870 8327 163926 8336
rect 163884 8090 163912 8327
rect 164252 8294 164280 9862
rect 164332 9716 164384 9722
rect 164332 9658 164384 9664
rect 164240 8288 164292 8294
rect 164240 8230 164292 8236
rect 163962 8120 164018 8129
rect 163872 8084 163924 8090
rect 163962 8055 163964 8064
rect 163872 8026 163924 8032
rect 164016 8055 164018 8064
rect 163964 8026 164016 8032
rect 163688 7880 163740 7886
rect 163688 7822 163740 7828
rect 164240 4684 164292 4690
rect 164240 4626 164292 4632
rect 163596 4208 163648 4214
rect 163596 4150 163648 4156
rect 163608 1970 163636 4150
rect 164252 3942 164280 4626
rect 164344 4622 164372 9658
rect 164528 9518 164556 10610
rect 164516 9512 164568 9518
rect 164516 9454 164568 9460
rect 164424 9376 164476 9382
rect 164424 9318 164476 9324
rect 164436 7886 164464 9318
rect 164528 8906 164556 9454
rect 164516 8900 164568 8906
rect 164516 8842 164568 8848
rect 164424 7880 164476 7886
rect 164424 7822 164476 7828
rect 164332 4616 164384 4622
rect 164332 4558 164384 4564
rect 164332 4140 164384 4146
rect 164332 4082 164384 4088
rect 164344 3942 164372 4082
rect 164240 3936 164292 3942
rect 164240 3878 164292 3884
rect 164332 3936 164384 3942
rect 164332 3878 164384 3884
rect 163964 2440 164016 2446
rect 163964 2382 164016 2388
rect 163872 2304 163924 2310
rect 163872 2246 163924 2252
rect 162676 1964 162728 1970
rect 162676 1906 162728 1912
rect 163596 1964 163648 1970
rect 163596 1906 163648 1912
rect 162860 1896 162912 1902
rect 162860 1838 162912 1844
rect 162584 1420 162636 1426
rect 162584 1362 162636 1368
rect 162872 1358 162900 1838
rect 163136 1760 163188 1766
rect 162950 1728 163006 1737
rect 163136 1702 163188 1708
rect 162950 1663 163006 1672
rect 162860 1352 162912 1358
rect 162860 1294 162912 1300
rect 162124 1216 162176 1222
rect 161296 1158 161348 1164
rect 161662 1184 161718 1193
rect 160834 1119 160890 1128
rect 160374 776 160430 785
rect 160192 740 160244 746
rect 160374 711 160430 720
rect 160558 776 160614 785
rect 160558 711 160614 720
rect 160192 682 160244 688
rect 160098 640 160154 649
rect 160098 575 160154 584
rect 160572 241 160600 711
rect 161308 377 161336 1158
rect 162124 1158 162176 1164
rect 161662 1119 161718 1128
rect 162136 649 162164 1158
rect 162964 814 162992 1663
rect 163148 1426 163176 1702
rect 163136 1420 163188 1426
rect 163136 1362 163188 1368
rect 163504 1216 163556 1222
rect 163884 1193 163912 2246
rect 163976 2106 164004 2382
rect 163964 2100 164016 2106
rect 163964 2042 164016 2048
rect 164528 1970 164556 8842
rect 165080 8498 165108 10678
rect 165344 10056 165396 10062
rect 165344 9998 165396 10004
rect 166172 10056 166224 10062
rect 166172 9998 166224 10004
rect 165356 9518 165384 9998
rect 165344 9512 165396 9518
rect 165344 9454 165396 9460
rect 165804 9512 165856 9518
rect 165804 9454 165856 9460
rect 165160 9376 165212 9382
rect 165160 9318 165212 9324
rect 165068 8492 165120 8498
rect 165068 8434 165120 8440
rect 165068 8356 165120 8362
rect 165068 8298 165120 8304
rect 164700 8288 164752 8294
rect 164700 8230 164752 8236
rect 164712 8022 164740 8230
rect 164700 8016 164752 8022
rect 164700 7958 164752 7964
rect 165080 2774 165108 8298
rect 165172 7886 165200 9318
rect 165356 8430 165384 9454
rect 165816 8838 165844 9454
rect 165896 9376 165948 9382
rect 165896 9318 165948 9324
rect 165804 8832 165856 8838
rect 165804 8774 165856 8780
rect 165344 8424 165396 8430
rect 165250 8392 165306 8401
rect 165344 8366 165396 8372
rect 165250 8327 165306 8336
rect 165160 7880 165212 7886
rect 165160 7822 165212 7828
rect 165264 7750 165292 8327
rect 165342 8120 165398 8129
rect 165342 8055 165344 8064
rect 165396 8055 165398 8064
rect 165344 8026 165396 8032
rect 165908 7886 165936 9318
rect 166184 8974 166212 9998
rect 166460 8974 166488 10814
rect 177580 10804 177632 10810
rect 177580 10746 177632 10752
rect 219900 10804 219952 10810
rect 219900 10746 219952 10752
rect 172242 10568 172298 10577
rect 172242 10503 172298 10512
rect 171690 10296 171746 10305
rect 166724 10260 166776 10266
rect 171690 10231 171746 10240
rect 166724 10202 166776 10208
rect 166736 9586 166764 10202
rect 168378 9752 168434 9761
rect 168378 9687 168380 9696
rect 168432 9687 168434 9696
rect 169482 9752 169538 9761
rect 169482 9687 169538 9696
rect 168380 9658 168432 9664
rect 168748 9648 168800 9654
rect 168748 9590 168800 9596
rect 166540 9580 166592 9586
rect 166540 9522 166592 9528
rect 166724 9580 166776 9586
rect 166724 9522 166776 9528
rect 166908 9580 166960 9586
rect 166908 9522 166960 9528
rect 166172 8968 166224 8974
rect 166448 8968 166500 8974
rect 166172 8910 166224 8916
rect 166368 8928 166448 8956
rect 166368 8498 166396 8928
rect 166448 8910 166500 8916
rect 166552 8498 166580 9522
rect 166724 9376 166776 9382
rect 166724 9318 166776 9324
rect 166356 8492 166408 8498
rect 166356 8434 166408 8440
rect 166540 8492 166592 8498
rect 166540 8434 166592 8440
rect 165896 7880 165948 7886
rect 165896 7822 165948 7828
rect 165252 7744 165304 7750
rect 165252 7686 165304 7692
rect 165712 6248 165764 6254
rect 165712 6190 165764 6196
rect 165620 5364 165672 5370
rect 165620 5306 165672 5312
rect 165632 5030 165660 5306
rect 165620 5024 165672 5030
rect 165620 4966 165672 4972
rect 165724 3058 165752 6190
rect 165988 4480 166040 4486
rect 165988 4422 166040 4428
rect 166000 4282 166028 4422
rect 165988 4276 166040 4282
rect 165988 4218 166040 4224
rect 165712 3052 165764 3058
rect 165712 2994 165764 3000
rect 166368 2774 166396 8434
rect 166538 8392 166594 8401
rect 166538 8327 166594 8336
rect 166552 7750 166580 8327
rect 166632 8288 166684 8294
rect 166632 8230 166684 8236
rect 166644 8022 166672 8230
rect 166632 8016 166684 8022
rect 166632 7958 166684 7964
rect 166540 7744 166592 7750
rect 166540 7686 166592 7692
rect 166736 7410 166764 9318
rect 166920 8514 166948 9522
rect 167092 9512 167144 9518
rect 167092 9454 167144 9460
rect 167104 8906 167132 9454
rect 168760 8974 168788 9590
rect 169208 9580 169260 9586
rect 169208 9522 169260 9528
rect 168748 8968 168800 8974
rect 168748 8910 168800 8916
rect 168932 8968 168984 8974
rect 168932 8910 168984 8916
rect 169024 8968 169076 8974
rect 169024 8910 169076 8916
rect 167092 8900 167144 8906
rect 167092 8842 167144 8848
rect 167828 8900 167880 8906
rect 167828 8842 167880 8848
rect 166920 8498 167040 8514
rect 166816 8492 166868 8498
rect 166816 8434 166868 8440
rect 166908 8492 167040 8498
rect 166960 8486 167040 8492
rect 166908 8434 166960 8440
rect 166828 7954 166856 8434
rect 166906 8392 166962 8401
rect 166906 8327 166962 8336
rect 166816 7948 166868 7954
rect 166816 7890 166868 7896
rect 166920 7546 166948 8327
rect 166908 7540 166960 7546
rect 166908 7482 166960 7488
rect 167012 7426 167040 8486
rect 166724 7404 166776 7410
rect 166724 7346 166776 7352
rect 166920 7398 167040 7426
rect 165080 2746 165200 2774
rect 165172 1970 165200 2746
rect 166276 2746 166396 2774
rect 165620 2440 165672 2446
rect 165620 2382 165672 2388
rect 165804 2440 165856 2446
rect 165804 2382 165856 2388
rect 165252 2304 165304 2310
rect 165252 2246 165304 2252
rect 164516 1964 164568 1970
rect 164516 1906 164568 1912
rect 165160 1964 165212 1970
rect 165160 1906 165212 1912
rect 164424 1760 164476 1766
rect 164424 1702 164476 1708
rect 164436 1358 164464 1702
rect 164424 1352 164476 1358
rect 164424 1294 164476 1300
rect 164608 1216 164660 1222
rect 163504 1158 163556 1164
rect 163870 1184 163926 1193
rect 162952 808 163004 814
rect 162952 750 163004 756
rect 163516 649 163544 1158
rect 165264 1193 165292 2246
rect 165632 2106 165660 2382
rect 165816 2106 165844 2382
rect 165988 2304 166040 2310
rect 165988 2246 166040 2252
rect 165620 2100 165672 2106
rect 165620 2042 165672 2048
rect 165804 2100 165856 2106
rect 165804 2042 165856 2048
rect 166000 1193 166028 2246
rect 166276 1970 166304 2746
rect 166540 2576 166592 2582
rect 166540 2518 166592 2524
rect 166264 1964 166316 1970
rect 166264 1906 166316 1912
rect 166552 1902 166580 2518
rect 166816 2304 166868 2310
rect 166816 2246 166868 2252
rect 166540 1896 166592 1902
rect 166540 1838 166592 1844
rect 166828 1193 166856 2246
rect 166920 1426 166948 7398
rect 167104 7290 167132 8842
rect 167840 7886 167868 8842
rect 168944 8838 168972 8910
rect 168840 8832 168892 8838
rect 168840 8774 168892 8780
rect 168932 8832 168984 8838
rect 168932 8774 168984 8780
rect 168656 8424 168708 8430
rect 168656 8366 168708 8372
rect 167828 7880 167880 7886
rect 167828 7822 167880 7828
rect 167012 7262 167132 7290
rect 167012 2774 167040 7262
rect 167736 6656 167788 6662
rect 167736 6598 167788 6604
rect 167748 6186 167776 6598
rect 167736 6180 167788 6186
rect 167736 6122 167788 6128
rect 167460 5568 167512 5574
rect 167460 5510 167512 5516
rect 167472 5234 167500 5510
rect 167460 5228 167512 5234
rect 167460 5170 167512 5176
rect 167184 4820 167236 4826
rect 167184 4762 167236 4768
rect 167196 4622 167224 4762
rect 167301 4684 167353 4690
rect 167288 4632 167301 4672
rect 167288 4626 167353 4632
rect 167184 4616 167236 4622
rect 167184 4558 167236 4564
rect 167288 4486 167316 4626
rect 167472 4622 167500 5170
rect 167460 4616 167512 4622
rect 167460 4558 167512 4564
rect 167184 4480 167236 4486
rect 167184 4422 167236 4428
rect 167276 4480 167328 4486
rect 167276 4422 167328 4428
rect 167196 4214 167224 4422
rect 167288 4282 167316 4422
rect 167276 4276 167328 4282
rect 167276 4218 167328 4224
rect 167368 4276 167420 4282
rect 167368 4218 167420 4224
rect 167184 4208 167236 4214
rect 167184 4150 167236 4156
rect 167380 3942 167408 4218
rect 167472 3942 167500 4558
rect 167748 4146 167776 6122
rect 167736 4140 167788 4146
rect 167736 4082 167788 4088
rect 167368 3936 167420 3942
rect 167368 3878 167420 3884
rect 167460 3936 167512 3942
rect 167460 3878 167512 3884
rect 167736 3392 167788 3398
rect 167736 3334 167788 3340
rect 167012 2746 167132 2774
rect 167104 1970 167132 2746
rect 167460 2440 167512 2446
rect 167460 2382 167512 2388
rect 167472 2106 167500 2382
rect 167748 2378 167776 3334
rect 167736 2372 167788 2378
rect 167736 2314 167788 2320
rect 167460 2100 167512 2106
rect 167460 2042 167512 2048
rect 167184 2032 167236 2038
rect 167184 1974 167236 1980
rect 167092 1964 167144 1970
rect 167092 1906 167144 1912
rect 166908 1420 166960 1426
rect 166908 1362 166960 1368
rect 167000 1420 167052 1426
rect 167000 1362 167052 1368
rect 167012 1329 167040 1362
rect 167196 1358 167224 1974
rect 167840 1902 167868 7822
rect 168668 7546 168696 8366
rect 168852 8362 168880 8774
rect 168932 8424 168984 8430
rect 168932 8366 168984 8372
rect 168840 8356 168892 8362
rect 168840 8298 168892 8304
rect 168944 7886 168972 8366
rect 169036 8022 169064 8910
rect 169220 8022 169248 9522
rect 169496 9518 169524 9687
rect 171232 9648 171284 9654
rect 171232 9590 171284 9596
rect 169484 9512 169536 9518
rect 171140 9512 171192 9518
rect 169484 9454 169536 9460
rect 169588 9450 169892 9466
rect 171140 9454 171192 9460
rect 169576 9444 169904 9450
rect 169628 9438 169852 9444
rect 169576 9386 169628 9392
rect 169852 9386 169904 9392
rect 169668 9376 169720 9382
rect 169668 9318 169720 9324
rect 169680 9110 169708 9318
rect 169942 9276 170250 9285
rect 169942 9274 169948 9276
rect 170004 9274 170028 9276
rect 170084 9274 170108 9276
rect 170164 9274 170188 9276
rect 170244 9274 170250 9276
rect 170004 9222 170006 9274
rect 170186 9222 170188 9274
rect 169942 9220 169948 9222
rect 170004 9220 170028 9222
rect 170084 9220 170108 9222
rect 170164 9220 170188 9222
rect 170244 9220 170250 9222
rect 169758 9208 169814 9217
rect 169942 9211 170250 9220
rect 169758 9143 169814 9152
rect 169772 9110 169800 9143
rect 169668 9104 169720 9110
rect 169668 9046 169720 9052
rect 169760 9104 169812 9110
rect 169760 9046 169812 9052
rect 171048 8832 171100 8838
rect 171048 8774 171100 8780
rect 169760 8424 169812 8430
rect 169760 8366 169812 8372
rect 169668 8356 169720 8362
rect 169668 8298 169720 8304
rect 169680 8022 169708 8298
rect 169024 8016 169076 8022
rect 169024 7958 169076 7964
rect 169208 8016 169260 8022
rect 169208 7958 169260 7964
rect 169668 8016 169720 8022
rect 169668 7958 169720 7964
rect 169772 7954 169800 8366
rect 171060 8265 171088 8774
rect 171046 8256 171102 8265
rect 169942 8188 170250 8197
rect 171046 8191 171102 8200
rect 169942 8186 169948 8188
rect 170004 8186 170028 8188
rect 170084 8186 170108 8188
rect 170164 8186 170188 8188
rect 170244 8186 170250 8188
rect 170004 8134 170006 8186
rect 170186 8134 170188 8186
rect 169942 8132 169948 8134
rect 170004 8132 170028 8134
rect 170084 8132 170108 8134
rect 170164 8132 170188 8134
rect 170244 8132 170250 8134
rect 169942 8123 170250 8132
rect 169760 7948 169812 7954
rect 169760 7890 169812 7896
rect 168932 7880 168984 7886
rect 168932 7822 168984 7828
rect 170588 7880 170640 7886
rect 170588 7822 170640 7828
rect 170770 7848 170826 7857
rect 169668 7744 169720 7750
rect 169668 7686 169720 7692
rect 168656 7540 168708 7546
rect 168656 7482 168708 7488
rect 169024 7404 169076 7410
rect 169024 7346 169076 7352
rect 168286 6760 168342 6769
rect 168286 6695 168342 6704
rect 168012 6384 168064 6390
rect 168012 6326 168064 6332
rect 167920 5364 167972 5370
rect 167920 5306 167972 5312
rect 167932 5166 167960 5306
rect 167920 5160 167972 5166
rect 167920 5102 167972 5108
rect 168024 4214 168052 6326
rect 168300 5817 168328 6695
rect 168840 6656 168892 6662
rect 168840 6598 168892 6604
rect 168656 6248 168708 6254
rect 168852 6225 168880 6598
rect 168656 6190 168708 6196
rect 168838 6216 168894 6225
rect 168286 5808 168342 5817
rect 168286 5743 168342 5752
rect 168300 5710 168328 5743
rect 168288 5704 168340 5710
rect 168288 5646 168340 5652
rect 168668 5642 168696 6190
rect 169036 6186 169064 7346
rect 169574 7168 169630 7177
rect 169574 7103 169630 7112
rect 168838 6151 168894 6160
rect 169024 6180 169076 6186
rect 168852 5710 168880 6151
rect 169024 6122 169076 6128
rect 169206 5808 169262 5817
rect 169206 5743 169262 5752
rect 169220 5710 169248 5743
rect 168840 5704 168892 5710
rect 168840 5646 168892 5652
rect 169208 5704 169260 5710
rect 169208 5646 169260 5652
rect 168656 5636 168708 5642
rect 168656 5578 168708 5584
rect 169392 5568 169444 5574
rect 169392 5510 169444 5516
rect 168104 5160 168156 5166
rect 168288 5160 168340 5166
rect 168104 5102 168156 5108
rect 168208 5108 168288 5114
rect 168208 5102 168340 5108
rect 168116 4826 168144 5102
rect 168208 5086 168328 5102
rect 168104 4820 168156 4826
rect 168104 4762 168156 4768
rect 168012 4208 168064 4214
rect 168012 4150 168064 4156
rect 168208 4078 168236 5086
rect 168288 5024 168340 5030
rect 168288 4966 168340 4972
rect 168300 4690 168328 4966
rect 168288 4684 168340 4690
rect 168288 4626 168340 4632
rect 169404 4622 169432 5510
rect 169588 5234 169616 7103
rect 169680 5778 169708 7686
rect 169942 7100 170250 7109
rect 169942 7098 169948 7100
rect 170004 7098 170028 7100
rect 170084 7098 170108 7100
rect 170164 7098 170188 7100
rect 170244 7098 170250 7100
rect 170004 7046 170006 7098
rect 170186 7046 170188 7098
rect 169942 7044 169948 7046
rect 170004 7044 170028 7046
rect 170084 7044 170108 7046
rect 170164 7044 170188 7046
rect 170244 7044 170250 7046
rect 169942 7035 170250 7044
rect 170600 6633 170628 7822
rect 170770 7783 170826 7792
rect 170586 6624 170642 6633
rect 170586 6559 170642 6568
rect 169758 6352 169814 6361
rect 169758 6287 169760 6296
rect 169812 6287 169814 6296
rect 169760 6258 169812 6264
rect 170784 6089 170812 7783
rect 171152 7449 171180 9454
rect 171138 7440 171194 7449
rect 171138 7375 171194 7384
rect 171244 6322 171272 9590
rect 171704 9586 171732 10231
rect 172256 9586 172284 10503
rect 173990 10432 174046 10441
rect 173990 10367 174046 10376
rect 173898 10296 173954 10305
rect 173898 10231 173954 10240
rect 171692 9580 171744 9586
rect 171692 9522 171744 9528
rect 172244 9580 172296 9586
rect 172244 9522 172296 9528
rect 172612 9512 172664 9518
rect 172612 9454 172664 9460
rect 171876 9036 171928 9042
rect 171876 8978 171928 8984
rect 171888 8566 171916 8978
rect 171876 8560 171928 8566
rect 171876 8502 171928 8508
rect 171784 8016 171836 8022
rect 171784 7958 171836 7964
rect 171796 7342 171824 7958
rect 172624 7886 172652 9454
rect 173912 8974 173940 10231
rect 174004 9586 174032 10367
rect 174268 10328 174320 10334
rect 174268 10270 174320 10276
rect 174450 10296 174506 10305
rect 173992 9580 174044 9586
rect 173992 9522 174044 9528
rect 174280 9110 174308 10270
rect 174450 10231 174506 10240
rect 175186 10296 175242 10305
rect 175186 10231 175242 10240
rect 175922 10296 175978 10305
rect 175922 10231 175978 10240
rect 176750 10296 176806 10305
rect 176750 10231 176806 10240
rect 177486 10296 177542 10305
rect 177486 10231 177542 10240
rect 174464 9654 174492 10231
rect 174452 9648 174504 9654
rect 174452 9590 174504 9596
rect 174268 9104 174320 9110
rect 174268 9046 174320 9052
rect 175200 8974 175228 10231
rect 175556 10192 175608 10198
rect 175556 10134 175608 10140
rect 175568 9654 175596 10134
rect 175556 9648 175608 9654
rect 175556 9590 175608 9596
rect 175936 9586 175964 10231
rect 175924 9580 175976 9586
rect 175924 9522 175976 9528
rect 175556 9376 175608 9382
rect 175556 9318 175608 9324
rect 175568 9178 175596 9318
rect 175556 9172 175608 9178
rect 175556 9114 175608 9120
rect 175280 9104 175332 9110
rect 175280 9046 175332 9052
rect 173900 8968 173952 8974
rect 173900 8910 173952 8916
rect 175188 8968 175240 8974
rect 175188 8910 175240 8916
rect 172704 8832 172756 8838
rect 172704 8774 172756 8780
rect 172612 7880 172664 7886
rect 172612 7822 172664 7828
rect 172518 7712 172574 7721
rect 172518 7647 172574 7656
rect 171784 7336 171836 7342
rect 171784 7278 171836 7284
rect 172532 7206 172560 7647
rect 172520 7200 172572 7206
rect 172520 7142 172572 7148
rect 172610 7168 172666 7177
rect 172610 7103 172666 7112
rect 171232 6316 171284 6322
rect 171232 6258 171284 6264
rect 170770 6080 170826 6089
rect 169942 6012 170250 6021
rect 170770 6015 170826 6024
rect 169942 6010 169948 6012
rect 170004 6010 170028 6012
rect 170084 6010 170108 6012
rect 170164 6010 170188 6012
rect 170244 6010 170250 6012
rect 170004 5958 170006 6010
rect 170186 5958 170188 6010
rect 169942 5956 169948 5958
rect 170004 5956 170028 5958
rect 170084 5956 170108 5958
rect 170164 5956 170188 5958
rect 170244 5956 170250 5958
rect 169942 5947 170250 5956
rect 169668 5772 169720 5778
rect 169668 5714 169720 5720
rect 169852 5704 169904 5710
rect 169852 5646 169904 5652
rect 172518 5672 172574 5681
rect 169576 5228 169628 5234
rect 169576 5170 169628 5176
rect 169392 4616 169444 4622
rect 169392 4558 169444 4564
rect 169588 4185 169616 5170
rect 169864 5166 169892 5646
rect 172518 5607 172574 5616
rect 171048 5568 171100 5574
rect 171048 5510 171100 5516
rect 171060 5370 171088 5510
rect 171048 5364 171100 5370
rect 171048 5306 171100 5312
rect 169852 5160 169904 5166
rect 169852 5102 169904 5108
rect 169864 4758 169892 5102
rect 172532 5030 172560 5607
rect 172624 5574 172652 7103
rect 172612 5568 172664 5574
rect 172612 5510 172664 5516
rect 172520 5024 172572 5030
rect 172520 4966 172572 4972
rect 169942 4924 170250 4933
rect 169942 4922 169948 4924
rect 170004 4922 170028 4924
rect 170084 4922 170108 4924
rect 170164 4922 170188 4924
rect 170244 4922 170250 4924
rect 170004 4870 170006 4922
rect 170186 4870 170188 4922
rect 169942 4868 169948 4870
rect 170004 4868 170028 4870
rect 170084 4868 170108 4870
rect 170164 4868 170188 4870
rect 170244 4868 170250 4870
rect 169942 4859 170250 4868
rect 169852 4752 169904 4758
rect 169852 4694 169904 4700
rect 170864 4752 170916 4758
rect 170864 4694 170916 4700
rect 169852 4548 169904 4554
rect 169852 4490 169904 4496
rect 169666 4448 169722 4457
rect 169666 4383 169722 4392
rect 169574 4176 169630 4185
rect 169574 4111 169630 4120
rect 168196 4072 168248 4078
rect 168196 4014 168248 4020
rect 168288 3936 168340 3942
rect 168288 3878 168340 3884
rect 168300 3534 168328 3878
rect 168380 3596 168432 3602
rect 168380 3538 168432 3544
rect 168288 3528 168340 3534
rect 168288 3470 168340 3476
rect 167920 2984 167972 2990
rect 167920 2926 167972 2932
rect 167932 2446 167960 2926
rect 168392 2582 168420 3538
rect 169680 2774 169708 4383
rect 169680 2746 169800 2774
rect 168380 2576 168432 2582
rect 168380 2518 168432 2524
rect 167920 2440 167972 2446
rect 167920 2382 167972 2388
rect 168012 2440 168064 2446
rect 168012 2382 168064 2388
rect 168288 2440 168340 2446
rect 168288 2382 168340 2388
rect 168024 1970 168052 2382
rect 168300 2310 168328 2382
rect 168196 2304 168248 2310
rect 168196 2246 168248 2252
rect 168288 2304 168340 2310
rect 168288 2246 168340 2252
rect 168012 1964 168064 1970
rect 168012 1906 168064 1912
rect 167828 1896 167880 1902
rect 167828 1838 167880 1844
rect 168208 1358 168236 2246
rect 169772 1970 169800 2746
rect 169760 1964 169812 1970
rect 169760 1906 169812 1912
rect 168380 1760 168432 1766
rect 168380 1702 168432 1708
rect 168392 1465 168420 1702
rect 168378 1456 168434 1465
rect 169864 1426 169892 4490
rect 170876 4282 170904 4694
rect 170864 4276 170916 4282
rect 170864 4218 170916 4224
rect 169942 3836 170250 3845
rect 169942 3834 169948 3836
rect 170004 3834 170028 3836
rect 170084 3834 170108 3836
rect 170164 3834 170188 3836
rect 170244 3834 170250 3836
rect 170004 3782 170006 3834
rect 170186 3782 170188 3834
rect 169942 3780 169948 3782
rect 170004 3780 170028 3782
rect 170084 3780 170108 3782
rect 170164 3780 170188 3782
rect 170244 3780 170250 3782
rect 169942 3771 170250 3780
rect 172716 3738 172744 8774
rect 175292 5409 175320 9046
rect 176764 8974 176792 10231
rect 176844 9920 176896 9926
rect 176844 9862 176896 9868
rect 176856 9178 176884 9862
rect 176844 9172 176896 9178
rect 176844 9114 176896 9120
rect 177500 8974 177528 10231
rect 177592 9178 177620 10746
rect 217876 10736 217928 10742
rect 217876 10678 217928 10684
rect 202328 10668 202380 10674
rect 202328 10610 202380 10616
rect 180708 10600 180760 10606
rect 180522 10568 180578 10577
rect 180708 10542 180760 10548
rect 200120 10600 200172 10606
rect 200120 10542 200172 10548
rect 180522 10503 180578 10512
rect 178040 10464 178092 10470
rect 178040 10406 178092 10412
rect 177946 10296 178002 10305
rect 177946 10231 178002 10240
rect 177960 9586 177988 10231
rect 178052 9586 178080 10406
rect 179142 10296 179198 10305
rect 179142 10231 179198 10240
rect 180430 10296 180486 10305
rect 180430 10231 180486 10240
rect 179156 9586 179184 10231
rect 177948 9580 178000 9586
rect 177948 9522 178000 9528
rect 178040 9580 178092 9586
rect 178040 9522 178092 9528
rect 179144 9580 179196 9586
rect 179144 9522 179196 9528
rect 178408 9376 178460 9382
rect 178408 9318 178460 9324
rect 177580 9172 177632 9178
rect 177580 9114 177632 9120
rect 176752 8968 176804 8974
rect 176752 8910 176804 8916
rect 177488 8968 177540 8974
rect 177488 8910 177540 8916
rect 177672 8832 177724 8838
rect 177672 8774 177724 8780
rect 177684 8090 177712 8774
rect 177672 8084 177724 8090
rect 177672 8026 177724 8032
rect 175278 5400 175334 5409
rect 175278 5335 175334 5344
rect 178420 4729 178448 9318
rect 180444 8974 180472 10231
rect 180536 9586 180564 10503
rect 180720 9586 180748 10542
rect 182088 10532 182140 10538
rect 182088 10474 182140 10480
rect 193312 10532 193364 10538
rect 193312 10474 193364 10480
rect 181810 10432 181866 10441
rect 181810 10367 181866 10376
rect 181824 9586 181852 10367
rect 181902 10296 181958 10305
rect 181902 10231 181958 10240
rect 180524 9580 180576 9586
rect 180524 9522 180576 9528
rect 180708 9580 180760 9586
rect 180708 9522 180760 9528
rect 181812 9580 181864 9586
rect 181812 9522 181864 9528
rect 181916 8974 181944 10231
rect 182100 9110 182128 10474
rect 191286 10432 191342 10441
rect 191286 10367 191342 10376
rect 192850 10432 192906 10441
rect 192850 10367 192906 10376
rect 182546 10296 182602 10305
rect 182546 10231 182602 10240
rect 183282 10296 183338 10305
rect 183282 10231 183338 10240
rect 184294 10296 184350 10305
rect 184294 10231 184350 10240
rect 184754 10296 184810 10305
rect 184754 10231 184810 10240
rect 185490 10296 185546 10305
rect 185490 10231 185546 10240
rect 186226 10296 186282 10305
rect 186226 10231 186282 10240
rect 186962 10296 187018 10305
rect 186962 10231 187018 10240
rect 187698 10296 187754 10305
rect 187698 10231 187754 10240
rect 188618 10296 188674 10305
rect 188618 10231 188674 10240
rect 189446 10296 189502 10305
rect 189446 10231 189502 10240
rect 189906 10296 189962 10305
rect 189906 10231 189962 10240
rect 182560 9586 182588 10231
rect 183296 9586 183324 10231
rect 182548 9580 182600 9586
rect 182548 9522 182600 9528
rect 183284 9580 183336 9586
rect 183284 9522 183336 9528
rect 182088 9104 182140 9110
rect 182088 9046 182140 9052
rect 184308 9042 184336 10231
rect 184572 9512 184624 9518
rect 184572 9454 184624 9460
rect 184584 9178 184612 9454
rect 184572 9172 184624 9178
rect 184572 9114 184624 9120
rect 184768 9042 184796 10231
rect 185504 9586 185532 10231
rect 185492 9580 185544 9586
rect 185492 9522 185544 9528
rect 184848 9444 184900 9450
rect 184848 9386 184900 9392
rect 184296 9036 184348 9042
rect 184296 8978 184348 8984
rect 184756 9036 184808 9042
rect 184756 8978 184808 8984
rect 180432 8968 180484 8974
rect 180432 8910 180484 8916
rect 181904 8968 181956 8974
rect 181904 8910 181956 8916
rect 182088 8832 182140 8838
rect 182088 8774 182140 8780
rect 179418 8256 179474 8265
rect 179418 8191 179474 8200
rect 179432 7546 179460 8191
rect 182100 8022 182128 8774
rect 182088 8016 182140 8022
rect 182088 7958 182140 7964
rect 179420 7540 179472 7546
rect 179420 7482 179472 7488
rect 184860 6458 184888 9386
rect 186240 9042 186268 10231
rect 186412 9512 186464 9518
rect 186412 9454 186464 9460
rect 186320 9376 186372 9382
rect 186320 9318 186372 9324
rect 186228 9036 186280 9042
rect 186228 8978 186280 8984
rect 185860 8968 185912 8974
rect 185860 8910 185912 8916
rect 185872 6497 185900 8910
rect 185858 6488 185914 6497
rect 184848 6452 184900 6458
rect 185858 6423 185914 6432
rect 184848 6394 184900 6400
rect 185492 6180 185544 6186
rect 185492 6122 185544 6128
rect 185504 5778 185532 6122
rect 185492 5772 185544 5778
rect 185492 5714 185544 5720
rect 184572 5024 184624 5030
rect 184572 4966 184624 4972
rect 178406 4720 178462 4729
rect 178406 4655 178462 4664
rect 173806 4312 173862 4321
rect 173806 4247 173862 4256
rect 176660 4276 176712 4282
rect 172704 3732 172756 3738
rect 172704 3674 172756 3680
rect 171784 3596 171836 3602
rect 171784 3538 171836 3544
rect 171796 3194 171824 3538
rect 171784 3188 171836 3194
rect 171784 3130 171836 3136
rect 170312 3052 170364 3058
rect 170312 2994 170364 3000
rect 169942 2748 170250 2757
rect 169942 2746 169948 2748
rect 170004 2746 170028 2748
rect 170084 2746 170108 2748
rect 170164 2746 170188 2748
rect 170244 2746 170250 2748
rect 170004 2694 170006 2746
rect 170186 2694 170188 2746
rect 169942 2692 169948 2694
rect 170004 2692 170028 2694
rect 170084 2692 170108 2694
rect 170164 2692 170188 2694
rect 170244 2692 170250 2694
rect 169942 2683 170250 2692
rect 169942 1660 170250 1669
rect 169942 1658 169948 1660
rect 170004 1658 170028 1660
rect 170084 1658 170108 1660
rect 170164 1658 170188 1660
rect 170244 1658 170250 1660
rect 170004 1606 170006 1658
rect 170186 1606 170188 1658
rect 169942 1604 169948 1606
rect 170004 1604 170028 1606
rect 170084 1604 170108 1606
rect 170164 1604 170188 1606
rect 170244 1604 170250 1606
rect 169942 1595 170250 1604
rect 168378 1391 168434 1400
rect 169852 1420 169904 1426
rect 169852 1362 169904 1368
rect 167184 1352 167236 1358
rect 166998 1320 167054 1329
rect 167184 1294 167236 1300
rect 168196 1352 168248 1358
rect 168196 1294 168248 1300
rect 166998 1255 167054 1264
rect 167920 1216 167972 1222
rect 164608 1158 164660 1164
rect 165250 1184 165306 1193
rect 163870 1119 163926 1128
rect 164620 649 164648 1158
rect 165250 1119 165306 1128
rect 165986 1184 166042 1193
rect 165986 1119 166042 1128
rect 166814 1184 166870 1193
rect 167920 1158 167972 1164
rect 169024 1216 169076 1222
rect 169024 1158 169076 1164
rect 166814 1119 166870 1128
rect 162122 640 162178 649
rect 162122 575 162178 584
rect 163502 640 163558 649
rect 163502 575 163558 584
rect 164606 640 164662 649
rect 164606 575 164662 584
rect 167932 377 167960 1158
rect 168378 1048 168434 1057
rect 168378 983 168434 992
rect 168392 678 168420 983
rect 168380 672 168432 678
rect 169036 649 169064 1158
rect 170324 1057 170352 2994
rect 172428 2372 172480 2378
rect 172428 2314 172480 2320
rect 171692 1420 171744 1426
rect 171692 1362 171744 1368
rect 170310 1048 170366 1057
rect 170310 983 170366 992
rect 171704 649 171732 1362
rect 172244 1352 172296 1358
rect 172244 1294 172296 1300
rect 172256 649 172284 1294
rect 168380 614 168432 620
rect 169022 640 169078 649
rect 169022 575 169078 584
rect 171690 640 171746 649
rect 171690 575 171746 584
rect 172242 640 172298 649
rect 172242 575 172298 584
rect 172440 474 172468 2314
rect 173820 2038 173848 4247
rect 176660 4218 176712 4224
rect 176672 3097 176700 4218
rect 182088 3664 182140 3670
rect 182088 3606 182140 3612
rect 176658 3088 176714 3097
rect 176658 3023 176714 3032
rect 176660 2440 176712 2446
rect 176660 2382 176712 2388
rect 176936 2440 176988 2446
rect 176936 2382 176988 2388
rect 179604 2440 179656 2446
rect 179604 2382 179656 2388
rect 181812 2440 181864 2446
rect 181812 2382 181864 2388
rect 173808 2032 173860 2038
rect 173808 1974 173860 1980
rect 172980 1896 173032 1902
rect 172980 1838 173032 1844
rect 174452 1896 174504 1902
rect 174728 1896 174780 1902
rect 174452 1838 174504 1844
rect 174726 1864 174728 1873
rect 176568 1896 176620 1902
rect 174780 1864 174782 1873
rect 172520 1352 172572 1358
rect 172520 1294 172572 1300
rect 172428 468 172480 474
rect 172428 410 172480 416
rect 172532 406 172560 1294
rect 172992 649 173020 1838
rect 173900 1352 173952 1358
rect 173900 1294 173952 1300
rect 174268 1352 174320 1358
rect 174268 1294 174320 1300
rect 173912 649 173940 1294
rect 172978 640 173034 649
rect 172978 575 173034 584
rect 173898 640 173954 649
rect 173898 575 173954 584
rect 172520 400 172572 406
rect 161294 368 161350 377
rect 161294 303 161350 312
rect 167918 368 167974 377
rect 172520 342 172572 348
rect 167918 303 167974 312
rect 174280 241 174308 1294
rect 174464 649 174492 1838
rect 176568 1838 176620 1844
rect 174726 1799 174782 1808
rect 175280 1352 175332 1358
rect 175280 1294 175332 1300
rect 175292 649 175320 1294
rect 174450 640 174506 649
rect 174450 575 174506 584
rect 175278 640 175334 649
rect 175278 575 175334 584
rect 176580 513 176608 1838
rect 176672 649 176700 2382
rect 176842 2272 176898 2281
rect 176842 2207 176898 2216
rect 176856 1970 176884 2207
rect 176844 1964 176896 1970
rect 176844 1906 176896 1912
rect 176948 1562 176976 2382
rect 179418 2136 179474 2145
rect 179418 2071 179474 2080
rect 179432 1970 179460 2071
rect 179420 1964 179472 1970
rect 179420 1906 179472 1912
rect 177856 1896 177908 1902
rect 177856 1838 177908 1844
rect 178132 1896 178184 1902
rect 178132 1838 178184 1844
rect 179144 1896 179196 1902
rect 179144 1838 179196 1844
rect 176936 1556 176988 1562
rect 176936 1498 176988 1504
rect 177028 1556 177080 1562
rect 177028 1498 177080 1504
rect 176844 1352 176896 1358
rect 176844 1294 176896 1300
rect 176658 640 176714 649
rect 176658 575 176714 584
rect 176566 504 176622 513
rect 176566 439 176622 448
rect 176856 377 176884 1294
rect 177040 610 177068 1498
rect 177868 649 177896 1838
rect 178144 1494 178172 1838
rect 178132 1488 178184 1494
rect 178132 1430 178184 1436
rect 178500 1352 178552 1358
rect 178500 1294 178552 1300
rect 178512 649 178540 1294
rect 179156 649 179184 1838
rect 179420 1352 179472 1358
rect 179420 1294 179472 1300
rect 179432 1018 179460 1294
rect 179420 1012 179472 1018
rect 179420 954 179472 960
rect 179616 649 179644 2382
rect 181720 1896 181772 1902
rect 181720 1838 181772 1844
rect 180340 1352 180392 1358
rect 180340 1294 180392 1300
rect 180352 649 180380 1294
rect 180522 1048 180578 1057
rect 180522 983 180578 992
rect 180536 649 180564 983
rect 177854 640 177910 649
rect 177028 604 177080 610
rect 177854 575 177910 584
rect 178498 640 178554 649
rect 178498 575 178554 584
rect 179142 640 179198 649
rect 179142 575 179198 584
rect 179602 640 179658 649
rect 179602 575 179658 584
rect 180338 640 180394 649
rect 180338 575 180394 584
rect 180522 640 180578 649
rect 180522 575 180578 584
rect 177028 546 177080 552
rect 181732 377 181760 1838
rect 181824 513 181852 2382
rect 182100 2038 182128 3606
rect 182088 2032 182140 2038
rect 182088 1974 182140 1980
rect 184584 1970 184612 4966
rect 186332 4826 186360 9318
rect 186320 4820 186372 4826
rect 186320 4762 186372 4768
rect 186424 3233 186452 9454
rect 186976 8498 187004 10231
rect 187712 9518 187740 10231
rect 188632 9586 188660 10231
rect 188620 9580 188672 9586
rect 188620 9522 188672 9528
rect 187700 9512 187752 9518
rect 187700 9454 187752 9460
rect 189460 9042 189488 10231
rect 189448 9036 189500 9042
rect 189448 8978 189500 8984
rect 189724 8968 189776 8974
rect 189724 8910 189776 8916
rect 186964 8492 187016 8498
rect 186964 8434 187016 8440
rect 189736 7750 189764 8910
rect 189920 8362 189948 10231
rect 190184 9580 190236 9586
rect 190184 9522 190236 9528
rect 190828 9580 190880 9586
rect 190828 9522 190880 9528
rect 189908 8356 189960 8362
rect 189908 8298 189960 8304
rect 189724 7744 189776 7750
rect 189724 7686 189776 7692
rect 190196 6934 190224 9522
rect 190840 9042 190868 9522
rect 190920 9376 190972 9382
rect 190920 9318 190972 9324
rect 190828 9036 190880 9042
rect 190828 8978 190880 8984
rect 190932 8974 190960 9318
rect 190644 8968 190696 8974
rect 190644 8910 190696 8916
rect 190920 8968 190972 8974
rect 190920 8910 190972 8916
rect 191012 8968 191064 8974
rect 191012 8910 191064 8916
rect 190368 8832 190420 8838
rect 190368 8774 190420 8780
rect 190380 8498 190408 8774
rect 190368 8492 190420 8498
rect 190368 8434 190420 8440
rect 190184 6928 190236 6934
rect 190184 6870 190236 6876
rect 188804 6792 188856 6798
rect 189724 6792 189776 6798
rect 188804 6734 188856 6740
rect 189446 6760 189502 6769
rect 188816 6458 188844 6734
rect 189356 6724 189408 6730
rect 189724 6734 189776 6740
rect 189446 6695 189502 6704
rect 189356 6666 189408 6672
rect 189368 6458 189396 6666
rect 189460 6458 189488 6695
rect 189736 6458 189764 6734
rect 189816 6724 189868 6730
rect 189816 6666 189868 6672
rect 189828 6458 189856 6666
rect 188804 6452 188856 6458
rect 188804 6394 188856 6400
rect 189356 6452 189408 6458
rect 189356 6394 189408 6400
rect 189448 6452 189500 6458
rect 189448 6394 189500 6400
rect 189724 6452 189776 6458
rect 189724 6394 189776 6400
rect 189816 6452 189868 6458
rect 189816 6394 189868 6400
rect 188816 5846 188844 6394
rect 188804 5840 188856 5846
rect 188804 5782 188856 5788
rect 188816 5710 188844 5782
rect 188804 5704 188856 5710
rect 188804 5646 188856 5652
rect 189368 5574 189396 6394
rect 190000 6384 190052 6390
rect 190000 6326 190052 6332
rect 189540 6316 189592 6322
rect 189540 6258 189592 6264
rect 189552 5642 189580 6258
rect 190012 6225 190040 6326
rect 189998 6216 190054 6225
rect 189998 6151 190054 6160
rect 190460 5840 190512 5846
rect 190460 5782 190512 5788
rect 189540 5636 189592 5642
rect 189540 5578 189592 5584
rect 189356 5568 189408 5574
rect 189356 5510 189408 5516
rect 187608 4480 187660 4486
rect 187608 4422 187660 4428
rect 187148 3460 187200 3466
rect 187148 3402 187200 3408
rect 186410 3224 186466 3233
rect 186410 3159 186466 3168
rect 184756 2440 184808 2446
rect 184756 2382 184808 2388
rect 186964 2440 187016 2446
rect 186964 2382 187016 2388
rect 184572 1964 184624 1970
rect 184572 1906 184624 1912
rect 183008 1896 183060 1902
rect 183008 1838 183060 1844
rect 184296 1896 184348 1902
rect 184296 1838 184348 1844
rect 181996 1352 182048 1358
rect 181996 1294 182048 1300
rect 181810 504 181866 513
rect 181810 439 181866 448
rect 176842 368 176898 377
rect 176842 303 176898 312
rect 181718 368 181774 377
rect 181718 303 181774 312
rect 160558 232 160614 241
rect 160558 167 160614 176
rect 174266 232 174322 241
rect 174266 167 174322 176
rect 160006 96 160062 105
rect 141238 31 141294 40
rect 149336 60 149388 66
rect 182008 66 182036 1294
rect 183020 513 183048 1838
rect 183284 1352 183336 1358
rect 183284 1294 183336 1300
rect 183296 513 183324 1294
rect 184308 513 184336 1838
rect 184572 1352 184624 1358
rect 184572 1294 184624 1300
rect 183006 504 183062 513
rect 183006 439 183062 448
rect 183282 504 183338 513
rect 183282 439 183338 448
rect 184294 504 184350 513
rect 184294 439 184350 448
rect 184584 338 184612 1294
rect 184768 513 184796 2382
rect 186320 1896 186372 1902
rect 186320 1838 186372 1844
rect 186332 1465 186360 1838
rect 186318 1456 186374 1465
rect 186318 1391 186374 1400
rect 185492 1352 185544 1358
rect 185492 1294 185544 1300
rect 185504 513 185532 1294
rect 186976 513 187004 2382
rect 187160 1970 187188 3402
rect 187148 1964 187200 1970
rect 187148 1906 187200 1912
rect 187148 1352 187200 1358
rect 187148 1294 187200 1300
rect 187160 542 187188 1294
rect 187620 1222 187648 4422
rect 190472 4146 190500 5782
rect 190460 4140 190512 4146
rect 190460 4082 190512 4088
rect 189724 3596 189776 3602
rect 189724 3538 189776 3544
rect 188160 1896 188212 1902
rect 188160 1838 188212 1844
rect 187608 1216 187660 1222
rect 187608 1158 187660 1164
rect 187148 536 187200 542
rect 184754 504 184810 513
rect 184754 439 184810 448
rect 185490 504 185546 513
rect 185490 439 185546 448
rect 186962 504 187018 513
rect 188172 513 188200 1838
rect 189736 1358 189764 3538
rect 190366 2816 190422 2825
rect 190422 2774 190500 2802
rect 190366 2751 190422 2760
rect 190472 2650 190500 2774
rect 190460 2644 190512 2650
rect 190460 2586 190512 2592
rect 190656 2038 190684 8910
rect 191024 2446 191052 8910
rect 191300 8362 191328 10367
rect 191378 10296 191434 10305
rect 191378 10231 191434 10240
rect 191392 9450 191420 10231
rect 192024 9580 192076 9586
rect 192024 9522 192076 9528
rect 192668 9580 192720 9586
rect 192668 9522 192720 9528
rect 191380 9444 191432 9450
rect 191380 9386 191432 9392
rect 192036 9178 192064 9522
rect 192024 9172 192076 9178
rect 192024 9114 192076 9120
rect 192116 8968 192168 8974
rect 192116 8910 192168 8916
rect 191932 8832 191984 8838
rect 191932 8774 191984 8780
rect 191944 8498 191972 8774
rect 191932 8492 191984 8498
rect 191932 8434 191984 8440
rect 191288 8356 191340 8362
rect 191288 8298 191340 8304
rect 191196 3936 191248 3942
rect 191196 3878 191248 3884
rect 191104 2848 191156 2854
rect 191104 2790 191156 2796
rect 190920 2440 190972 2446
rect 190920 2382 190972 2388
rect 191012 2440 191064 2446
rect 191012 2382 191064 2388
rect 190932 2106 190960 2382
rect 191012 2304 191064 2310
rect 191012 2246 191064 2252
rect 190920 2100 190972 2106
rect 190920 2042 190972 2048
rect 190644 2032 190696 2038
rect 190644 1974 190696 1980
rect 191024 1970 191052 2246
rect 191012 1964 191064 1970
rect 191012 1906 191064 1912
rect 191024 1358 191052 1906
rect 188620 1352 188672 1358
rect 188620 1294 188672 1300
rect 189448 1352 189500 1358
rect 189448 1294 189500 1300
rect 189724 1352 189776 1358
rect 189724 1294 189776 1300
rect 191012 1352 191064 1358
rect 191012 1294 191064 1300
rect 188632 513 188660 1294
rect 189460 513 189488 1294
rect 191116 513 191144 2790
rect 191208 2378 191236 3878
rect 191288 3052 191340 3058
rect 191288 2994 191340 3000
rect 191196 2372 191248 2378
rect 191196 2314 191248 2320
rect 191208 1834 191236 2314
rect 191196 1828 191248 1834
rect 191196 1770 191248 1776
rect 191300 1358 191328 2994
rect 191746 2816 191802 2825
rect 191802 2774 191880 2802
rect 191746 2751 191802 2760
rect 191852 2650 191880 2774
rect 191840 2644 191892 2650
rect 191840 2586 191892 2592
rect 191380 2372 191432 2378
rect 191380 2314 191432 2320
rect 191392 1426 191420 2314
rect 192128 2009 192156 8910
rect 192484 8900 192536 8906
rect 192484 8842 192536 8848
rect 192496 8498 192524 8842
rect 192680 8498 192708 9522
rect 192392 8492 192444 8498
rect 192392 8434 192444 8440
rect 192484 8492 192536 8498
rect 192484 8434 192536 8440
rect 192668 8492 192720 8498
rect 192668 8434 192720 8440
rect 192404 2582 192432 8434
rect 192864 8362 192892 10367
rect 192942 10296 192998 10305
rect 192942 10231 192998 10240
rect 192956 9450 192984 10231
rect 192944 9444 192996 9450
rect 192944 9386 192996 9392
rect 193324 8974 193352 10474
rect 196164 10328 196216 10334
rect 194046 10296 194102 10305
rect 194046 10231 194102 10240
rect 194322 10296 194378 10305
rect 194322 10231 194378 10240
rect 195518 10296 195574 10305
rect 195518 10231 195574 10240
rect 195794 10296 195850 10305
rect 196164 10270 196216 10276
rect 196530 10296 196586 10305
rect 195794 10231 195850 10240
rect 193312 8968 193364 8974
rect 193312 8910 193364 8916
rect 193128 8832 193180 8838
rect 193128 8774 193180 8780
rect 193140 8498 193168 8774
rect 193128 8492 193180 8498
rect 193128 8434 193180 8440
rect 192852 8356 192904 8362
rect 192852 8298 192904 8304
rect 193324 6914 193352 8910
rect 193864 8832 193916 8838
rect 193864 8774 193916 8780
rect 193876 8498 193904 8774
rect 193864 8492 193916 8498
rect 193864 8434 193916 8440
rect 194060 8362 194088 10231
rect 194336 9450 194364 10231
rect 194600 9580 194652 9586
rect 194600 9522 194652 9528
rect 194324 9444 194376 9450
rect 194324 9386 194376 9392
rect 194508 9376 194560 9382
rect 194508 9318 194560 9324
rect 194520 9110 194548 9318
rect 194612 9178 194640 9522
rect 195532 9450 195560 10231
rect 195612 9580 195664 9586
rect 195612 9522 195664 9528
rect 195520 9444 195572 9450
rect 195520 9386 195572 9392
rect 194600 9172 194652 9178
rect 194600 9114 194652 9120
rect 194508 9104 194560 9110
rect 194508 9046 194560 9052
rect 194692 9104 194744 9110
rect 194692 9046 194744 9052
rect 195336 9104 195388 9110
rect 195336 9046 195388 9052
rect 195520 9104 195572 9110
rect 195520 9046 195572 9052
rect 194704 8974 194732 9046
rect 194692 8968 194744 8974
rect 194692 8910 194744 8916
rect 194048 8356 194100 8362
rect 194048 8298 194100 8304
rect 194704 6914 194732 8910
rect 195348 8838 195376 9046
rect 195532 8974 195560 9046
rect 195520 8968 195572 8974
rect 195520 8910 195572 8916
rect 195336 8832 195388 8838
rect 195336 8774 195388 8780
rect 195348 8265 195376 8774
rect 195334 8256 195390 8265
rect 195334 8191 195390 8200
rect 195532 6914 195560 8910
rect 195624 8498 195652 9522
rect 195612 8492 195664 8498
rect 195612 8434 195664 8440
rect 195808 8362 195836 10231
rect 195980 8900 196032 8906
rect 195980 8842 196032 8848
rect 195992 8430 196020 8842
rect 196072 8832 196124 8838
rect 196072 8774 196124 8780
rect 196084 8498 196112 8774
rect 196072 8492 196124 8498
rect 196072 8434 196124 8440
rect 195980 8424 196032 8430
rect 195980 8366 196032 8372
rect 195796 8356 195848 8362
rect 195796 8298 195848 8304
rect 196176 8294 196204 10270
rect 196530 10231 196586 10240
rect 197266 10296 197322 10305
rect 197266 10231 197322 10240
rect 198002 10296 198058 10305
rect 198002 10231 198058 10240
rect 199106 10296 199162 10305
rect 199106 10231 199162 10240
rect 199934 10296 199990 10305
rect 199934 10231 199990 10240
rect 196348 9920 196400 9926
rect 196348 9862 196400 9868
rect 196360 8974 196388 9862
rect 196544 9450 196572 10231
rect 197084 10192 197136 10198
rect 197084 10134 197136 10140
rect 196532 9444 196584 9450
rect 196532 9386 196584 9392
rect 196348 8968 196400 8974
rect 196348 8910 196400 8916
rect 195980 8288 196032 8294
rect 195980 8230 196032 8236
rect 196164 8288 196216 8294
rect 196164 8230 196216 8236
rect 193324 6886 193536 6914
rect 194704 6886 194824 6914
rect 192392 2576 192444 2582
rect 192392 2518 192444 2524
rect 192852 2576 192904 2582
rect 192852 2518 192904 2524
rect 192208 2440 192260 2446
rect 192208 2382 192260 2388
rect 192220 2106 192248 2382
rect 192208 2100 192260 2106
rect 192208 2042 192260 2048
rect 191838 2000 191894 2009
rect 191838 1935 191894 1944
rect 192114 2000 192170 2009
rect 192114 1935 192170 1944
rect 191852 1902 191880 1935
rect 192864 1902 192892 2518
rect 193508 1970 193536 6886
rect 194600 2304 194652 2310
rect 194600 2246 194652 2252
rect 193496 1964 193548 1970
rect 193496 1906 193548 1912
rect 191840 1896 191892 1902
rect 191840 1838 191892 1844
rect 192852 1896 192904 1902
rect 194612 1873 194640 2246
rect 194796 1902 194824 6886
rect 195348 6886 195560 6914
rect 195348 1970 195376 6886
rect 195704 2440 195756 2446
rect 195704 2382 195756 2388
rect 195716 1970 195744 2382
rect 195992 1970 196020 8230
rect 196360 2774 196388 8910
rect 197096 8430 197124 10134
rect 197280 9450 197308 10231
rect 197544 9580 197596 9586
rect 197544 9522 197596 9528
rect 197728 9580 197780 9586
rect 197728 9522 197780 9528
rect 197268 9444 197320 9450
rect 197268 9386 197320 9392
rect 197176 9376 197228 9382
rect 197176 9318 197228 9324
rect 197084 8424 197136 8430
rect 197084 8366 197136 8372
rect 196268 2746 196388 2774
rect 197096 2774 197124 8366
rect 197188 8090 197216 9318
rect 197556 8498 197584 9522
rect 197740 9042 197768 9522
rect 197912 9512 197964 9518
rect 197912 9454 197964 9460
rect 197728 9036 197780 9042
rect 197728 8978 197780 8984
rect 197740 8498 197768 8978
rect 197544 8492 197596 8498
rect 197544 8434 197596 8440
rect 197728 8492 197780 8498
rect 197728 8434 197780 8440
rect 197176 8084 197228 8090
rect 197176 8026 197228 8032
rect 197096 2746 197216 2774
rect 196164 2440 196216 2446
rect 196164 2382 196216 2388
rect 196072 2304 196124 2310
rect 196072 2246 196124 2252
rect 195336 1964 195388 1970
rect 195336 1906 195388 1912
rect 195704 1964 195756 1970
rect 195704 1906 195756 1912
rect 195980 1964 196032 1970
rect 195980 1906 196032 1912
rect 194784 1896 194836 1902
rect 192852 1838 192904 1844
rect 194598 1864 194654 1873
rect 196084 1873 196112 2246
rect 194784 1838 194836 1844
rect 196070 1864 196126 1873
rect 194598 1799 194654 1808
rect 196070 1799 196126 1808
rect 193220 1760 193272 1766
rect 193220 1702 193272 1708
rect 194048 1760 194100 1766
rect 194048 1702 194100 1708
rect 194600 1760 194652 1766
rect 194600 1702 194652 1708
rect 196072 1760 196124 1766
rect 196072 1702 196124 1708
rect 191380 1420 191432 1426
rect 191380 1362 191432 1368
rect 191288 1352 191340 1358
rect 191288 1294 191340 1300
rect 193232 1290 193260 1702
rect 194060 1358 194088 1702
rect 194612 1358 194640 1702
rect 196084 1358 196112 1702
rect 196176 1494 196204 2382
rect 196164 1488 196216 1494
rect 196164 1430 196216 1436
rect 196268 1426 196296 2746
rect 196624 2304 196676 2310
rect 196624 2246 196676 2252
rect 196440 2032 196492 2038
rect 196440 1974 196492 1980
rect 196256 1420 196308 1426
rect 196256 1362 196308 1368
rect 196452 1358 196480 1974
rect 194048 1352 194100 1358
rect 194048 1294 194100 1300
rect 194600 1352 194652 1358
rect 194600 1294 194652 1300
rect 196072 1352 196124 1358
rect 196072 1294 196124 1300
rect 196440 1352 196492 1358
rect 196440 1294 196492 1300
rect 193220 1284 193272 1290
rect 193220 1226 193272 1232
rect 192576 1216 192628 1222
rect 192576 1158 192628 1164
rect 192852 1216 192904 1222
rect 192852 1158 192904 1164
rect 193588 1216 193640 1222
rect 193588 1158 193640 1164
rect 195612 1216 195664 1222
rect 195612 1158 195664 1164
rect 187148 478 187200 484
rect 188158 504 188214 513
rect 186962 439 187018 448
rect 188158 439 188214 448
rect 188618 504 188674 513
rect 188618 439 188674 448
rect 189446 504 189502 513
rect 189446 439 189502 448
rect 191102 504 191158 513
rect 191102 439 191158 448
rect 192588 377 192616 1158
rect 192864 513 192892 1158
rect 193600 513 193628 1158
rect 195624 513 195652 1158
rect 196636 513 196664 2246
rect 197188 1970 197216 2746
rect 197544 2440 197596 2446
rect 197544 2382 197596 2388
rect 197360 2304 197412 2310
rect 197360 2246 197412 2252
rect 197176 1964 197228 1970
rect 197176 1906 197228 1912
rect 197372 1465 197400 2246
rect 197556 2106 197584 2382
rect 197544 2100 197596 2106
rect 197544 2042 197596 2048
rect 197358 1456 197414 1465
rect 197924 1426 197952 9454
rect 198016 9178 198044 10231
rect 198004 9172 198056 9178
rect 198004 9114 198056 9120
rect 198556 8968 198608 8974
rect 198556 8910 198608 8916
rect 198568 8498 198596 8910
rect 198556 8492 198608 8498
rect 198556 8434 198608 8440
rect 198740 8424 198792 8430
rect 198740 8366 198792 8372
rect 198752 8022 198780 8366
rect 199120 8362 199148 10231
rect 199752 9172 199804 9178
rect 199752 9114 199804 9120
rect 199764 8974 199792 9114
rect 199752 8968 199804 8974
rect 199752 8910 199804 8916
rect 199200 8832 199252 8838
rect 199200 8774 199252 8780
rect 199212 8498 199240 8774
rect 199200 8492 199252 8498
rect 199200 8434 199252 8440
rect 199948 8362 199976 10231
rect 200132 9178 200160 10542
rect 200762 10296 200818 10305
rect 200762 10231 200818 10240
rect 200946 10296 201002 10305
rect 200946 10231 201002 10240
rect 200120 9172 200172 9178
rect 200120 9114 200172 9120
rect 200672 9172 200724 9178
rect 200672 9114 200724 9120
rect 199108 8356 199160 8362
rect 199108 8298 199160 8304
rect 199936 8356 199988 8362
rect 199936 8298 199988 8304
rect 198740 8016 198792 8022
rect 198740 7958 198792 7964
rect 199384 8016 199436 8022
rect 199384 7958 199436 7964
rect 198646 2816 198702 2825
rect 198702 2774 198780 2802
rect 198646 2751 198702 2760
rect 198752 2650 198780 2774
rect 198740 2644 198792 2650
rect 198740 2586 198792 2592
rect 198280 2440 198332 2446
rect 198280 2382 198332 2388
rect 198292 1494 198320 2382
rect 199396 1970 199424 7958
rect 200132 7426 200160 9114
rect 200684 8974 200712 9114
rect 200672 8968 200724 8974
rect 200672 8910 200724 8916
rect 200212 8832 200264 8838
rect 200212 8774 200264 8780
rect 200224 8498 200252 8774
rect 200212 8492 200264 8498
rect 200212 8434 200264 8440
rect 200132 7398 200344 7426
rect 200026 2816 200082 2825
rect 200082 2760 200252 2774
rect 200026 2751 200252 2760
rect 200040 2746 200252 2751
rect 200224 2582 200252 2746
rect 200212 2576 200264 2582
rect 200212 2518 200264 2524
rect 199752 2440 199804 2446
rect 199752 2382 199804 2388
rect 200212 2440 200264 2446
rect 200212 2382 200264 2388
rect 199764 2106 199792 2382
rect 199752 2100 199804 2106
rect 199752 2042 199804 2048
rect 200224 2038 200252 2382
rect 200212 2032 200264 2038
rect 200212 1974 200264 1980
rect 200316 1970 200344 7398
rect 200684 1970 200712 8910
rect 200776 8362 200804 10231
rect 200960 8362 200988 10231
rect 201316 9104 201368 9110
rect 201316 9046 201368 9052
rect 201328 8974 201356 9046
rect 202340 8974 202368 10610
rect 208306 10568 208362 10577
rect 208306 10503 208362 10512
rect 213458 10568 213514 10577
rect 213458 10503 213514 10512
rect 202418 10432 202474 10441
rect 202418 10367 202474 10376
rect 202432 9382 202460 10367
rect 202510 10296 202566 10305
rect 204074 10296 204130 10305
rect 202510 10231 202566 10240
rect 203064 10260 203116 10266
rect 202524 9450 202552 10231
rect 204074 10231 204130 10240
rect 205822 10296 205878 10305
rect 205822 10231 205878 10240
rect 203064 10202 203116 10208
rect 202696 9580 202748 9586
rect 202696 9522 202748 9528
rect 202512 9444 202564 9450
rect 202512 9386 202564 9392
rect 202420 9376 202472 9382
rect 202420 9318 202472 9324
rect 201316 8968 201368 8974
rect 201316 8910 201368 8916
rect 202328 8968 202380 8974
rect 202328 8910 202380 8916
rect 201040 8832 201092 8838
rect 201040 8774 201092 8780
rect 201052 8498 201080 8774
rect 201040 8492 201092 8498
rect 201040 8434 201092 8440
rect 200764 8356 200816 8362
rect 200764 8298 200816 8304
rect 200948 8356 201000 8362
rect 200948 8298 201000 8304
rect 200764 6112 200816 6118
rect 200764 6054 200816 6060
rect 200776 5574 200804 6054
rect 200764 5568 200816 5574
rect 200764 5510 200816 5516
rect 201040 2440 201092 2446
rect 201040 2382 201092 2388
rect 199384 1964 199436 1970
rect 199384 1906 199436 1912
rect 200304 1964 200356 1970
rect 200304 1906 200356 1912
rect 200672 1964 200724 1970
rect 200672 1906 200724 1912
rect 198372 1896 198424 1902
rect 198372 1838 198424 1844
rect 198280 1488 198332 1494
rect 198280 1430 198332 1436
rect 197358 1391 197414 1400
rect 197912 1420 197964 1426
rect 197912 1362 197964 1368
rect 198384 1358 198412 1838
rect 200580 1760 200632 1766
rect 200580 1702 200632 1708
rect 200592 1358 200620 1702
rect 198372 1352 198424 1358
rect 198372 1294 198424 1300
rect 200580 1352 200632 1358
rect 200580 1294 200632 1300
rect 201052 1290 201080 2382
rect 201224 2304 201276 2310
rect 201224 2246 201276 2252
rect 201040 1284 201092 1290
rect 201040 1226 201092 1232
rect 199936 1216 199988 1222
rect 199936 1158 199988 1164
rect 199948 513 199976 1158
rect 201236 513 201264 2246
rect 201328 1426 201356 8910
rect 201868 8832 201920 8838
rect 201868 8774 201920 8780
rect 201880 8498 201908 8774
rect 201868 8492 201920 8498
rect 201868 8434 201920 8440
rect 201406 2816 201462 2825
rect 201462 2774 201540 2802
rect 201406 2751 201462 2760
rect 201512 2582 201540 2774
rect 201500 2576 201552 2582
rect 201500 2518 201552 2524
rect 202340 1970 202368 8910
rect 202512 8900 202564 8906
rect 202512 8842 202564 8848
rect 202524 8498 202552 8842
rect 202708 8498 202736 9522
rect 203076 8974 203104 10202
rect 203740 9820 204048 9829
rect 203740 9818 203746 9820
rect 203802 9818 203826 9820
rect 203882 9818 203906 9820
rect 203962 9818 203986 9820
rect 204042 9818 204048 9820
rect 203802 9766 203804 9818
rect 203984 9766 203986 9818
rect 203740 9764 203746 9766
rect 203802 9764 203826 9766
rect 203882 9764 203906 9766
rect 203962 9764 203986 9766
rect 204042 9764 204048 9766
rect 203740 9755 204048 9764
rect 203432 9580 203484 9586
rect 203432 9522 203484 9528
rect 203444 9178 203472 9522
rect 204088 9178 204116 10231
rect 204352 10192 204404 10198
rect 204352 10134 204404 10140
rect 204364 9926 204392 10134
rect 204260 9920 204312 9926
rect 204260 9862 204312 9868
rect 204352 9920 204404 9926
rect 204352 9862 204404 9868
rect 203340 9172 203392 9178
rect 203340 9114 203392 9120
rect 203432 9172 203484 9178
rect 203432 9114 203484 9120
rect 204076 9172 204128 9178
rect 204076 9114 204128 9120
rect 203064 8968 203116 8974
rect 203064 8910 203116 8916
rect 202512 8492 202564 8498
rect 202512 8434 202564 8440
rect 202696 8492 202748 8498
rect 202696 8434 202748 8440
rect 202972 8424 203024 8430
rect 202972 8366 203024 8372
rect 202984 7886 203012 8366
rect 202972 7880 203024 7886
rect 202972 7822 203024 7828
rect 202788 2508 202840 2514
rect 202788 2450 202840 2456
rect 202696 2440 202748 2446
rect 202696 2382 202748 2388
rect 202708 2038 202736 2382
rect 202696 2032 202748 2038
rect 202696 1974 202748 1980
rect 202328 1964 202380 1970
rect 202328 1906 202380 1912
rect 202800 1902 202828 2450
rect 201500 1896 201552 1902
rect 201500 1838 201552 1844
rect 202788 1896 202840 1902
rect 202788 1838 202840 1844
rect 201316 1420 201368 1426
rect 201316 1362 201368 1368
rect 201512 1358 201540 1838
rect 202880 1760 202932 1766
rect 202880 1702 202932 1708
rect 202892 1465 202920 1702
rect 203076 1494 203104 8910
rect 203352 8906 203380 9114
rect 204272 9110 204300 9862
rect 205836 9586 205864 10231
rect 206558 10160 206614 10169
rect 206558 10095 206614 10104
rect 207662 10160 207718 10169
rect 207662 10095 207718 10104
rect 206572 9586 206600 10095
rect 207676 9586 207704 10095
rect 208320 9586 208348 10503
rect 210882 10432 210938 10441
rect 210882 10367 210938 10376
rect 208950 10160 209006 10169
rect 208950 10095 209006 10104
rect 209318 10160 209374 10169
rect 209318 10095 209374 10104
rect 208964 9586 208992 10095
rect 209332 9586 209360 10095
rect 210896 9586 210924 10367
rect 211252 10192 211304 10198
rect 211158 10160 211214 10169
rect 211252 10134 211304 10140
rect 212538 10160 212594 10169
rect 211158 10095 211214 10104
rect 211172 9586 211200 10095
rect 205824 9580 205876 9586
rect 205824 9522 205876 9528
rect 206560 9580 206612 9586
rect 206560 9522 206612 9528
rect 207664 9580 207716 9586
rect 207664 9522 207716 9528
rect 208308 9580 208360 9586
rect 208308 9522 208360 9528
rect 208952 9580 209004 9586
rect 208952 9522 209004 9528
rect 209320 9580 209372 9586
rect 209320 9522 209372 9528
rect 210884 9580 210936 9586
rect 210884 9522 210936 9528
rect 211160 9580 211212 9586
rect 211160 9522 211212 9528
rect 207020 9444 207072 9450
rect 207020 9386 207072 9392
rect 206836 9376 206888 9382
rect 206836 9318 206888 9324
rect 204260 9104 204312 9110
rect 204260 9046 204312 9052
rect 203524 8968 203576 8974
rect 203524 8910 203576 8916
rect 203340 8900 203392 8906
rect 203340 8842 203392 8848
rect 203536 8498 203564 8910
rect 203740 8732 204048 8741
rect 203740 8730 203746 8732
rect 203802 8730 203826 8732
rect 203882 8730 203906 8732
rect 203962 8730 203986 8732
rect 204042 8730 204048 8732
rect 203802 8678 203804 8730
rect 203984 8678 203986 8730
rect 203740 8676 203746 8678
rect 203802 8676 203826 8678
rect 203882 8676 203906 8678
rect 203962 8676 203986 8678
rect 204042 8676 204048 8678
rect 203740 8667 204048 8676
rect 203524 8492 203576 8498
rect 203524 8434 203576 8440
rect 203248 8356 203300 8362
rect 203248 8298 203300 8304
rect 203156 2984 203208 2990
rect 203156 2926 203208 2932
rect 203168 2446 203196 2926
rect 203156 2440 203208 2446
rect 203156 2382 203208 2388
rect 203260 1970 203288 8298
rect 203740 7644 204048 7653
rect 203740 7642 203746 7644
rect 203802 7642 203826 7644
rect 203882 7642 203906 7644
rect 203962 7642 203986 7644
rect 204042 7642 204048 7644
rect 203802 7590 203804 7642
rect 203984 7590 203986 7642
rect 203740 7588 203746 7590
rect 203802 7588 203826 7590
rect 203882 7588 203906 7590
rect 203962 7588 203986 7590
rect 204042 7588 204048 7590
rect 203740 7579 204048 7588
rect 203740 6556 204048 6565
rect 203740 6554 203746 6556
rect 203802 6554 203826 6556
rect 203882 6554 203906 6556
rect 203962 6554 203986 6556
rect 204042 6554 204048 6556
rect 203802 6502 203804 6554
rect 203984 6502 203986 6554
rect 203740 6500 203746 6502
rect 203802 6500 203826 6502
rect 203882 6500 203906 6502
rect 203962 6500 203986 6502
rect 204042 6500 204048 6502
rect 203740 6491 204048 6500
rect 206744 5636 206796 5642
rect 206744 5578 206796 5584
rect 206190 5536 206246 5545
rect 203740 5468 204048 5477
rect 206190 5471 206246 5480
rect 203740 5466 203746 5468
rect 203802 5466 203826 5468
rect 203882 5466 203906 5468
rect 203962 5466 203986 5468
rect 204042 5466 204048 5468
rect 203802 5414 203804 5466
rect 203984 5414 203986 5466
rect 203740 5412 203746 5414
rect 203802 5412 203826 5414
rect 203882 5412 203906 5414
rect 203962 5412 203986 5414
rect 204042 5412 204048 5414
rect 203740 5403 204048 5412
rect 205640 5228 205692 5234
rect 205640 5170 205692 5176
rect 205652 4758 205680 5170
rect 205824 5160 205876 5166
rect 205824 5102 205876 5108
rect 205640 4752 205692 4758
rect 205640 4694 205692 4700
rect 205652 4622 205680 4694
rect 205836 4622 205864 5102
rect 205640 4616 205692 4622
rect 205640 4558 205692 4564
rect 205824 4616 205876 4622
rect 205824 4558 205876 4564
rect 203740 4380 204048 4389
rect 203740 4378 203746 4380
rect 203802 4378 203826 4380
rect 203882 4378 203906 4380
rect 203962 4378 203986 4380
rect 204042 4378 204048 4380
rect 203802 4326 203804 4378
rect 203984 4326 203986 4378
rect 203740 4324 203746 4326
rect 203802 4324 203826 4326
rect 203882 4324 203906 4326
rect 203962 4324 203986 4326
rect 204042 4324 204048 4326
rect 203740 4315 204048 4324
rect 205652 4214 205680 4558
rect 205640 4208 205692 4214
rect 205640 4150 205692 4156
rect 203740 3292 204048 3301
rect 203740 3290 203746 3292
rect 203802 3290 203826 3292
rect 203882 3290 203906 3292
rect 203962 3290 203986 3292
rect 204042 3290 204048 3292
rect 203802 3238 203804 3290
rect 203984 3238 203986 3290
rect 203740 3236 203746 3238
rect 203802 3236 203826 3238
rect 203882 3236 203906 3238
rect 203962 3236 203986 3238
rect 204042 3236 204048 3238
rect 203740 3227 204048 3236
rect 206204 2922 206232 5471
rect 206756 5370 206784 5578
rect 206744 5364 206796 5370
rect 206744 5306 206796 5312
rect 206848 5234 206876 9318
rect 206652 5228 206704 5234
rect 206652 5170 206704 5176
rect 206836 5228 206888 5234
rect 206836 5170 206888 5176
rect 206468 5024 206520 5030
rect 206468 4966 206520 4972
rect 206480 4690 206508 4966
rect 206664 4758 206692 5170
rect 206652 4752 206704 4758
rect 206652 4694 206704 4700
rect 206468 4684 206520 4690
rect 206468 4626 206520 4632
rect 206560 4140 206612 4146
rect 206560 4082 206612 4088
rect 206652 4140 206704 4146
rect 206652 4082 206704 4088
rect 206744 4140 206796 4146
rect 206744 4082 206796 4088
rect 206572 3058 206600 4082
rect 206664 3126 206692 4082
rect 206756 3398 206784 4082
rect 207032 3602 207060 9386
rect 207480 9376 207532 9382
rect 207480 9318 207532 9324
rect 208768 9376 208820 9382
rect 208768 9318 208820 9324
rect 210056 9376 210108 9382
rect 210056 9318 210108 9324
rect 210700 9376 210752 9382
rect 210700 9318 210752 9324
rect 207110 7712 207166 7721
rect 207110 7647 207166 7656
rect 207124 5642 207152 7647
rect 207492 6322 207520 9318
rect 207480 6316 207532 6322
rect 207480 6258 207532 6264
rect 208492 6248 208544 6254
rect 208492 6190 208544 6196
rect 207756 6180 207808 6186
rect 207756 6122 207808 6128
rect 207296 6112 207348 6118
rect 207296 6054 207348 6060
rect 207308 5710 207336 6054
rect 207296 5704 207348 5710
rect 207296 5646 207348 5652
rect 207112 5636 207164 5642
rect 207112 5578 207164 5584
rect 207480 5636 207532 5642
rect 207480 5578 207532 5584
rect 207492 5370 207520 5578
rect 207480 5364 207532 5370
rect 207480 5306 207532 5312
rect 207112 5160 207164 5166
rect 207112 5102 207164 5108
rect 207020 3596 207072 3602
rect 207020 3538 207072 3544
rect 206744 3392 206796 3398
rect 206744 3334 206796 3340
rect 206652 3120 206704 3126
rect 206652 3062 206704 3068
rect 206560 3052 206612 3058
rect 206560 2994 206612 3000
rect 206192 2916 206244 2922
rect 206192 2858 206244 2864
rect 204076 2304 204128 2310
rect 204076 2246 204128 2252
rect 203740 2204 204048 2213
rect 203740 2202 203746 2204
rect 203802 2202 203826 2204
rect 203882 2202 203906 2204
rect 203962 2202 203986 2204
rect 204042 2202 204048 2204
rect 203802 2150 203804 2202
rect 203984 2150 203986 2202
rect 203740 2148 203746 2150
rect 203802 2148 203826 2150
rect 203882 2148 203906 2150
rect 203962 2148 203986 2150
rect 204042 2148 204048 2150
rect 203740 2139 204048 2148
rect 203248 1964 203300 1970
rect 203248 1906 203300 1912
rect 203064 1488 203116 1494
rect 202878 1456 202934 1465
rect 203064 1430 203116 1436
rect 202878 1391 202934 1400
rect 201500 1352 201552 1358
rect 201500 1294 201552 1300
rect 202420 1216 202472 1222
rect 202420 1158 202472 1164
rect 202432 513 202460 1158
rect 203740 1116 204048 1125
rect 203740 1114 203746 1116
rect 203802 1114 203826 1116
rect 203882 1114 203906 1116
rect 203962 1114 203986 1116
rect 204042 1114 204048 1116
rect 203802 1062 203804 1114
rect 203984 1062 203986 1114
rect 203740 1060 203746 1062
rect 203802 1060 203826 1062
rect 203882 1060 203906 1062
rect 203962 1060 203986 1062
rect 204042 1060 204048 1062
rect 203740 1051 204048 1060
rect 204088 513 204116 2246
rect 205824 1420 205876 1426
rect 205824 1362 205876 1368
rect 205836 921 205864 1362
rect 206560 1352 206612 1358
rect 206560 1294 206612 1300
rect 206572 921 206600 1294
rect 207124 1222 207152 5102
rect 207768 5098 207796 6122
rect 208400 5160 208452 5166
rect 208398 5128 208400 5137
rect 208452 5128 208454 5137
rect 207572 5092 207624 5098
rect 207756 5092 207808 5098
rect 207572 5034 207624 5040
rect 207676 5052 207756 5080
rect 207584 4554 207612 5034
rect 207572 4548 207624 4554
rect 207572 4490 207624 4496
rect 207480 4072 207532 4078
rect 207480 4014 207532 4020
rect 207492 3738 207520 4014
rect 207480 3732 207532 3738
rect 207480 3674 207532 3680
rect 207676 3602 207704 5052
rect 208398 5063 208454 5072
rect 207756 5034 207808 5040
rect 207940 4616 207992 4622
rect 207940 4558 207992 4564
rect 207572 3596 207624 3602
rect 207572 3538 207624 3544
rect 207664 3596 207716 3602
rect 207664 3538 207716 3544
rect 207584 1222 207612 3538
rect 207676 2854 207704 3538
rect 207952 3534 207980 4558
rect 208308 4004 208360 4010
rect 208308 3946 208360 3952
rect 207940 3528 207992 3534
rect 207940 3470 207992 3476
rect 208216 3528 208268 3534
rect 208320 3516 208348 3946
rect 208268 3488 208348 3516
rect 208216 3470 208268 3476
rect 207940 3392 207992 3398
rect 207940 3334 207992 3340
rect 207952 3058 207980 3334
rect 207940 3052 207992 3058
rect 207940 2994 207992 3000
rect 208308 2916 208360 2922
rect 208308 2858 208360 2864
rect 207664 2848 207716 2854
rect 207664 2790 207716 2796
rect 208124 2304 208176 2310
rect 208124 2246 208176 2252
rect 207664 1352 207716 1358
rect 207664 1294 207716 1300
rect 207112 1216 207164 1222
rect 207112 1158 207164 1164
rect 207572 1216 207624 1222
rect 207572 1158 207624 1164
rect 207676 921 207704 1294
rect 205822 912 205878 921
rect 205822 847 205878 856
rect 206558 912 206614 921
rect 206558 847 206614 856
rect 207662 912 207718 921
rect 207662 847 207718 856
rect 208136 610 208164 2246
rect 208320 1902 208348 2858
rect 208504 2088 208532 6190
rect 208584 5160 208636 5166
rect 208584 5102 208636 5108
rect 208596 4826 208624 5102
rect 208584 4820 208636 4826
rect 208584 4762 208636 4768
rect 208676 4616 208728 4622
rect 208676 4558 208728 4564
rect 208584 4548 208636 4554
rect 208584 4490 208636 4496
rect 208596 2292 208624 4490
rect 208688 3670 208716 4558
rect 208676 3664 208728 3670
rect 208676 3606 208728 3612
rect 208688 2990 208716 3606
rect 208780 3058 208808 9318
rect 209318 6624 209374 6633
rect 209318 6559 209374 6568
rect 209134 6488 209190 6497
rect 209134 6423 209190 6432
rect 209148 6322 209176 6423
rect 209332 6322 209360 6559
rect 209136 6316 209188 6322
rect 209136 6258 209188 6264
rect 209320 6316 209372 6322
rect 209320 6258 209372 6264
rect 209412 6248 209464 6254
rect 209240 6196 209412 6202
rect 209240 6190 209464 6196
rect 209240 6174 209452 6190
rect 209136 5636 209188 5642
rect 209136 5578 209188 5584
rect 209148 5545 209176 5578
rect 209134 5536 209190 5545
rect 209134 5471 209190 5480
rect 209240 5166 209268 6174
rect 209228 5160 209280 5166
rect 209228 5102 209280 5108
rect 209044 4616 209096 4622
rect 209044 4558 209096 4564
rect 208860 4480 208912 4486
rect 208860 4422 208912 4428
rect 208872 3126 208900 4422
rect 209056 3398 209084 4558
rect 209240 4010 209268 5102
rect 209964 5024 210016 5030
rect 209964 4966 210016 4972
rect 209976 4622 210004 4966
rect 209964 4616 210016 4622
rect 209964 4558 210016 4564
rect 209964 4480 210016 4486
rect 209964 4422 210016 4428
rect 209320 4276 209372 4282
rect 209320 4218 209372 4224
rect 209332 4078 209360 4218
rect 209976 4078 210004 4422
rect 209320 4072 209372 4078
rect 209320 4014 209372 4020
rect 209780 4072 209832 4078
rect 209780 4014 209832 4020
rect 209964 4072 210016 4078
rect 209964 4014 210016 4020
rect 209228 4004 209280 4010
rect 209228 3946 209280 3952
rect 209240 3466 209268 3946
rect 209332 3913 209360 4014
rect 209688 3936 209740 3942
rect 209318 3904 209374 3913
rect 209688 3878 209740 3884
rect 209318 3839 209374 3848
rect 209228 3460 209280 3466
rect 209228 3402 209280 3408
rect 209044 3392 209096 3398
rect 209044 3334 209096 3340
rect 208860 3120 208912 3126
rect 208860 3062 208912 3068
rect 208768 3052 208820 3058
rect 208768 2994 208820 3000
rect 208676 2984 208728 2990
rect 208676 2926 208728 2932
rect 208688 2446 208716 2926
rect 208872 2774 208900 3062
rect 208872 2746 208992 2774
rect 208964 2446 208992 2746
rect 209056 2446 209084 3334
rect 209700 3194 209728 3878
rect 209792 3194 209820 4014
rect 209872 3596 209924 3602
rect 209872 3538 209924 3544
rect 209688 3188 209740 3194
rect 209688 3130 209740 3136
rect 209780 3188 209832 3194
rect 209780 3130 209832 3136
rect 209136 2984 209188 2990
rect 209136 2926 209188 2932
rect 208676 2440 208728 2446
rect 208676 2382 208728 2388
rect 208952 2440 209004 2446
rect 208952 2382 209004 2388
rect 209044 2440 209096 2446
rect 209044 2382 209096 2388
rect 208596 2264 208716 2292
rect 208412 2060 208532 2088
rect 208308 1896 208360 1902
rect 208308 1838 208360 1844
rect 208308 1352 208360 1358
rect 208308 1294 208360 1300
rect 208124 604 208176 610
rect 208124 546 208176 552
rect 192850 504 192906 513
rect 192850 439 192906 448
rect 193586 504 193642 513
rect 193586 439 193642 448
rect 195610 504 195666 513
rect 195610 439 195666 448
rect 196622 504 196678 513
rect 196622 439 196678 448
rect 199934 504 199990 513
rect 199934 439 199990 448
rect 201222 504 201278 513
rect 201222 439 201278 448
rect 202418 504 202474 513
rect 202418 439 202474 448
rect 204074 504 204130 513
rect 204074 439 204130 448
rect 208320 377 208348 1294
rect 208412 1290 208440 2060
rect 208492 1964 208544 1970
rect 208492 1906 208544 1912
rect 208400 1284 208452 1290
rect 208400 1226 208452 1232
rect 208504 513 208532 1906
rect 208582 1592 208638 1601
rect 208582 1527 208638 1536
rect 208596 746 208624 1527
rect 208584 740 208636 746
rect 208584 682 208636 688
rect 208490 504 208546 513
rect 208688 474 208716 2264
rect 208952 1964 209004 1970
rect 208952 1906 209004 1912
rect 208964 1442 208992 1906
rect 208964 1414 209084 1442
rect 208952 1352 209004 1358
rect 208952 1294 209004 1300
rect 208964 921 208992 1294
rect 209056 1290 209084 1414
rect 209044 1284 209096 1290
rect 209044 1226 209096 1232
rect 209148 1222 209176 2926
rect 209596 2916 209648 2922
rect 209596 2858 209648 2864
rect 209608 1494 209636 2858
rect 209686 2816 209742 2825
rect 209686 2751 209742 2760
rect 209700 2514 209728 2751
rect 209688 2508 209740 2514
rect 209688 2450 209740 2456
rect 209688 2032 209740 2038
rect 209688 1974 209740 1980
rect 209596 1488 209648 1494
rect 209700 1465 209728 1974
rect 209780 1896 209832 1902
rect 209780 1838 209832 1844
rect 209596 1430 209648 1436
rect 209686 1456 209742 1465
rect 209686 1391 209742 1400
rect 209136 1216 209188 1222
rect 209136 1158 209188 1164
rect 209504 1216 209556 1222
rect 209504 1158 209556 1164
rect 208950 912 209006 921
rect 208950 847 209006 856
rect 208490 439 208546 448
rect 208676 468 208728 474
rect 208676 410 208728 416
rect 192574 368 192630 377
rect 184572 332 184624 338
rect 192574 303 192630 312
rect 208306 368 208362 377
rect 208306 303 208362 312
rect 184572 274 184624 280
rect 209516 202 209544 1158
rect 209792 1057 209820 1838
rect 209778 1048 209834 1057
rect 209778 983 209834 992
rect 209884 542 209912 3538
rect 209962 3224 210018 3233
rect 209962 3159 210018 3168
rect 209976 3058 210004 3159
rect 209964 3052 210016 3058
rect 209964 2994 210016 3000
rect 209976 2854 210004 2994
rect 209964 2848 210016 2854
rect 209964 2790 210016 2796
rect 210068 1358 210096 9318
rect 210332 7812 210384 7818
rect 210332 7754 210384 7760
rect 210344 6662 210372 7754
rect 210424 7744 210476 7750
rect 210424 7686 210476 7692
rect 210436 7546 210464 7686
rect 210424 7540 210476 7546
rect 210424 7482 210476 7488
rect 210516 7472 210568 7478
rect 210516 7414 210568 7420
rect 210424 7200 210476 7206
rect 210424 7142 210476 7148
rect 210436 6934 210464 7142
rect 210528 6934 210556 7414
rect 210424 6928 210476 6934
rect 210424 6870 210476 6876
rect 210516 6928 210568 6934
rect 210516 6870 210568 6876
rect 210332 6656 210384 6662
rect 210332 6598 210384 6604
rect 210424 5908 210476 5914
rect 210424 5850 210476 5856
rect 210436 5574 210464 5850
rect 210424 5568 210476 5574
rect 210424 5510 210476 5516
rect 210332 5228 210384 5234
rect 210332 5170 210384 5176
rect 210148 4752 210200 4758
rect 210148 4694 210200 4700
rect 210160 4554 210188 4694
rect 210148 4548 210200 4554
rect 210148 4490 210200 4496
rect 210160 4282 210188 4490
rect 210344 4486 210372 5170
rect 210516 4616 210568 4622
rect 210516 4558 210568 4564
rect 210240 4480 210292 4486
rect 210240 4422 210292 4428
rect 210332 4480 210384 4486
rect 210332 4422 210384 4428
rect 210148 4276 210200 4282
rect 210148 4218 210200 4224
rect 210252 3516 210280 4422
rect 210528 3534 210556 4558
rect 210332 3528 210384 3534
rect 210252 3488 210332 3516
rect 210332 3470 210384 3476
rect 210516 3528 210568 3534
rect 210516 3470 210568 3476
rect 210148 3460 210200 3466
rect 210148 3402 210200 3408
rect 210160 3058 210188 3402
rect 210148 3052 210200 3058
rect 210148 2994 210200 3000
rect 210160 1426 210188 2994
rect 210712 2038 210740 9318
rect 211264 8022 211292 10134
rect 212538 10095 212594 10104
rect 211710 9888 211766 9897
rect 211710 9823 211766 9832
rect 211724 8974 211752 9823
rect 212552 9586 212580 10095
rect 213472 9586 213500 10503
rect 216586 10432 216642 10441
rect 216586 10367 216588 10376
rect 216640 10367 216642 10376
rect 216588 10338 216640 10344
rect 213918 10160 213974 10169
rect 213918 10095 213974 10104
rect 214470 10160 214526 10169
rect 214470 10095 214526 10104
rect 216678 10160 216734 10169
rect 216678 10095 216734 10104
rect 213932 9586 213960 10095
rect 214484 9586 214512 10095
rect 216588 9988 216640 9994
rect 216588 9930 216640 9936
rect 215206 9752 215262 9761
rect 215206 9687 215208 9696
rect 215260 9687 215262 9696
rect 215208 9658 215260 9664
rect 215482 9616 215538 9625
rect 212540 9580 212592 9586
rect 212540 9522 212592 9528
rect 213460 9580 213512 9586
rect 213460 9522 213512 9528
rect 213920 9580 213972 9586
rect 213920 9522 213972 9528
rect 214472 9580 214524 9586
rect 215482 9551 215484 9560
rect 214472 9522 214524 9528
rect 215536 9551 215538 9560
rect 215484 9522 215536 9528
rect 215024 9444 215076 9450
rect 215024 9386 215076 9392
rect 215116 9444 215168 9450
rect 215116 9386 215168 9392
rect 212448 9376 212500 9382
rect 212448 9318 212500 9324
rect 212632 9376 212684 9382
rect 212632 9318 212684 9324
rect 213276 9376 213328 9382
rect 213276 9318 213328 9324
rect 214840 9376 214892 9382
rect 214840 9318 214892 9324
rect 211712 8968 211764 8974
rect 211712 8910 211764 8916
rect 211804 8968 211856 8974
rect 211804 8910 211856 8916
rect 211816 8362 211844 8910
rect 211804 8356 211856 8362
rect 211804 8298 211856 8304
rect 211252 8016 211304 8022
rect 211252 7958 211304 7964
rect 211160 7880 211212 7886
rect 211160 7822 211212 7828
rect 210976 3528 211028 3534
rect 210976 3470 211028 3476
rect 210988 3194 211016 3470
rect 210976 3188 211028 3194
rect 210976 3130 211028 3136
rect 211172 2922 211200 7822
rect 211436 7472 211488 7478
rect 211436 7414 211488 7420
rect 211448 4690 211476 7414
rect 212172 4752 212224 4758
rect 212170 4720 212172 4729
rect 212224 4720 212226 4729
rect 211436 4684 211488 4690
rect 212170 4655 212226 4664
rect 211436 4626 211488 4632
rect 211344 4616 211396 4622
rect 211620 4616 211672 4622
rect 211344 4558 211396 4564
rect 211540 4576 211620 4604
rect 211356 3738 211384 4558
rect 211344 3732 211396 3738
rect 211344 3674 211396 3680
rect 211356 3534 211384 3674
rect 211540 3534 211568 4576
rect 211620 4558 211672 4564
rect 211712 4616 211764 4622
rect 211712 4558 211764 4564
rect 211724 3534 211752 4558
rect 212080 4072 212132 4078
rect 212080 4014 212132 4020
rect 211804 4004 211856 4010
rect 211804 3946 211856 3952
rect 211344 3528 211396 3534
rect 211528 3528 211580 3534
rect 211344 3470 211396 3476
rect 211448 3488 211528 3516
rect 211356 3058 211384 3470
rect 211448 3398 211476 3488
rect 211528 3470 211580 3476
rect 211712 3528 211764 3534
rect 211712 3470 211764 3476
rect 211436 3392 211488 3398
rect 211436 3334 211488 3340
rect 211528 3392 211580 3398
rect 211724 3346 211752 3470
rect 211528 3334 211580 3340
rect 211448 3058 211476 3334
rect 211540 3097 211568 3334
rect 211632 3318 211752 3346
rect 211632 3194 211660 3318
rect 211620 3188 211672 3194
rect 211620 3130 211672 3136
rect 211526 3088 211582 3097
rect 211344 3052 211396 3058
rect 211344 2994 211396 3000
rect 211436 3052 211488 3058
rect 211632 3058 211660 3130
rect 211526 3023 211582 3032
rect 211620 3052 211672 3058
rect 211436 2994 211488 3000
rect 211620 2994 211672 3000
rect 211160 2916 211212 2922
rect 211160 2858 211212 2864
rect 210700 2032 210752 2038
rect 210700 1974 210752 1980
rect 211356 1970 211384 2994
rect 211448 1970 211476 2994
rect 211632 1970 211660 2994
rect 211344 1964 211396 1970
rect 211344 1906 211396 1912
rect 211436 1964 211488 1970
rect 211436 1906 211488 1912
rect 211620 1964 211672 1970
rect 211620 1906 211672 1912
rect 210240 1760 210292 1766
rect 210240 1702 210292 1708
rect 210700 1760 210752 1766
rect 210700 1702 210752 1708
rect 210148 1420 210200 1426
rect 210148 1362 210200 1368
rect 210252 1358 210280 1702
rect 210712 1494 210740 1702
rect 210700 1488 210752 1494
rect 210700 1430 210752 1436
rect 210056 1352 210108 1358
rect 210056 1294 210108 1300
rect 210240 1352 210292 1358
rect 210240 1294 210292 1300
rect 210976 1352 211028 1358
rect 210976 1294 211028 1300
rect 211068 1352 211120 1358
rect 211068 1294 211120 1300
rect 209872 536 209924 542
rect 209872 478 209924 484
rect 210988 241 211016 1294
rect 210974 232 211030 241
rect 209504 196 209556 202
rect 211080 202 211108 1294
rect 211816 1193 211844 3946
rect 212092 3670 212120 4014
rect 212080 3664 212132 3670
rect 212080 3606 212132 3612
rect 212356 3460 212408 3466
rect 212356 3402 212408 3408
rect 211988 3120 212040 3126
rect 211988 3062 212040 3068
rect 211896 2372 211948 2378
rect 211896 2314 211948 2320
rect 211908 1562 211936 2314
rect 212000 2038 212028 3062
rect 212368 3058 212396 3402
rect 212356 3052 212408 3058
rect 212356 2994 212408 3000
rect 212356 2440 212408 2446
rect 212356 2382 212408 2388
rect 211988 2032 212040 2038
rect 211988 1974 212040 1980
rect 211896 1556 211948 1562
rect 211896 1498 211948 1504
rect 211802 1184 211858 1193
rect 211802 1119 211858 1128
rect 211908 1057 211936 1498
rect 212368 1222 212396 2382
rect 212460 1358 212488 9318
rect 212644 4690 212672 9318
rect 213182 7304 213238 7313
rect 213182 7239 213238 7248
rect 213196 6798 213224 7239
rect 213184 6792 213236 6798
rect 213184 6734 213236 6740
rect 213090 6352 213146 6361
rect 213090 6287 213092 6296
rect 213144 6287 213146 6296
rect 213092 6258 213144 6264
rect 212816 6248 212868 6254
rect 212816 6190 212868 6196
rect 212828 5817 212856 6190
rect 212814 5808 212870 5817
rect 212814 5743 212870 5752
rect 212828 5710 212856 5743
rect 212816 5704 212868 5710
rect 212816 5646 212868 5652
rect 213182 5536 213238 5545
rect 213182 5471 213238 5480
rect 213196 5234 213224 5471
rect 213288 5234 213316 9318
rect 214010 9208 214066 9217
rect 214010 9143 214066 9152
rect 213920 8560 213972 8566
rect 213920 8502 213972 8508
rect 213552 7948 213604 7954
rect 213552 7890 213604 7896
rect 213458 7440 213514 7449
rect 213458 7375 213460 7384
rect 213512 7375 213514 7384
rect 213460 7346 213512 7352
rect 213368 7336 213420 7342
rect 213368 7278 213420 7284
rect 213380 5846 213408 7278
rect 213564 6798 213592 7890
rect 213932 7857 213960 8502
rect 214024 8265 214052 9143
rect 214564 8832 214616 8838
rect 214564 8774 214616 8780
rect 214010 8256 214066 8265
rect 214010 8191 214066 8200
rect 214194 8120 214250 8129
rect 214194 8055 214250 8064
rect 213918 7848 213974 7857
rect 213828 7812 213880 7818
rect 213918 7783 213974 7792
rect 213828 7754 213880 7760
rect 213734 7032 213790 7041
rect 213734 6967 213790 6976
rect 213552 6792 213604 6798
rect 213552 6734 213604 6740
rect 213644 6724 213696 6730
rect 213644 6666 213696 6672
rect 213460 6180 213512 6186
rect 213460 6122 213512 6128
rect 213472 5846 213500 6122
rect 213368 5840 213420 5846
rect 213368 5782 213420 5788
rect 213460 5840 213512 5846
rect 213460 5782 213512 5788
rect 213380 5710 213408 5782
rect 213656 5710 213684 6666
rect 213368 5704 213420 5710
rect 213368 5646 213420 5652
rect 213644 5704 213696 5710
rect 213644 5646 213696 5652
rect 213184 5228 213236 5234
rect 213184 5170 213236 5176
rect 213276 5228 213328 5234
rect 213276 5170 213328 5176
rect 213552 5160 213604 5166
rect 213552 5102 213604 5108
rect 213460 5092 213512 5098
rect 213460 5034 213512 5040
rect 213472 4690 213500 5034
rect 212632 4684 212684 4690
rect 212632 4626 212684 4632
rect 213460 4684 213512 4690
rect 213460 4626 213512 4632
rect 213000 4616 213052 4622
rect 213000 4558 213052 4564
rect 213012 3738 213040 4558
rect 213184 4140 213236 4146
rect 213184 4082 213236 4088
rect 213196 4010 213224 4082
rect 213184 4004 213236 4010
rect 213184 3946 213236 3952
rect 213000 3732 213052 3738
rect 213000 3674 213052 3680
rect 213000 3528 213052 3534
rect 213000 3470 213052 3476
rect 213012 3194 213040 3470
rect 213000 3188 213052 3194
rect 213000 3130 213052 3136
rect 213460 3188 213512 3194
rect 213460 3130 213512 3136
rect 212540 3052 212592 3058
rect 212540 2994 212592 3000
rect 212552 2514 212580 2994
rect 213000 2984 213052 2990
rect 213000 2926 213052 2932
rect 213012 2854 213040 2926
rect 213000 2848 213052 2854
rect 213000 2790 213052 2796
rect 212540 2508 212592 2514
rect 212540 2450 212592 2456
rect 213368 1896 213420 1902
rect 213472 1884 213500 3130
rect 213420 1856 213500 1884
rect 213368 1838 213420 1844
rect 213092 1828 213144 1834
rect 213092 1770 213144 1776
rect 213104 1426 213132 1770
rect 213564 1442 213592 5102
rect 213748 4622 213776 6967
rect 213736 4616 213788 4622
rect 213736 4558 213788 4564
rect 213736 3392 213788 3398
rect 213736 3334 213788 3340
rect 213642 2272 213698 2281
rect 213642 2207 213698 2216
rect 213656 1970 213684 2207
rect 213644 1964 213696 1970
rect 213644 1906 213696 1912
rect 213748 1766 213776 3334
rect 213840 3194 213868 7754
rect 213920 6996 213972 7002
rect 213920 6938 213972 6944
rect 213932 6662 213960 6938
rect 213920 6656 213972 6662
rect 213920 6598 213972 6604
rect 214104 5364 214156 5370
rect 214104 5306 214156 5312
rect 214116 5166 214144 5306
rect 214104 5160 214156 5166
rect 214104 5102 214156 5108
rect 214012 5024 214064 5030
rect 214012 4966 214064 4972
rect 214024 4622 214052 4966
rect 214012 4616 214064 4622
rect 214012 4558 214064 4564
rect 213920 4072 213972 4078
rect 213920 4014 213972 4020
rect 213828 3188 213880 3194
rect 213828 3130 213880 3136
rect 213828 2984 213880 2990
rect 213828 2926 213880 2932
rect 213840 2514 213868 2926
rect 213828 2508 213880 2514
rect 213828 2450 213880 2456
rect 213828 1964 213880 1970
rect 213828 1906 213880 1912
rect 213736 1760 213788 1766
rect 213736 1702 213788 1708
rect 213092 1420 213144 1426
rect 213564 1414 213684 1442
rect 213840 1426 213868 1906
rect 213092 1362 213144 1368
rect 212448 1352 212500 1358
rect 212448 1294 212500 1300
rect 212632 1352 212684 1358
rect 212632 1294 212684 1300
rect 213368 1352 213420 1358
rect 213368 1294 213420 1300
rect 213552 1352 213604 1358
rect 213552 1294 213604 1300
rect 212356 1216 212408 1222
rect 212356 1158 212408 1164
rect 211894 1048 211950 1057
rect 211894 983 211950 992
rect 212644 610 212672 1294
rect 212632 604 212684 610
rect 212632 546 212684 552
rect 212998 368 213054 377
rect 212998 303 213000 312
rect 213052 303 213054 312
rect 213000 274 213052 280
rect 210974 167 211030 176
rect 211068 196 211120 202
rect 209504 138 209556 144
rect 211068 138 211120 144
rect 213380 105 213408 1294
rect 213564 882 213592 1294
rect 213460 876 213512 882
rect 213460 818 213512 824
rect 213552 876 213604 882
rect 213552 818 213604 824
rect 213472 610 213500 818
rect 213656 814 213684 1414
rect 213828 1420 213880 1426
rect 213828 1362 213880 1368
rect 213644 808 213696 814
rect 213644 750 213696 756
rect 213460 604 213512 610
rect 213460 546 213512 552
rect 213932 270 213960 4014
rect 214208 3670 214236 8055
rect 214288 7268 214340 7274
rect 214288 7210 214340 7216
rect 214196 3664 214248 3670
rect 214196 3606 214248 3612
rect 214012 3528 214064 3534
rect 214012 3470 214064 3476
rect 214024 1873 214052 3470
rect 214300 2990 214328 7210
rect 214470 5536 214526 5545
rect 214470 5471 214526 5480
rect 214378 5400 214434 5409
rect 214378 5335 214434 5344
rect 214392 5234 214420 5335
rect 214484 5234 214512 5471
rect 214380 5228 214432 5234
rect 214380 5170 214432 5176
rect 214472 5228 214524 5234
rect 214472 5170 214524 5176
rect 214378 4856 214434 4865
rect 214576 4842 214604 8774
rect 214576 4814 214696 4842
rect 214378 4791 214434 4800
rect 214288 2984 214340 2990
rect 214288 2926 214340 2932
rect 214392 2446 214420 4791
rect 214564 4752 214616 4758
rect 214564 4694 214616 4700
rect 214576 2553 214604 4694
rect 214562 2544 214618 2553
rect 214562 2479 214618 2488
rect 214380 2440 214432 2446
rect 214378 2408 214380 2417
rect 214432 2408 214434 2417
rect 214378 2343 214434 2352
rect 214472 2304 214524 2310
rect 214472 2246 214524 2252
rect 214484 2038 214512 2246
rect 214472 2032 214524 2038
rect 214472 1974 214524 1980
rect 214668 1970 214696 4814
rect 214746 4720 214802 4729
rect 214746 4655 214748 4664
rect 214800 4655 214802 4664
rect 214748 4626 214800 4632
rect 214656 1964 214708 1970
rect 214656 1906 214708 1912
rect 214010 1864 214066 1873
rect 214010 1799 214066 1808
rect 214852 1766 214880 9318
rect 214932 2984 214984 2990
rect 214932 2926 214984 2932
rect 214840 1760 214892 1766
rect 214562 1728 214618 1737
rect 214840 1702 214892 1708
rect 214562 1663 214618 1672
rect 214576 474 214604 1663
rect 214656 1216 214708 1222
rect 214656 1158 214708 1164
rect 214668 950 214696 1158
rect 214944 1018 214972 2926
rect 215036 1358 215064 9386
rect 215128 8974 215156 9386
rect 215116 8968 215168 8974
rect 215116 8910 215168 8916
rect 216404 8628 216456 8634
rect 216404 8570 216456 8576
rect 215484 8560 215536 8566
rect 215484 8502 215536 8508
rect 215208 8492 215260 8498
rect 215208 8434 215260 8440
rect 215220 6202 215248 8434
rect 215300 7200 215352 7206
rect 215300 7142 215352 7148
rect 215128 6174 215248 6202
rect 215128 5574 215156 6174
rect 215312 5896 215340 7142
rect 215312 5868 215432 5896
rect 215208 5704 215260 5710
rect 215208 5646 215260 5652
rect 215116 5568 215168 5574
rect 215116 5510 215168 5516
rect 215116 5092 215168 5098
rect 215116 5034 215168 5040
rect 215128 4486 215156 5034
rect 215116 4480 215168 4486
rect 215116 4422 215168 4428
rect 215220 4049 215248 5646
rect 215404 5166 215432 5868
rect 215392 5160 215444 5166
rect 215392 5102 215444 5108
rect 215300 5024 215352 5030
rect 215300 4966 215352 4972
rect 215206 4040 215262 4049
rect 215312 4010 215340 4966
rect 215206 3975 215262 3984
rect 215300 4004 215352 4010
rect 215300 3946 215352 3952
rect 215392 3664 215444 3670
rect 215392 3606 215444 3612
rect 215116 3460 215168 3466
rect 215116 3402 215168 3408
rect 215128 3126 215156 3402
rect 215116 3120 215168 3126
rect 215116 3062 215168 3068
rect 215404 2990 215432 3606
rect 215392 2984 215444 2990
rect 215392 2926 215444 2932
rect 215496 1902 215524 8502
rect 216128 6792 216180 6798
rect 216128 6734 216180 6740
rect 216036 6384 216088 6390
rect 216036 6326 216088 6332
rect 215852 6112 215904 6118
rect 215852 6054 215904 6060
rect 215864 5778 215892 6054
rect 215852 5772 215904 5778
rect 215852 5714 215904 5720
rect 216048 5642 216076 6326
rect 216036 5636 216088 5642
rect 216036 5578 216088 5584
rect 216140 5302 216168 6734
rect 216312 6724 216364 6730
rect 216312 6666 216364 6672
rect 216324 6322 216352 6666
rect 216312 6316 216364 6322
rect 216312 6258 216364 6264
rect 216416 6225 216444 8570
rect 216600 8265 216628 9930
rect 216692 9586 216720 10095
rect 216862 9888 216918 9897
rect 216862 9823 216918 9832
rect 216680 9580 216732 9586
rect 216680 9522 216732 9528
rect 216770 9072 216826 9081
rect 216770 9007 216826 9016
rect 216586 8256 216642 8265
rect 216586 8191 216642 8200
rect 216496 6656 216548 6662
rect 216496 6598 216548 6604
rect 216508 6458 216536 6598
rect 216496 6452 216548 6458
rect 216496 6394 216548 6400
rect 216588 6452 216640 6458
rect 216588 6394 216640 6400
rect 216402 6216 216458 6225
rect 216402 6151 216458 6160
rect 216600 6089 216628 6394
rect 216784 6186 216812 9007
rect 216876 8974 216904 9823
rect 217508 9376 217560 9382
rect 217508 9318 217560 9324
rect 217784 9376 217836 9382
rect 217784 9318 217836 9324
rect 216864 8968 216916 8974
rect 216864 8910 216916 8916
rect 217322 8392 217378 8401
rect 217322 8327 217378 8336
rect 216864 7404 216916 7410
rect 216864 7346 216916 7352
rect 216876 6866 216904 7346
rect 216864 6860 216916 6866
rect 216864 6802 216916 6808
rect 217336 6798 217364 8327
rect 217324 6792 217376 6798
rect 217324 6734 217376 6740
rect 217048 6656 217100 6662
rect 217048 6598 217100 6604
rect 217060 6254 217088 6598
rect 217336 6390 217364 6734
rect 217324 6384 217376 6390
rect 217324 6326 217376 6332
rect 217048 6248 217100 6254
rect 217048 6190 217100 6196
rect 216772 6180 216824 6186
rect 216772 6122 216824 6128
rect 216586 6080 216642 6089
rect 216586 6015 216642 6024
rect 216680 5908 216732 5914
rect 216680 5850 216732 5856
rect 216586 5808 216642 5817
rect 216586 5743 216642 5752
rect 216496 5704 216548 5710
rect 216402 5672 216458 5681
rect 216496 5646 216548 5652
rect 216402 5607 216458 5616
rect 216220 5568 216272 5574
rect 216220 5510 216272 5516
rect 216128 5296 216180 5302
rect 216128 5238 216180 5244
rect 215576 5228 215628 5234
rect 215576 5170 215628 5176
rect 215944 5228 215996 5234
rect 215944 5170 215996 5176
rect 215588 4214 215616 5170
rect 215850 4992 215906 5001
rect 215850 4927 215906 4936
rect 215576 4208 215628 4214
rect 215576 4150 215628 4156
rect 215588 3534 215616 4150
rect 215576 3528 215628 3534
rect 215576 3470 215628 3476
rect 215864 1970 215892 4927
rect 215956 4282 215984 5170
rect 216232 4486 216260 5510
rect 216312 5228 216364 5234
rect 216312 5170 216364 5176
rect 216324 5098 216352 5170
rect 216312 5092 216364 5098
rect 216312 5034 216364 5040
rect 216220 4480 216272 4486
rect 216220 4422 216272 4428
rect 215944 4276 215996 4282
rect 215944 4218 215996 4224
rect 216324 4214 216352 5034
rect 216416 4554 216444 5607
rect 216508 5302 216536 5646
rect 216600 5522 216628 5743
rect 216692 5642 216720 5850
rect 217060 5778 217088 6190
rect 217140 6180 217192 6186
rect 217140 6122 217192 6128
rect 217048 5772 217100 5778
rect 217048 5714 217100 5720
rect 216680 5636 216732 5642
rect 216680 5578 216732 5584
rect 217152 5574 217180 6122
rect 217232 5636 217284 5642
rect 217232 5578 217284 5584
rect 217140 5568 217192 5574
rect 216600 5494 216904 5522
rect 217140 5510 217192 5516
rect 216496 5296 216548 5302
rect 216496 5238 216548 5244
rect 216772 4820 216824 4826
rect 216772 4762 216824 4768
rect 216404 4548 216456 4554
rect 216404 4490 216456 4496
rect 216784 4282 216812 4762
rect 216772 4276 216824 4282
rect 216772 4218 216824 4224
rect 216312 4208 216364 4214
rect 216312 4150 216364 4156
rect 216588 4072 216640 4078
rect 216588 4014 216640 4020
rect 216680 4072 216732 4078
rect 216680 4014 216732 4020
rect 216036 3936 216088 3942
rect 216036 3878 216088 3884
rect 216048 3670 216076 3878
rect 216036 3664 216088 3670
rect 216036 3606 216088 3612
rect 216496 3528 216548 3534
rect 216496 3470 216548 3476
rect 216508 2854 216536 3470
rect 216600 3398 216628 4014
rect 216692 3534 216720 4014
rect 216680 3528 216732 3534
rect 216680 3470 216732 3476
rect 216588 3392 216640 3398
rect 216588 3334 216640 3340
rect 216772 3120 216824 3126
rect 216772 3062 216824 3068
rect 216680 2916 216732 2922
rect 216680 2858 216732 2864
rect 216496 2848 216548 2854
rect 216496 2790 216548 2796
rect 215942 2408 215998 2417
rect 215942 2343 215998 2352
rect 215852 1964 215904 1970
rect 215852 1906 215904 1912
rect 215484 1896 215536 1902
rect 215484 1838 215536 1844
rect 215576 1828 215628 1834
rect 215576 1770 215628 1776
rect 215588 1426 215616 1770
rect 215576 1420 215628 1426
rect 215576 1362 215628 1368
rect 215024 1352 215076 1358
rect 215024 1294 215076 1300
rect 214932 1012 214984 1018
rect 214932 954 214984 960
rect 214656 944 214708 950
rect 214656 886 214708 892
rect 215956 746 215984 2343
rect 216034 2136 216090 2145
rect 216692 2106 216720 2858
rect 216784 2514 216812 3062
rect 216876 2553 216904 5494
rect 217152 5370 217180 5510
rect 217140 5364 217192 5370
rect 217140 5306 217192 5312
rect 217140 5228 217192 5234
rect 217140 5170 217192 5176
rect 216956 5024 217008 5030
rect 216956 4966 217008 4972
rect 216968 4146 216996 4966
rect 217048 4548 217100 4554
rect 217048 4490 217100 4496
rect 216956 4140 217008 4146
rect 216956 4082 217008 4088
rect 217060 3505 217088 4490
rect 217046 3496 217102 3505
rect 217046 3431 217102 3440
rect 217152 2961 217180 5170
rect 217244 4826 217272 5578
rect 217232 4820 217284 4826
rect 217232 4762 217284 4768
rect 217416 3936 217468 3942
rect 217416 3878 217468 3884
rect 217428 3602 217456 3878
rect 217416 3596 217468 3602
rect 217416 3538 217468 3544
rect 217138 2952 217194 2961
rect 217138 2887 217194 2896
rect 216862 2544 216918 2553
rect 216772 2508 216824 2514
rect 217520 2514 217548 9318
rect 217692 8832 217744 8838
rect 217692 8774 217744 8780
rect 217704 4078 217732 8774
rect 217796 5234 217824 9318
rect 217888 6866 217916 10678
rect 218796 10668 218848 10674
rect 218796 10610 218848 10616
rect 218610 10568 218666 10577
rect 218610 10503 218666 10512
rect 217966 10160 218022 10169
rect 217966 10095 218022 10104
rect 217980 9586 218008 10095
rect 218520 9716 218572 9722
rect 218520 9658 218572 9664
rect 217968 9580 218020 9586
rect 217968 9522 218020 9528
rect 218428 9376 218480 9382
rect 218428 9318 218480 9324
rect 217968 8832 218020 8838
rect 217968 8774 218020 8780
rect 217980 8566 218008 8774
rect 217968 8560 218020 8566
rect 217968 8502 218020 8508
rect 217968 7336 218020 7342
rect 217968 7278 218020 7284
rect 217876 6860 217928 6866
rect 217876 6802 217928 6808
rect 217876 6316 217928 6322
rect 217876 6258 217928 6264
rect 217888 5710 217916 6258
rect 217980 5914 218008 7278
rect 218058 6896 218114 6905
rect 218058 6831 218114 6840
rect 218244 6860 218296 6866
rect 218072 6322 218100 6831
rect 218244 6802 218296 6808
rect 218060 6316 218112 6322
rect 218060 6258 218112 6264
rect 217968 5908 218020 5914
rect 217968 5850 218020 5856
rect 217876 5704 217928 5710
rect 217876 5646 217928 5652
rect 218072 5642 218100 6258
rect 218152 6112 218204 6118
rect 218152 6054 218204 6060
rect 218060 5636 218112 5642
rect 218060 5578 218112 5584
rect 217784 5228 217836 5234
rect 217784 5170 217836 5176
rect 218072 5114 218100 5578
rect 217888 5086 218100 5114
rect 217888 4214 217916 5086
rect 217968 5024 218020 5030
rect 217968 4966 218020 4972
rect 217980 4690 218008 4966
rect 218164 4690 218192 6054
rect 217968 4684 218020 4690
rect 217968 4626 218020 4632
rect 218152 4684 218204 4690
rect 218152 4626 218204 4632
rect 217968 4548 218020 4554
rect 217968 4490 218020 4496
rect 217876 4208 217928 4214
rect 217876 4150 217928 4156
rect 217692 4072 217744 4078
rect 217692 4014 217744 4020
rect 217980 4010 218008 4490
rect 218152 4072 218204 4078
rect 218256 4049 218284 6802
rect 218334 6760 218390 6769
rect 218334 6695 218390 6704
rect 218348 6254 218376 6695
rect 218440 6322 218468 9318
rect 218428 6316 218480 6322
rect 218428 6258 218480 6264
rect 218336 6248 218388 6254
rect 218336 6190 218388 6196
rect 218348 5710 218376 6190
rect 218428 5908 218480 5914
rect 218428 5850 218480 5856
rect 218336 5704 218388 5710
rect 218336 5646 218388 5652
rect 218440 5250 218468 5850
rect 218348 5222 218468 5250
rect 218348 4554 218376 5222
rect 218428 5160 218480 5166
rect 218428 5102 218480 5108
rect 218440 4690 218468 5102
rect 218428 4684 218480 4690
rect 218428 4626 218480 4632
rect 218336 4548 218388 4554
rect 218336 4490 218388 4496
rect 218428 4548 218480 4554
rect 218428 4490 218480 4496
rect 218440 4078 218468 4490
rect 218428 4072 218480 4078
rect 218152 4014 218204 4020
rect 218242 4040 218298 4049
rect 217968 4004 218020 4010
rect 217968 3946 218020 3952
rect 217968 3664 218020 3670
rect 217968 3606 218020 3612
rect 217692 3460 217744 3466
rect 217692 3402 217744 3408
rect 217704 3233 217732 3402
rect 217690 3224 217746 3233
rect 217690 3159 217746 3168
rect 217876 2848 217928 2854
rect 217876 2790 217928 2796
rect 217600 2644 217652 2650
rect 217600 2586 217652 2592
rect 217612 2514 217640 2586
rect 216862 2479 216918 2488
rect 217508 2508 217560 2514
rect 216772 2450 216824 2456
rect 217508 2450 217560 2456
rect 217600 2508 217652 2514
rect 217600 2450 217652 2456
rect 216034 2071 216090 2080
rect 216588 2100 216640 2106
rect 216048 1970 216076 2071
rect 216588 2042 216640 2048
rect 216680 2100 216732 2106
rect 216680 2042 216732 2048
rect 216036 1964 216088 1970
rect 216036 1906 216088 1912
rect 216128 1896 216180 1902
rect 216126 1864 216128 1873
rect 216180 1864 216182 1873
rect 216126 1799 216182 1808
rect 216402 1864 216458 1873
rect 216402 1799 216458 1808
rect 216416 1358 216444 1799
rect 216600 1562 216628 2042
rect 216588 1556 216640 1562
rect 216588 1498 216640 1504
rect 216128 1352 216180 1358
rect 216128 1294 216180 1300
rect 216312 1352 216364 1358
rect 216312 1294 216364 1300
rect 216404 1352 216456 1358
rect 216404 1294 216456 1300
rect 216140 950 216168 1294
rect 216128 944 216180 950
rect 216128 886 216180 892
rect 216140 746 216168 886
rect 215944 740 215996 746
rect 215944 682 215996 688
rect 216128 740 216180 746
rect 216128 682 216180 688
rect 215574 640 215630 649
rect 215574 575 215630 584
rect 214564 468 214616 474
rect 214564 410 214616 416
rect 214472 400 214524 406
rect 214470 368 214472 377
rect 215588 377 215616 575
rect 216324 474 216352 1294
rect 216680 944 216732 950
rect 216680 886 216732 892
rect 216692 513 216720 886
rect 216784 610 216812 2450
rect 217692 2440 217744 2446
rect 217692 2382 217744 2388
rect 217048 1216 217100 1222
rect 217048 1158 217100 1164
rect 217060 1018 217088 1158
rect 217048 1012 217100 1018
rect 217048 954 217100 960
rect 217704 610 217732 2382
rect 217888 1358 217916 2790
rect 217980 1494 218008 3606
rect 218164 2582 218192 4014
rect 218428 4014 218480 4020
rect 218242 3975 218298 3984
rect 218532 3670 218560 9658
rect 218624 9586 218652 10503
rect 218612 9580 218664 9586
rect 218612 9522 218664 9528
rect 218704 6656 218756 6662
rect 218704 6598 218756 6604
rect 218612 6180 218664 6186
rect 218612 6122 218664 6128
rect 218624 5166 218652 6122
rect 218716 6118 218744 6598
rect 218704 6112 218756 6118
rect 218704 6054 218756 6060
rect 218612 5160 218664 5166
rect 218612 5102 218664 5108
rect 218716 4554 218744 6054
rect 218808 5914 218836 10610
rect 219072 10396 219124 10402
rect 219072 10338 219124 10344
rect 219084 8090 219112 10338
rect 219254 10160 219310 10169
rect 219254 10095 219310 10104
rect 219268 9586 219296 10095
rect 219256 9580 219308 9586
rect 219256 9522 219308 9528
rect 219912 9518 219940 10746
rect 220084 10532 220136 10538
rect 220084 10474 220136 10480
rect 219992 10056 220044 10062
rect 219992 9998 220044 10004
rect 220004 9518 220032 9998
rect 220096 9994 220124 10474
rect 220084 9988 220136 9994
rect 220084 9930 220136 9936
rect 220188 9926 220216 10814
rect 223486 10568 223542 10577
rect 223486 10503 223488 10512
rect 223540 10503 223542 10512
rect 223488 10474 223540 10480
rect 223580 10464 223632 10470
rect 221830 10432 221886 10441
rect 223580 10406 223632 10412
rect 221830 10367 221886 10376
rect 220358 10296 220414 10305
rect 220358 10231 220414 10240
rect 220176 9920 220228 9926
rect 220176 9862 220228 9868
rect 220268 9920 220320 9926
rect 220268 9862 220320 9868
rect 220084 9716 220136 9722
rect 220084 9658 220136 9664
rect 219900 9512 219952 9518
rect 219900 9454 219952 9460
rect 219992 9512 220044 9518
rect 219992 9454 220044 9460
rect 219348 9376 219400 9382
rect 219348 9318 219400 9324
rect 219256 8560 219308 8566
rect 219256 8502 219308 8508
rect 219164 8356 219216 8362
rect 219164 8298 219216 8304
rect 219072 8084 219124 8090
rect 219072 8026 219124 8032
rect 218980 8016 219032 8022
rect 218980 7958 219032 7964
rect 218992 6633 219020 7958
rect 219070 7712 219126 7721
rect 219070 7647 219126 7656
rect 219084 7041 219112 7647
rect 219176 7478 219204 8298
rect 219268 7886 219296 8502
rect 219256 7880 219308 7886
rect 219256 7822 219308 7828
rect 219164 7472 219216 7478
rect 219164 7414 219216 7420
rect 219256 7472 219308 7478
rect 219256 7414 219308 7420
rect 219070 7032 219126 7041
rect 219070 6967 219126 6976
rect 219164 6792 219216 6798
rect 219164 6734 219216 6740
rect 218978 6624 219034 6633
rect 218978 6559 219034 6568
rect 218980 6248 219032 6254
rect 218980 6190 219032 6196
rect 218992 5914 219020 6190
rect 218796 5908 218848 5914
rect 218796 5850 218848 5856
rect 218980 5908 219032 5914
rect 218980 5850 219032 5856
rect 218796 5704 218848 5710
rect 218796 5646 218848 5652
rect 218808 5234 218836 5646
rect 218796 5228 218848 5234
rect 218796 5170 218848 5176
rect 218980 5160 219032 5166
rect 218980 5102 219032 5108
rect 218992 4729 219020 5102
rect 218978 4720 219034 4729
rect 218978 4655 219034 4664
rect 219072 4684 219124 4690
rect 219072 4626 219124 4632
rect 218704 4548 218756 4554
rect 218704 4490 218756 4496
rect 218888 4548 218940 4554
rect 218888 4490 218940 4496
rect 218704 4072 218756 4078
rect 218704 4014 218756 4020
rect 218796 4072 218848 4078
rect 218796 4014 218848 4020
rect 218716 3738 218744 4014
rect 218704 3732 218756 3738
rect 218704 3674 218756 3680
rect 218520 3664 218572 3670
rect 218520 3606 218572 3612
rect 218808 3194 218836 4014
rect 218900 3777 218928 4490
rect 219084 4321 219112 4626
rect 219070 4312 219126 4321
rect 219070 4247 219126 4256
rect 219176 4078 219204 6734
rect 219268 6730 219296 7414
rect 219256 6724 219308 6730
rect 219256 6666 219308 6672
rect 219254 5944 219310 5953
rect 219254 5879 219310 5888
rect 219268 4185 219296 5879
rect 219254 4176 219310 4185
rect 219254 4111 219310 4120
rect 219360 4078 219388 9318
rect 220096 9042 220124 9658
rect 220176 9648 220228 9654
rect 220176 9590 220228 9596
rect 220188 9042 220216 9590
rect 220280 9110 220308 9862
rect 220372 9654 220400 10231
rect 220542 10160 220598 10169
rect 220542 10095 220598 10104
rect 220452 10056 220504 10062
rect 220452 9998 220504 10004
rect 220360 9648 220412 9654
rect 220360 9590 220412 9596
rect 220360 9376 220412 9382
rect 220360 9318 220412 9324
rect 220268 9104 220320 9110
rect 220268 9046 220320 9052
rect 220084 9036 220136 9042
rect 220084 8978 220136 8984
rect 220176 9036 220228 9042
rect 220176 8978 220228 8984
rect 219440 8628 219492 8634
rect 219440 8570 219492 8576
rect 219452 7857 219480 8570
rect 219438 7848 219494 7857
rect 219438 7783 219494 7792
rect 220082 7576 220138 7585
rect 220082 7511 220138 7520
rect 219440 7268 219492 7274
rect 219440 7210 219492 7216
rect 219452 6089 219480 7210
rect 220096 7177 220124 7511
rect 220082 7168 220138 7177
rect 220082 7103 220138 7112
rect 219624 6860 219676 6866
rect 219624 6802 219676 6808
rect 219532 6656 219584 6662
rect 219532 6598 219584 6604
rect 219544 6254 219572 6598
rect 219532 6248 219584 6254
rect 219532 6190 219584 6196
rect 219438 6080 219494 6089
rect 219438 6015 219494 6024
rect 219532 5704 219584 5710
rect 219532 5646 219584 5652
rect 219438 5264 219494 5273
rect 219438 5199 219494 5208
rect 219452 4690 219480 5199
rect 219544 5098 219572 5646
rect 219532 5092 219584 5098
rect 219532 5034 219584 5040
rect 219440 4684 219492 4690
rect 219440 4626 219492 4632
rect 219452 4457 219480 4626
rect 219532 4548 219584 4554
rect 219532 4490 219584 4496
rect 219438 4448 219494 4457
rect 219438 4383 219494 4392
rect 219544 4162 219572 4490
rect 219452 4134 219572 4162
rect 218980 4072 219032 4078
rect 218980 4014 219032 4020
rect 219164 4072 219216 4078
rect 219164 4014 219216 4020
rect 219348 4072 219400 4078
rect 219348 4014 219400 4020
rect 218886 3768 218942 3777
rect 218886 3703 218942 3712
rect 218796 3188 218848 3194
rect 218796 3130 218848 3136
rect 218428 3120 218480 3126
rect 218428 3062 218480 3068
rect 218440 2990 218468 3062
rect 218336 2984 218388 2990
rect 218336 2926 218388 2932
rect 218428 2984 218480 2990
rect 218992 2972 219020 4014
rect 219452 3890 219480 4134
rect 219360 3862 219480 3890
rect 219164 3460 219216 3466
rect 219164 3402 219216 3408
rect 219176 3369 219204 3402
rect 219162 3360 219218 3369
rect 219162 3295 219218 3304
rect 218428 2926 218480 2932
rect 218716 2944 219020 2972
rect 218152 2576 218204 2582
rect 218152 2518 218204 2524
rect 218164 1834 218192 2518
rect 218152 1828 218204 1834
rect 218152 1770 218204 1776
rect 217968 1488 218020 1494
rect 217968 1430 218020 1436
rect 217980 1358 218008 1430
rect 218164 1426 218192 1770
rect 218348 1578 218376 2926
rect 218716 2446 218744 2944
rect 218428 2440 218480 2446
rect 218428 2382 218480 2388
rect 218612 2440 218664 2446
rect 218612 2382 218664 2388
rect 218704 2440 218756 2446
rect 218704 2382 218756 2388
rect 218440 2106 218468 2382
rect 218428 2100 218480 2106
rect 218428 2042 218480 2048
rect 218348 1550 218468 1578
rect 218334 1456 218390 1465
rect 218152 1420 218204 1426
rect 218334 1391 218336 1400
rect 218152 1362 218204 1368
rect 218388 1391 218390 1400
rect 218336 1362 218388 1368
rect 217876 1352 217928 1358
rect 217876 1294 217928 1300
rect 217968 1352 218020 1358
rect 218060 1352 218112 1358
rect 217968 1294 218020 1300
rect 218058 1320 218060 1329
rect 218244 1352 218296 1358
rect 218112 1320 218114 1329
rect 218244 1294 218296 1300
rect 218058 1255 218114 1264
rect 218060 1012 218112 1018
rect 218060 954 218112 960
rect 218072 785 218100 954
rect 218058 776 218114 785
rect 218058 711 218114 720
rect 216772 604 216824 610
rect 216772 546 216824 552
rect 217692 604 217744 610
rect 217692 546 217744 552
rect 216678 504 216734 513
rect 216312 468 216364 474
rect 216678 439 216734 448
rect 216312 410 216364 416
rect 214524 368 214526 377
rect 214470 303 214526 312
rect 215574 368 215630 377
rect 218256 338 218284 1294
rect 218440 1222 218468 1550
rect 218428 1216 218480 1222
rect 218428 1158 218480 1164
rect 215574 303 215630 312
rect 218244 332 218296 338
rect 218244 274 218296 280
rect 218624 270 218652 2382
rect 218704 1964 218756 1970
rect 218900 1952 218928 2944
rect 218980 1964 219032 1970
rect 218756 1924 218836 1952
rect 218704 1906 218756 1912
rect 218704 1216 218756 1222
rect 218704 1158 218756 1164
rect 218716 814 218744 1158
rect 218704 808 218756 814
rect 218704 750 218756 756
rect 218808 338 218836 1924
rect 218900 1924 218980 1952
rect 218900 1873 218928 1924
rect 218980 1906 219032 1912
rect 218886 1864 218942 1873
rect 218886 1799 218942 1808
rect 219176 649 219204 3295
rect 219360 2990 219388 3862
rect 219532 3664 219584 3670
rect 219532 3606 219584 3612
rect 219348 2984 219400 2990
rect 219348 2926 219400 2932
rect 219256 2916 219308 2922
rect 219256 2858 219308 2864
rect 219268 2650 219296 2858
rect 219256 2644 219308 2650
rect 219256 2586 219308 2592
rect 219544 1902 219572 3606
rect 219636 3466 219664 6802
rect 219900 6248 219952 6254
rect 219898 6216 219900 6225
rect 219952 6216 219954 6225
rect 219898 6151 219954 6160
rect 219808 6112 219860 6118
rect 219808 6054 219860 6060
rect 220176 6112 220228 6118
rect 220176 6054 220228 6060
rect 219716 5568 219768 5574
rect 219716 5510 219768 5516
rect 219728 5302 219756 5510
rect 219716 5296 219768 5302
rect 219716 5238 219768 5244
rect 219820 4010 219848 6054
rect 219990 5672 220046 5681
rect 219990 5607 220046 5616
rect 220084 5636 220136 5642
rect 219900 5364 219952 5370
rect 219900 5306 219952 5312
rect 219808 4004 219860 4010
rect 219808 3946 219860 3952
rect 219912 3670 219940 5306
rect 220004 4758 220032 5607
rect 220084 5578 220136 5584
rect 220096 5302 220124 5578
rect 220084 5296 220136 5302
rect 220084 5238 220136 5244
rect 220188 5234 220216 6054
rect 220176 5228 220228 5234
rect 220176 5170 220228 5176
rect 219992 4752 220044 4758
rect 219992 4694 220044 4700
rect 220372 4690 220400 9318
rect 220464 8498 220492 9998
rect 220556 9586 220584 10095
rect 221844 9586 221872 10367
rect 223118 10160 223174 10169
rect 223118 10095 223174 10104
rect 222014 9888 222070 9897
rect 222014 9823 222070 9832
rect 220544 9580 220596 9586
rect 220544 9522 220596 9528
rect 221832 9580 221884 9586
rect 221832 9522 221884 9528
rect 221004 9376 221056 9382
rect 221004 9318 221056 9324
rect 221648 9376 221700 9382
rect 221648 9318 221700 9324
rect 220542 8800 220598 8809
rect 220542 8735 220598 8744
rect 220452 8492 220504 8498
rect 220452 8434 220504 8440
rect 220450 6760 220506 6769
rect 220450 6695 220506 6704
rect 220464 6186 220492 6695
rect 220452 6180 220504 6186
rect 220452 6122 220504 6128
rect 220556 4865 220584 8735
rect 220912 8628 220964 8634
rect 220912 8570 220964 8576
rect 220818 8528 220874 8537
rect 220818 8463 220874 8472
rect 220832 7750 220860 8463
rect 220820 7744 220872 7750
rect 220820 7686 220872 7692
rect 220924 7562 220952 8570
rect 220832 7534 220952 7562
rect 220832 7002 220860 7534
rect 220820 6996 220872 7002
rect 220820 6938 220872 6944
rect 220728 6248 220780 6254
rect 220728 6190 220780 6196
rect 220636 5296 220688 5302
rect 220636 5238 220688 5244
rect 220542 4856 220598 4865
rect 220542 4791 220598 4800
rect 220360 4684 220412 4690
rect 220360 4626 220412 4632
rect 220648 4554 220676 5238
rect 220740 5166 220768 6190
rect 220832 5778 220860 6938
rect 220820 5772 220872 5778
rect 220820 5714 220872 5720
rect 220728 5160 220780 5166
rect 220728 5102 220780 5108
rect 220820 5160 220872 5166
rect 220820 5102 220872 5108
rect 220832 4758 220860 5102
rect 220912 5092 220964 5098
rect 220912 5034 220964 5040
rect 220820 4752 220872 4758
rect 220820 4694 220872 4700
rect 220728 4616 220780 4622
rect 220832 4593 220860 4694
rect 220728 4558 220780 4564
rect 220818 4584 220874 4593
rect 220636 4548 220688 4554
rect 220636 4490 220688 4496
rect 220176 4480 220228 4486
rect 220176 4422 220228 4428
rect 220268 4480 220320 4486
rect 220268 4422 220320 4428
rect 219900 3664 219952 3670
rect 219900 3606 219952 3612
rect 219624 3460 219676 3466
rect 219624 3402 219676 3408
rect 219636 2990 219664 3402
rect 219624 2984 219676 2990
rect 219624 2926 219676 2932
rect 219898 2680 219954 2689
rect 219898 2615 219954 2624
rect 219624 2304 219676 2310
rect 219624 2246 219676 2252
rect 219716 2304 219768 2310
rect 219716 2246 219768 2252
rect 219636 2106 219664 2246
rect 219624 2100 219676 2106
rect 219624 2042 219676 2048
rect 219348 1896 219400 1902
rect 219346 1864 219348 1873
rect 219532 1896 219584 1902
rect 219400 1864 219402 1873
rect 219532 1838 219584 1844
rect 219346 1799 219402 1808
rect 219440 1828 219492 1834
rect 219440 1770 219492 1776
rect 219452 1562 219480 1770
rect 219532 1760 219584 1766
rect 219532 1702 219584 1708
rect 219544 1562 219572 1702
rect 219440 1556 219492 1562
rect 219440 1498 219492 1504
rect 219532 1556 219584 1562
rect 219532 1498 219584 1504
rect 219728 1465 219756 2246
rect 219912 2009 219940 2615
rect 219898 2000 219954 2009
rect 219898 1935 219954 1944
rect 220082 2000 220138 2009
rect 220188 1970 220216 4422
rect 220280 4146 220308 4422
rect 220268 4140 220320 4146
rect 220268 4082 220320 4088
rect 220740 4010 220768 4558
rect 220818 4519 220874 4528
rect 220924 4282 220952 5034
rect 221016 4282 221044 9318
rect 221660 9042 221688 9318
rect 221648 9036 221700 9042
rect 221648 8978 221700 8984
rect 222028 8974 222056 9823
rect 223132 9586 223160 10095
rect 223120 9580 223172 9586
rect 223120 9522 223172 9528
rect 222936 9376 222988 9382
rect 222936 9318 222988 9324
rect 222016 8968 222068 8974
rect 222016 8910 222068 8916
rect 221280 8832 221332 8838
rect 221280 8774 221332 8780
rect 221292 8430 221320 8774
rect 221464 8492 221516 8498
rect 221464 8434 221516 8440
rect 221280 8424 221332 8430
rect 221280 8366 221332 8372
rect 221096 8084 221148 8090
rect 221096 8026 221148 8032
rect 221108 6662 221136 8026
rect 221476 7546 221504 8434
rect 221464 7540 221516 7546
rect 221464 7482 221516 7488
rect 221924 7540 221976 7546
rect 221924 7482 221976 7488
rect 221280 6996 221332 7002
rect 221280 6938 221332 6944
rect 221096 6656 221148 6662
rect 221096 6598 221148 6604
rect 220912 4276 220964 4282
rect 220912 4218 220964 4224
rect 221004 4276 221056 4282
rect 221004 4218 221056 4224
rect 221004 4072 221056 4078
rect 221004 4014 221056 4020
rect 221188 4072 221240 4078
rect 221188 4014 221240 4020
rect 220360 4004 220412 4010
rect 220360 3946 220412 3952
rect 220728 4004 220780 4010
rect 220728 3946 220780 3952
rect 220082 1935 220138 1944
rect 220176 1964 220228 1970
rect 220096 1737 220124 1935
rect 220176 1906 220228 1912
rect 220372 1902 220400 3946
rect 220818 3768 220874 3777
rect 220818 3703 220874 3712
rect 220832 3466 220860 3703
rect 220820 3460 220872 3466
rect 220820 3402 220872 3408
rect 220912 3460 220964 3466
rect 220912 3402 220964 3408
rect 220924 3194 220952 3402
rect 220912 3188 220964 3194
rect 220912 3130 220964 3136
rect 220636 3052 220688 3058
rect 220636 2994 220688 3000
rect 220544 2916 220596 2922
rect 220544 2858 220596 2864
rect 220556 2446 220584 2858
rect 220648 2854 220676 2994
rect 220820 2984 220872 2990
rect 221016 2961 221044 4014
rect 221096 3936 221148 3942
rect 221096 3878 221148 3884
rect 221108 3602 221136 3878
rect 221200 3670 221228 4014
rect 221188 3664 221240 3670
rect 221188 3606 221240 3612
rect 221096 3596 221148 3602
rect 221096 3538 221148 3544
rect 220820 2926 220872 2932
rect 221002 2952 221058 2961
rect 220636 2848 220688 2854
rect 220636 2790 220688 2796
rect 220648 2446 220676 2790
rect 220832 2446 220860 2926
rect 221002 2887 221058 2896
rect 221292 2774 221320 6938
rect 221830 6896 221886 6905
rect 221830 6831 221886 6840
rect 221556 6384 221608 6390
rect 221556 6326 221608 6332
rect 221372 6316 221424 6322
rect 221372 6258 221424 6264
rect 221384 5370 221412 6258
rect 221372 5364 221424 5370
rect 221372 5306 221424 5312
rect 221384 3602 221412 5306
rect 221372 3596 221424 3602
rect 221372 3538 221424 3544
rect 221384 3058 221412 3538
rect 221464 3460 221516 3466
rect 221464 3402 221516 3408
rect 221476 3233 221504 3402
rect 221462 3224 221518 3233
rect 221462 3159 221518 3168
rect 221372 3052 221424 3058
rect 221372 2994 221424 3000
rect 221384 2922 221412 2994
rect 221372 2916 221424 2922
rect 221424 2876 221504 2904
rect 221372 2858 221424 2864
rect 221016 2746 221320 2774
rect 220544 2440 220596 2446
rect 220544 2382 220596 2388
rect 220636 2440 220688 2446
rect 220636 2382 220688 2388
rect 220820 2440 220872 2446
rect 220820 2382 220872 2388
rect 220360 1896 220412 1902
rect 220360 1838 220412 1844
rect 220452 1828 220504 1834
rect 220452 1770 220504 1776
rect 220082 1728 220138 1737
rect 220082 1663 220138 1672
rect 220464 1562 220492 1770
rect 220452 1556 220504 1562
rect 220452 1498 220504 1504
rect 220648 1494 220676 2382
rect 220728 2100 220780 2106
rect 220728 2042 220780 2048
rect 220740 1494 220768 2042
rect 220636 1488 220688 1494
rect 219714 1456 219770 1465
rect 220636 1430 220688 1436
rect 220728 1488 220780 1494
rect 220728 1430 220780 1436
rect 219714 1391 219770 1400
rect 219532 1352 219584 1358
rect 219532 1294 219584 1300
rect 220544 1352 220596 1358
rect 220832 1329 220860 2382
rect 221016 1968 221044 2746
rect 221094 2544 221150 2553
rect 221094 2479 221150 2488
rect 221004 1962 221056 1968
rect 221004 1904 221056 1910
rect 220544 1294 220596 1300
rect 220818 1320 220874 1329
rect 219544 950 219572 1294
rect 219532 944 219584 950
rect 219532 886 219584 892
rect 219162 640 219218 649
rect 219162 575 219218 584
rect 220556 406 220584 1294
rect 220818 1255 220820 1264
rect 220872 1255 220874 1264
rect 220820 1226 220872 1232
rect 220820 808 220872 814
rect 220820 750 220872 756
rect 220544 400 220596 406
rect 220832 377 220860 750
rect 221108 377 221136 2479
rect 221372 2440 221424 2446
rect 221372 2382 221424 2388
rect 221384 2106 221412 2382
rect 221372 2100 221424 2106
rect 221372 2042 221424 2048
rect 221280 1964 221332 1970
rect 221332 1924 221412 1952
rect 221280 1906 221332 1912
rect 221384 1766 221412 1924
rect 221372 1760 221424 1766
rect 221372 1702 221424 1708
rect 221476 1358 221504 2876
rect 221568 2854 221596 6326
rect 221844 6322 221872 6831
rect 221740 6316 221792 6322
rect 221660 6276 221740 6304
rect 221660 6186 221688 6276
rect 221740 6258 221792 6264
rect 221832 6316 221884 6322
rect 221832 6258 221884 6264
rect 221648 6180 221700 6186
rect 221648 6122 221700 6128
rect 221660 3058 221688 6122
rect 221740 5160 221792 5166
rect 221740 5102 221792 5108
rect 221752 4690 221780 5102
rect 221740 4684 221792 4690
rect 221740 4626 221792 4632
rect 221738 4040 221794 4049
rect 221738 3975 221794 3984
rect 221648 3052 221700 3058
rect 221648 2994 221700 3000
rect 221660 2854 221688 2994
rect 221556 2848 221608 2854
rect 221556 2790 221608 2796
rect 221648 2848 221700 2854
rect 221648 2790 221700 2796
rect 221464 1352 221516 1358
rect 221660 1340 221688 2790
rect 221752 1737 221780 3975
rect 221844 3058 221872 6258
rect 221936 6236 221964 7482
rect 222014 7168 222070 7177
rect 222014 7103 222070 7112
rect 222028 6304 222056 7103
rect 222198 6488 222254 6497
rect 222198 6423 222200 6432
rect 222252 6423 222254 6432
rect 222200 6394 222252 6400
rect 222028 6276 222148 6304
rect 221936 6208 222056 6236
rect 222028 4622 222056 6208
rect 222120 4622 222148 6276
rect 222292 6248 222344 6254
rect 222292 6190 222344 6196
rect 222752 6248 222804 6254
rect 222752 6190 222804 6196
rect 222304 4622 222332 6190
rect 222764 5914 222792 6190
rect 222844 6180 222896 6186
rect 222844 6122 222896 6128
rect 222660 5908 222712 5914
rect 222660 5850 222712 5856
rect 222752 5908 222804 5914
rect 222752 5850 222804 5856
rect 222384 5092 222436 5098
rect 222384 5034 222436 5040
rect 222016 4616 222068 4622
rect 222016 4558 222068 4564
rect 222108 4616 222160 4622
rect 222108 4558 222160 4564
rect 222292 4616 222344 4622
rect 222292 4558 222344 4564
rect 222304 4486 222332 4558
rect 222108 4480 222160 4486
rect 222108 4422 222160 4428
rect 222292 4480 222344 4486
rect 222292 4422 222344 4428
rect 221924 4072 221976 4078
rect 221924 4014 221976 4020
rect 221832 3052 221884 3058
rect 221832 2994 221884 3000
rect 221832 2508 221884 2514
rect 221832 2450 221884 2456
rect 221844 2038 221872 2450
rect 221832 2032 221884 2038
rect 221832 1974 221884 1980
rect 221936 1766 221964 4014
rect 222120 3942 222148 4422
rect 222304 4078 222332 4422
rect 222292 4072 222344 4078
rect 222198 4040 222254 4049
rect 222292 4014 222344 4020
rect 222198 3975 222254 3984
rect 222108 3936 222160 3942
rect 222108 3878 222160 3884
rect 222106 3768 222162 3777
rect 222212 3754 222240 3975
rect 222162 3726 222240 3754
rect 222106 3703 222162 3712
rect 222014 3632 222070 3641
rect 222014 3567 222070 3576
rect 222028 2582 222056 3567
rect 222108 3392 222160 3398
rect 222108 3334 222160 3340
rect 222120 2774 222148 3334
rect 222120 2746 222240 2774
rect 222016 2576 222068 2582
rect 222016 2518 222068 2524
rect 222016 1964 222068 1970
rect 222016 1906 222068 1912
rect 221924 1760 221976 1766
rect 221738 1728 221794 1737
rect 221924 1702 221976 1708
rect 221738 1663 221794 1672
rect 222028 1426 222056 1906
rect 222016 1420 222068 1426
rect 222016 1362 222068 1368
rect 221740 1352 221792 1358
rect 221660 1312 221740 1340
rect 221464 1294 221516 1300
rect 222212 1329 222240 2746
rect 221740 1294 221792 1300
rect 222198 1320 222254 1329
rect 222198 1255 222254 1264
rect 222396 406 222424 5034
rect 222568 3596 222620 3602
rect 222568 3538 222620 3544
rect 222580 3233 222608 3538
rect 222566 3224 222622 3233
rect 222566 3159 222622 3168
rect 222580 2825 222608 3159
rect 222566 2816 222622 2825
rect 222566 2751 222622 2760
rect 222568 2372 222620 2378
rect 222568 2314 222620 2320
rect 222580 1465 222608 2314
rect 222672 2106 222700 5850
rect 222856 4826 222884 6122
rect 222948 5778 222976 9318
rect 223028 8968 223080 8974
rect 223028 8910 223080 8916
rect 222936 5772 222988 5778
rect 222936 5714 222988 5720
rect 222936 5160 222988 5166
rect 222936 5102 222988 5108
rect 222948 4826 222976 5102
rect 222844 4820 222896 4826
rect 222844 4762 222896 4768
rect 222936 4820 222988 4826
rect 222936 4762 222988 4768
rect 222856 4554 222884 4762
rect 222844 4548 222896 4554
rect 222844 4490 222896 4496
rect 222752 3596 222804 3602
rect 222752 3538 222804 3544
rect 222764 2854 222792 3538
rect 222752 2848 222804 2854
rect 222752 2790 222804 2796
rect 222660 2100 222712 2106
rect 222660 2042 222712 2048
rect 223040 1562 223068 8910
rect 223396 8832 223448 8838
rect 223396 8774 223448 8780
rect 223212 8560 223264 8566
rect 223212 8502 223264 8508
rect 223224 8129 223252 8502
rect 223302 8392 223358 8401
rect 223302 8327 223358 8336
rect 223210 8120 223266 8129
rect 223210 8055 223266 8064
rect 223316 6254 223344 8327
rect 223304 6248 223356 6254
rect 223304 6190 223356 6196
rect 223120 6112 223172 6118
rect 223120 6054 223172 6060
rect 223212 6112 223264 6118
rect 223212 6054 223264 6060
rect 223132 5302 223160 6054
rect 223224 5846 223252 6054
rect 223316 5846 223344 6190
rect 223212 5840 223264 5846
rect 223212 5782 223264 5788
rect 223304 5840 223356 5846
rect 223304 5782 223356 5788
rect 223212 5704 223264 5710
rect 223212 5646 223264 5652
rect 223304 5704 223356 5710
rect 223304 5646 223356 5652
rect 223120 5296 223172 5302
rect 223120 5238 223172 5244
rect 223120 4820 223172 4826
rect 223120 4762 223172 4768
rect 223132 4486 223160 4762
rect 223224 4622 223252 5646
rect 223212 4616 223264 4622
rect 223212 4558 223264 4564
rect 223120 4480 223172 4486
rect 223120 4422 223172 4428
rect 223118 4312 223174 4321
rect 223316 4282 223344 5646
rect 223118 4247 223174 4256
rect 223304 4276 223356 4282
rect 223132 2514 223160 4247
rect 223304 4218 223356 4224
rect 223304 4072 223356 4078
rect 223304 4014 223356 4020
rect 223120 2508 223172 2514
rect 223120 2450 223172 2456
rect 223028 1556 223080 1562
rect 223028 1498 223080 1504
rect 222566 1456 222622 1465
rect 222566 1391 222622 1400
rect 223120 1352 223172 1358
rect 223120 1294 223172 1300
rect 222936 1216 222988 1222
rect 222936 1158 222988 1164
rect 222948 610 222976 1158
rect 223132 1018 223160 1294
rect 223316 1018 223344 4014
rect 223408 3058 223436 8774
rect 223488 8628 223540 8634
rect 223488 8570 223540 8576
rect 223500 7041 223528 8570
rect 223592 7478 223620 10406
rect 223946 10160 224002 10169
rect 223946 10095 224002 10104
rect 223960 9586 223988 10095
rect 224776 9716 224828 9722
rect 224776 9658 224828 9664
rect 223764 9580 223816 9586
rect 223764 9522 223816 9528
rect 223948 9580 224000 9586
rect 224788 9568 224816 9658
rect 224868 9580 224920 9586
rect 224788 9540 224868 9568
rect 223948 9522 224000 9528
rect 224868 9522 224920 9528
rect 223776 9110 223804 9522
rect 224038 9480 224094 9489
rect 224038 9415 224094 9424
rect 224052 9382 224080 9415
rect 224040 9376 224092 9382
rect 224040 9318 224092 9324
rect 223672 9104 223724 9110
rect 223672 9046 223724 9052
rect 223764 9104 223816 9110
rect 223764 9046 223816 9052
rect 223684 7818 223712 9046
rect 224592 9036 224644 9042
rect 224592 8978 224644 8984
rect 224316 8968 224368 8974
rect 224316 8910 224368 8916
rect 224408 8968 224460 8974
rect 224408 8910 224460 8916
rect 224040 8492 224092 8498
rect 224040 8434 224092 8440
rect 223764 8424 223816 8430
rect 224052 8378 224080 8434
rect 223816 8372 224080 8378
rect 223764 8366 224080 8372
rect 224224 8424 224276 8430
rect 224328 8401 224356 8910
rect 224420 8566 224448 8910
rect 224500 8832 224552 8838
rect 224500 8774 224552 8780
rect 224408 8560 224460 8566
rect 224408 8502 224460 8508
rect 224512 8498 224540 8774
rect 224500 8492 224552 8498
rect 224500 8434 224552 8440
rect 224224 8366 224276 8372
rect 224314 8392 224370 8401
rect 223776 8350 224080 8366
rect 224236 8242 224264 8366
rect 224604 8378 224632 8978
rect 224682 8664 224738 8673
rect 224972 8634 225000 10814
rect 225144 10804 225196 10810
rect 225144 10746 225196 10752
rect 225052 9716 225104 9722
rect 225052 9658 225104 9664
rect 224682 8599 224684 8608
rect 224736 8599 224738 8608
rect 224960 8628 225012 8634
rect 224684 8570 224736 8576
rect 224960 8570 225012 8576
rect 225064 8480 225092 9658
rect 225156 8906 225184 10746
rect 226708 10668 226760 10674
rect 226708 10610 226760 10616
rect 226984 10668 227036 10674
rect 226984 10610 227036 10616
rect 229100 10668 229152 10674
rect 229100 10610 229152 10616
rect 225236 9376 225288 9382
rect 225236 9318 225288 9324
rect 225144 8900 225196 8906
rect 225144 8842 225196 8848
rect 224314 8327 224370 8336
rect 224512 8350 224632 8378
rect 224788 8452 225092 8480
rect 224788 8362 224816 8452
rect 224776 8356 224828 8362
rect 224512 8242 224540 8350
rect 224776 8298 224828 8304
rect 224868 8356 224920 8362
rect 224868 8298 224920 8304
rect 224236 8214 224540 8242
rect 224592 8288 224644 8294
rect 224592 8230 224644 8236
rect 224684 8288 224736 8294
rect 224880 8265 224908 8298
rect 224684 8230 224736 8236
rect 224866 8256 224922 8265
rect 224604 8129 224632 8230
rect 224590 8120 224646 8129
rect 224590 8055 224646 8064
rect 223762 7984 223818 7993
rect 223762 7919 223818 7928
rect 223856 7948 223908 7954
rect 223672 7812 223724 7818
rect 223672 7754 223724 7760
rect 223580 7472 223632 7478
rect 223580 7414 223632 7420
rect 223672 7200 223724 7206
rect 223672 7142 223724 7148
rect 223486 7032 223542 7041
rect 223486 6967 223542 6976
rect 223488 6656 223540 6662
rect 223488 6598 223540 6604
rect 223500 5778 223528 6598
rect 223488 5772 223540 5778
rect 223488 5714 223540 5720
rect 223500 5098 223528 5714
rect 223578 5672 223634 5681
rect 223578 5607 223634 5616
rect 223592 5098 223620 5607
rect 223488 5092 223540 5098
rect 223488 5034 223540 5040
rect 223580 5092 223632 5098
rect 223580 5034 223632 5040
rect 223500 4978 223528 5034
rect 223500 4950 223620 4978
rect 223488 4548 223540 4554
rect 223488 4490 223540 4496
rect 223500 3777 223528 4490
rect 223592 4078 223620 4950
rect 223684 4865 223712 7142
rect 223776 5370 223804 7919
rect 223856 7890 223908 7896
rect 223764 5364 223816 5370
rect 223764 5306 223816 5312
rect 223762 5264 223818 5273
rect 223762 5199 223818 5208
rect 223776 5166 223804 5199
rect 223764 5160 223816 5166
rect 223764 5102 223816 5108
rect 223670 4856 223726 4865
rect 223670 4791 223726 4800
rect 223764 4752 223816 4758
rect 223764 4694 223816 4700
rect 223776 4622 223804 4694
rect 223764 4616 223816 4622
rect 223764 4558 223816 4564
rect 223868 4112 223896 7890
rect 224040 7880 224092 7886
rect 224040 7822 224092 7828
rect 224052 5778 224080 7822
rect 224696 7546 224724 8230
rect 224866 8191 224922 8200
rect 224776 7812 224828 7818
rect 224880 7806 225092 7834
rect 224880 7800 224908 7806
rect 224828 7772 224908 7800
rect 224776 7754 224828 7760
rect 224960 7744 225012 7750
rect 224960 7686 225012 7692
rect 224684 7540 224736 7546
rect 224684 7482 224736 7488
rect 224592 7404 224644 7410
rect 224592 7346 224644 7352
rect 224604 7206 224632 7346
rect 224592 7200 224644 7206
rect 224592 7142 224644 7148
rect 224868 6928 224920 6934
rect 224868 6870 224920 6876
rect 224316 6860 224368 6866
rect 224316 6802 224368 6808
rect 224224 6792 224276 6798
rect 224224 6734 224276 6740
rect 224132 6724 224184 6730
rect 224132 6666 224184 6672
rect 224040 5772 224092 5778
rect 224040 5714 224092 5720
rect 224144 4758 224172 6666
rect 224132 4752 224184 4758
rect 224132 4694 224184 4700
rect 223960 4554 224172 4570
rect 223960 4548 224184 4554
rect 223960 4542 224132 4548
rect 223856 4106 223908 4112
rect 223580 4072 223632 4078
rect 223856 4048 223908 4054
rect 223580 4014 223632 4020
rect 223592 3924 223620 4014
rect 223592 3896 223712 3924
rect 223486 3768 223542 3777
rect 223486 3703 223542 3712
rect 223578 3496 223634 3505
rect 223578 3431 223634 3440
rect 223396 3052 223448 3058
rect 223396 2994 223448 3000
rect 223592 2774 223620 3431
rect 223684 2990 223712 3896
rect 223960 3602 223988 4542
rect 224132 4490 224184 4496
rect 224040 4480 224092 4486
rect 224040 4422 224092 4428
rect 223948 3596 224000 3602
rect 223948 3538 224000 3544
rect 224052 3534 224080 4422
rect 224132 4140 224184 4146
rect 224236 4128 224264 6734
rect 224328 5710 224356 6802
rect 224776 6792 224828 6798
rect 224880 6769 224908 6870
rect 224972 6798 225000 7686
rect 225064 7342 225092 7806
rect 225052 7336 225104 7342
rect 225052 7278 225104 7284
rect 224960 6792 225012 6798
rect 224776 6734 224828 6740
rect 224866 6760 224922 6769
rect 224788 6440 224816 6734
rect 224960 6734 225012 6740
rect 224866 6695 224922 6704
rect 224788 6412 225092 6440
rect 224408 6384 224460 6390
rect 224408 6326 224460 6332
rect 224316 5704 224368 5710
rect 224316 5646 224368 5652
rect 224328 4826 224356 5646
rect 224420 5234 224448 6326
rect 224592 6316 224644 6322
rect 224592 6258 224644 6264
rect 224880 6310 225000 6338
rect 224604 5953 224632 6258
rect 224776 6180 224828 6186
rect 224776 6122 224828 6128
rect 224590 5944 224646 5953
rect 224590 5879 224646 5888
rect 224788 5846 224816 6122
rect 224880 6118 224908 6310
rect 224868 6112 224920 6118
rect 224868 6054 224920 6060
rect 224776 5840 224828 5846
rect 224776 5782 224828 5788
rect 224972 5710 225000 6310
rect 225064 5914 225092 6412
rect 225248 6254 225276 9318
rect 225420 9104 225472 9110
rect 225420 9046 225472 9052
rect 225328 8832 225380 8838
rect 225328 8774 225380 8780
rect 225340 8498 225368 8774
rect 225328 8492 225380 8498
rect 225328 8434 225380 8440
rect 225432 7290 225460 9046
rect 225604 8968 225656 8974
rect 225604 8910 225656 8916
rect 226432 8968 226484 8974
rect 226432 8910 226484 8916
rect 225510 8664 225566 8673
rect 225510 8599 225512 8608
rect 225564 8599 225566 8608
rect 225512 8570 225564 8576
rect 225512 7880 225564 7886
rect 225510 7848 225512 7857
rect 225564 7848 225566 7857
rect 225510 7783 225566 7792
rect 225524 7478 225552 7783
rect 225512 7472 225564 7478
rect 225512 7414 225564 7420
rect 225432 7262 225552 7290
rect 225236 6248 225288 6254
rect 225236 6190 225288 6196
rect 225420 6248 225472 6254
rect 225420 6190 225472 6196
rect 225052 5908 225104 5914
rect 225052 5850 225104 5856
rect 224960 5704 225012 5710
rect 224960 5646 225012 5652
rect 224960 5296 225012 5302
rect 224960 5238 225012 5244
rect 224408 5228 224460 5234
rect 224408 5170 224460 5176
rect 224972 4826 225000 5238
rect 225144 5160 225196 5166
rect 225144 5102 225196 5108
rect 225236 5160 225288 5166
rect 225236 5102 225288 5108
rect 224316 4820 224368 4826
rect 224316 4762 224368 4768
rect 224960 4820 225012 4826
rect 224960 4762 225012 4768
rect 224684 4752 224736 4758
rect 224684 4694 224736 4700
rect 224592 4480 224644 4486
rect 224184 4100 224264 4128
rect 224328 4440 224592 4468
rect 224132 4082 224184 4088
rect 224224 3596 224276 3602
rect 224224 3538 224276 3544
rect 223764 3528 223816 3534
rect 223764 3470 223816 3476
rect 224040 3528 224092 3534
rect 224040 3470 224092 3476
rect 223776 3058 223804 3470
rect 223948 3392 224000 3398
rect 223948 3334 224000 3340
rect 223764 3052 223816 3058
rect 223764 2994 223816 3000
rect 223672 2984 223724 2990
rect 223672 2926 223724 2932
rect 223500 2746 223620 2774
rect 223396 1896 223448 1902
rect 223396 1838 223448 1844
rect 223408 1766 223436 1838
rect 223396 1760 223448 1766
rect 223396 1702 223448 1708
rect 223408 1562 223436 1702
rect 223396 1556 223448 1562
rect 223396 1498 223448 1504
rect 223500 1193 223528 2746
rect 223578 2544 223634 2553
rect 223578 2479 223634 2488
rect 223486 1184 223542 1193
rect 223486 1119 223542 1128
rect 223120 1012 223172 1018
rect 223120 954 223172 960
rect 223304 1012 223356 1018
rect 223304 954 223356 960
rect 223592 785 223620 2479
rect 223960 1358 223988 3334
rect 224132 2984 224184 2990
rect 224236 2972 224264 3538
rect 224328 3058 224356 4440
rect 224592 4422 224644 4428
rect 224696 4298 224724 4694
rect 224776 4616 224828 4622
rect 224776 4558 224828 4564
rect 224604 4270 224724 4298
rect 224604 3058 224632 4270
rect 224788 4146 224816 4558
rect 225156 4282 225184 5102
rect 225144 4276 225196 4282
rect 225144 4218 225196 4224
rect 224776 4140 224828 4146
rect 224776 4082 224828 4088
rect 224682 4040 224738 4049
rect 224682 3975 224738 3984
rect 224696 3738 224724 3975
rect 224776 3936 224828 3942
rect 224776 3878 224828 3884
rect 224684 3732 224736 3738
rect 224684 3674 224736 3680
rect 224316 3052 224368 3058
rect 224316 2994 224368 3000
rect 224592 3052 224644 3058
rect 224592 2994 224644 3000
rect 224184 2944 224264 2972
rect 224132 2926 224184 2932
rect 224498 2816 224554 2825
rect 224498 2751 224554 2760
rect 224512 2650 224540 2751
rect 224500 2644 224552 2650
rect 224500 2586 224552 2592
rect 224132 2440 224184 2446
rect 224132 2382 224184 2388
rect 224144 2106 224172 2382
rect 224224 2304 224276 2310
rect 224224 2246 224276 2252
rect 224132 2100 224184 2106
rect 224132 2042 224184 2048
rect 223948 1352 224000 1358
rect 223948 1294 224000 1300
rect 224236 1193 224264 2246
rect 224512 2106 224540 2586
rect 224788 2310 224816 3878
rect 224958 3768 225014 3777
rect 224958 3703 225014 3712
rect 224866 2952 224922 2961
rect 224866 2887 224922 2896
rect 224776 2304 224828 2310
rect 224776 2246 224828 2252
rect 224500 2100 224552 2106
rect 224500 2042 224552 2048
rect 224408 1964 224460 1970
rect 224408 1906 224460 1912
rect 224420 1426 224448 1906
rect 224512 1902 224540 2042
rect 224880 2009 224908 2887
rect 224866 2000 224922 2009
rect 224866 1935 224922 1944
rect 224500 1896 224552 1902
rect 224500 1838 224552 1844
rect 224408 1420 224460 1426
rect 224408 1362 224460 1368
rect 224776 1216 224828 1222
rect 224222 1184 224278 1193
rect 224776 1158 224828 1164
rect 224222 1119 224278 1128
rect 224788 785 224816 1158
rect 223578 776 223634 785
rect 223578 711 223634 720
rect 224774 776 224830 785
rect 224774 711 224830 720
rect 222936 604 222988 610
rect 222936 546 222988 552
rect 223028 604 223080 610
rect 223028 546 223080 552
rect 222384 400 222436 406
rect 220544 342 220596 348
rect 220818 368 220874 377
rect 218796 332 218848 338
rect 220818 303 220874 312
rect 221094 368 221150 377
rect 222384 342 222436 348
rect 221094 303 221150 312
rect 218796 274 218848 280
rect 223040 270 223068 546
rect 224972 270 225000 3703
rect 225248 3126 225276 5102
rect 225432 4758 225460 6190
rect 225420 4752 225472 4758
rect 225420 4694 225472 4700
rect 225420 4072 225472 4078
rect 225420 4014 225472 4020
rect 225236 3120 225288 3126
rect 225236 3062 225288 3068
rect 225432 2774 225460 4014
rect 225524 3534 225552 7262
rect 225512 3528 225564 3534
rect 225512 3470 225564 3476
rect 225340 2746 225460 2774
rect 225340 1290 225368 2746
rect 225418 2680 225474 2689
rect 225616 2666 225644 8910
rect 226064 8832 226116 8838
rect 226064 8774 226116 8780
rect 226076 8498 226104 8774
rect 226246 8664 226302 8673
rect 226246 8599 226248 8608
rect 226300 8599 226302 8608
rect 226248 8570 226300 8576
rect 226064 8492 226116 8498
rect 226064 8434 226116 8440
rect 226248 8424 226300 8430
rect 226248 8366 226300 8372
rect 226064 8016 226116 8022
rect 226064 7958 226116 7964
rect 226154 7984 226210 7993
rect 225696 7744 225748 7750
rect 225696 7686 225748 7692
rect 225708 5710 225736 7686
rect 225970 7576 226026 7585
rect 225970 7511 226026 7520
rect 225984 7177 226012 7511
rect 225786 7168 225842 7177
rect 225786 7103 225842 7112
rect 225970 7168 226026 7177
rect 225970 7103 226026 7112
rect 225800 6730 225828 7103
rect 225788 6724 225840 6730
rect 225788 6666 225840 6672
rect 225880 6180 225932 6186
rect 225880 6122 225932 6128
rect 225696 5704 225748 5710
rect 225696 5646 225748 5652
rect 225892 3602 225920 6122
rect 226076 6100 226104 7958
rect 226154 7919 226210 7928
rect 226168 7585 226196 7919
rect 226260 7857 226288 8366
rect 226340 8016 226392 8022
rect 226340 7958 226392 7964
rect 226246 7848 226302 7857
rect 226246 7783 226302 7792
rect 226154 7576 226210 7585
rect 226154 7511 226210 7520
rect 226156 6656 226208 6662
rect 226156 6598 226208 6604
rect 226168 6458 226196 6598
rect 226246 6488 226302 6497
rect 226156 6452 226208 6458
rect 226246 6423 226248 6432
rect 226156 6394 226208 6400
rect 226300 6423 226302 6432
rect 226248 6394 226300 6400
rect 226168 6322 226196 6394
rect 226156 6316 226208 6322
rect 226156 6258 226208 6264
rect 226248 6248 226300 6254
rect 226248 6190 226300 6196
rect 226156 6112 226208 6118
rect 226076 6072 226156 6100
rect 226156 6054 226208 6060
rect 226260 5817 226288 6190
rect 226246 5808 226302 5817
rect 226064 5772 226116 5778
rect 226246 5743 226302 5752
rect 226064 5714 226116 5720
rect 226076 5098 226104 5714
rect 226064 5092 226116 5098
rect 226064 5034 226116 5040
rect 225880 3596 225932 3602
rect 225880 3538 225932 3544
rect 226248 3596 226300 3602
rect 226352 3584 226380 7958
rect 226444 6440 226472 8910
rect 226720 6905 226748 10610
rect 226996 10334 227024 10610
rect 228640 10600 228692 10606
rect 228692 10548 228864 10554
rect 228640 10542 228864 10548
rect 228652 10538 228864 10542
rect 228652 10532 228876 10538
rect 228652 10526 228824 10532
rect 228824 10474 228876 10480
rect 226984 10328 227036 10334
rect 226984 10270 227036 10276
rect 227076 10328 227128 10334
rect 227076 10270 227128 10276
rect 227088 10198 227116 10270
rect 227076 10192 227128 10198
rect 227076 10134 227128 10140
rect 227168 10192 227220 10198
rect 227168 10134 227220 10140
rect 227180 9994 227208 10134
rect 229008 10124 229060 10130
rect 229008 10066 229060 10072
rect 229112 10112 229140 10610
rect 229192 10124 229244 10130
rect 229112 10084 229192 10112
rect 228732 10056 228784 10062
rect 228732 9998 228784 10004
rect 227168 9988 227220 9994
rect 227168 9930 227220 9936
rect 227812 9988 227864 9994
rect 227812 9930 227864 9936
rect 227180 8974 227208 9930
rect 227824 9586 227852 9930
rect 227812 9580 227864 9586
rect 227812 9522 227864 9528
rect 228364 9580 228416 9586
rect 228364 9522 228416 9528
rect 228456 9580 228508 9586
rect 228456 9522 228508 9528
rect 227258 9072 227314 9081
rect 227258 9007 227314 9016
rect 227168 8968 227220 8974
rect 227168 8910 227220 8916
rect 226800 8832 226852 8838
rect 226800 8774 226852 8780
rect 226812 8498 226840 8774
rect 226982 8664 227038 8673
rect 226982 8599 226984 8608
rect 227036 8599 227038 8608
rect 226984 8570 227036 8576
rect 226800 8492 226852 8498
rect 226800 8434 226852 8440
rect 226984 7200 227036 7206
rect 226984 7142 227036 7148
rect 226706 6896 226762 6905
rect 226616 6860 226668 6866
rect 226996 6866 227024 7142
rect 226706 6831 226762 6840
rect 226984 6860 227036 6866
rect 226616 6802 226668 6808
rect 226444 6412 226564 6440
rect 226432 6316 226484 6322
rect 226432 6258 226484 6264
rect 226444 5846 226472 6258
rect 226432 5840 226484 5846
rect 226432 5782 226484 5788
rect 226300 3556 226380 3584
rect 226248 3538 226300 3544
rect 225696 3528 225748 3534
rect 225696 3470 225748 3476
rect 225708 3194 225736 3470
rect 225880 3392 225932 3398
rect 225880 3334 225932 3340
rect 225696 3188 225748 3194
rect 225696 3130 225748 3136
rect 225788 3188 225840 3194
rect 225788 3130 225840 3136
rect 225474 2638 225644 2666
rect 225418 2615 225474 2624
rect 225432 2378 225460 2615
rect 225800 2582 225828 3130
rect 225892 3058 225920 3334
rect 225880 3052 225932 3058
rect 225880 2994 225932 3000
rect 225972 3052 226024 3058
rect 225972 2994 226024 3000
rect 225788 2576 225840 2582
rect 225788 2518 225840 2524
rect 225788 2440 225840 2446
rect 225788 2382 225840 2388
rect 225420 2372 225472 2378
rect 225420 2314 225472 2320
rect 225432 1902 225460 2314
rect 225696 2304 225748 2310
rect 225696 2246 225748 2252
rect 225420 1896 225472 1902
rect 225420 1838 225472 1844
rect 225512 1760 225564 1766
rect 225512 1702 225564 1708
rect 225524 1358 225552 1702
rect 225512 1352 225564 1358
rect 225512 1294 225564 1300
rect 225328 1284 225380 1290
rect 225328 1226 225380 1232
rect 225708 1193 225736 2246
rect 225800 2106 225828 2382
rect 225788 2100 225840 2106
rect 225788 2042 225840 2048
rect 225694 1184 225750 1193
rect 225694 1119 225750 1128
rect 225984 649 226012 2994
rect 226536 2774 226564 6412
rect 226628 5846 226656 6802
rect 226616 5840 226668 5846
rect 226616 5782 226668 5788
rect 226628 3516 226656 5782
rect 226720 4078 226748 6831
rect 226984 6802 227036 6808
rect 226800 6656 226852 6662
rect 226800 6598 226852 6604
rect 226812 6254 226840 6598
rect 226800 6248 226852 6254
rect 226800 6190 226852 6196
rect 227076 6112 227128 6118
rect 227076 6054 227128 6060
rect 226892 5908 226944 5914
rect 226892 5850 226944 5856
rect 226708 4072 226760 4078
rect 226708 4014 226760 4020
rect 226708 3528 226760 3534
rect 226628 3488 226708 3516
rect 226708 3470 226760 3476
rect 226444 2746 226564 2774
rect 226340 2304 226392 2310
rect 226340 2246 226392 2252
rect 226352 1465 226380 2246
rect 226444 2038 226472 2746
rect 226800 2440 226852 2446
rect 226800 2382 226852 2388
rect 226812 2106 226840 2382
rect 226800 2100 226852 2106
rect 226800 2042 226852 2048
rect 226432 2032 226484 2038
rect 226430 2000 226432 2009
rect 226484 2000 226486 2009
rect 226430 1935 226486 1944
rect 226444 1902 226472 1935
rect 226432 1896 226484 1902
rect 226432 1838 226484 1844
rect 226522 1728 226578 1737
rect 226522 1663 226578 1672
rect 226536 1465 226564 1663
rect 226338 1456 226394 1465
rect 226338 1391 226394 1400
rect 226522 1456 226578 1465
rect 226522 1391 226578 1400
rect 226432 1352 226484 1358
rect 226246 1320 226302 1329
rect 226302 1278 226380 1306
rect 226432 1294 226484 1300
rect 226246 1255 226302 1264
rect 226352 1222 226380 1278
rect 226248 1216 226300 1222
rect 226248 1158 226300 1164
rect 226340 1216 226392 1222
rect 226340 1158 226392 1164
rect 226260 1018 226288 1158
rect 226248 1012 226300 1018
rect 226248 954 226300 960
rect 226444 814 226472 1294
rect 226432 808 226484 814
rect 226432 750 226484 756
rect 226904 746 226932 5850
rect 227088 5642 227116 6054
rect 227076 5636 227128 5642
rect 227076 5578 227128 5584
rect 226984 4208 227036 4214
rect 226984 4150 227036 4156
rect 226996 2650 227024 4150
rect 226984 2644 227036 2650
rect 226984 2586 227036 2592
rect 227076 2644 227128 2650
rect 227076 2586 227128 2592
rect 227088 2417 227116 2586
rect 227074 2408 227130 2417
rect 227074 2343 227130 2352
rect 227076 1896 227128 1902
rect 227076 1838 227128 1844
rect 227088 1358 227116 1838
rect 227180 1426 227208 8910
rect 227272 4146 227300 9007
rect 227824 8498 227852 9522
rect 228270 9480 228326 9489
rect 228270 9415 228272 9424
rect 228324 9415 228326 9424
rect 228272 9386 228324 9392
rect 228086 9208 228142 9217
rect 228376 9178 228404 9522
rect 228086 9143 228142 9152
rect 228364 9172 228416 9178
rect 228100 8974 228128 9143
rect 228364 9114 228416 9120
rect 228088 8968 228140 8974
rect 228088 8910 228140 8916
rect 228100 8838 228128 8910
rect 228272 8900 228324 8906
rect 228272 8842 228324 8848
rect 228088 8832 228140 8838
rect 228008 8792 228088 8820
rect 227812 8492 227864 8498
rect 227812 8434 227864 8440
rect 227352 7880 227404 7886
rect 227352 7822 227404 7828
rect 227364 7546 227392 7822
rect 227352 7540 227404 7546
rect 227352 7482 227404 7488
rect 227536 7540 227588 7546
rect 227536 7482 227588 7488
rect 227350 7168 227406 7177
rect 227350 7103 227406 7112
rect 227364 4622 227392 7103
rect 227442 7032 227498 7041
rect 227442 6967 227498 6976
rect 227456 6186 227484 6967
rect 227444 6180 227496 6186
rect 227444 6122 227496 6128
rect 227444 5160 227496 5166
rect 227444 5102 227496 5108
rect 227352 4616 227404 4622
rect 227352 4558 227404 4564
rect 227260 4140 227312 4146
rect 227260 4082 227312 4088
rect 227456 4010 227484 5102
rect 227548 4486 227576 7482
rect 227628 6928 227680 6934
rect 227680 6888 227852 6916
rect 227628 6870 227680 6876
rect 227626 6760 227682 6769
rect 227626 6695 227682 6704
rect 227640 5846 227668 6695
rect 227628 5840 227680 5846
rect 227628 5782 227680 5788
rect 227720 5636 227772 5642
rect 227720 5578 227772 5584
rect 227628 5160 227680 5166
rect 227628 5102 227680 5108
rect 227640 4593 227668 5102
rect 227626 4584 227682 4593
rect 227626 4519 227682 4528
rect 227536 4480 227588 4486
rect 227536 4422 227588 4428
rect 227732 4321 227760 5578
rect 227824 4758 227852 6888
rect 227902 5944 227958 5953
rect 227902 5879 227958 5888
rect 227812 4752 227864 4758
rect 227812 4694 227864 4700
rect 227812 4616 227864 4622
rect 227810 4584 227812 4593
rect 227864 4584 227866 4593
rect 227810 4519 227866 4528
rect 227718 4312 227774 4321
rect 227718 4247 227774 4256
rect 227628 4072 227680 4078
rect 227628 4014 227680 4020
rect 227352 4004 227404 4010
rect 227352 3946 227404 3952
rect 227444 4004 227496 4010
rect 227444 3946 227496 3952
rect 227364 3670 227392 3946
rect 227352 3664 227404 3670
rect 227352 3606 227404 3612
rect 227456 3194 227484 3946
rect 227640 3777 227668 4014
rect 227626 3768 227682 3777
rect 227626 3703 227682 3712
rect 227628 3664 227680 3670
rect 227628 3606 227680 3612
rect 227718 3632 227774 3641
rect 227640 3369 227668 3606
rect 227718 3567 227774 3576
rect 227732 3534 227760 3567
rect 227720 3528 227772 3534
rect 227720 3470 227772 3476
rect 227720 3392 227772 3398
rect 227626 3360 227682 3369
rect 227720 3334 227772 3340
rect 227626 3295 227682 3304
rect 227444 3188 227496 3194
rect 227444 3130 227496 3136
rect 227732 3058 227760 3334
rect 227720 3052 227772 3058
rect 227720 2994 227772 3000
rect 227916 2417 227944 5879
rect 228008 3194 228036 8792
rect 228088 8774 228140 8780
rect 228284 8498 228312 8842
rect 228468 8634 228496 9522
rect 228548 9172 228600 9178
rect 228548 9114 228600 9120
rect 228560 8838 228588 9114
rect 228548 8832 228600 8838
rect 228548 8774 228600 8780
rect 228456 8628 228508 8634
rect 228456 8570 228508 8576
rect 228272 8492 228324 8498
rect 228272 8434 228324 8440
rect 228364 8356 228416 8362
rect 228364 8298 228416 8304
rect 228456 8356 228508 8362
rect 228456 8298 228508 8304
rect 228376 7993 228404 8298
rect 228362 7984 228418 7993
rect 228362 7919 228418 7928
rect 228088 4820 228140 4826
rect 228088 4762 228140 4768
rect 228272 4820 228324 4826
rect 228272 4762 228324 4768
rect 227996 3188 228048 3194
rect 227996 3130 228048 3136
rect 227902 2408 227958 2417
rect 227902 2343 227958 2352
rect 227996 2304 228048 2310
rect 227996 2246 228048 2252
rect 227260 1964 227312 1970
rect 227260 1906 227312 1912
rect 227272 1426 227300 1906
rect 227444 1760 227496 1766
rect 227444 1702 227496 1708
rect 227168 1420 227220 1426
rect 227168 1362 227220 1368
rect 227260 1420 227312 1426
rect 227260 1362 227312 1368
rect 227076 1352 227128 1358
rect 227076 1294 227128 1300
rect 226892 740 226944 746
rect 226892 682 226944 688
rect 227456 649 227484 1702
rect 228008 1193 228036 2246
rect 227994 1184 228050 1193
rect 227994 1119 228050 1128
rect 228100 814 228128 4762
rect 228180 3936 228232 3942
rect 228180 3878 228232 3884
rect 228192 3738 228220 3878
rect 228180 3732 228232 3738
rect 228180 3674 228232 3680
rect 228284 3618 228312 4762
rect 228192 3590 228312 3618
rect 228088 808 228140 814
rect 228088 750 228140 756
rect 225970 640 226026 649
rect 225970 575 226026 584
rect 227442 640 227498 649
rect 227442 575 227498 584
rect 228192 338 228220 3590
rect 228468 3516 228496 8298
rect 228640 5228 228692 5234
rect 228640 5170 228692 5176
rect 228546 3904 228602 3913
rect 228546 3839 228602 3848
rect 228284 3488 228496 3516
rect 228284 2650 228312 3488
rect 228364 3188 228416 3194
rect 228364 3130 228416 3136
rect 228272 2644 228324 2650
rect 228272 2586 228324 2592
rect 228376 2038 228404 3130
rect 228560 2774 228588 3839
rect 228468 2746 228588 2774
rect 228468 2582 228496 2746
rect 228456 2576 228508 2582
rect 228456 2518 228508 2524
rect 228456 2440 228508 2446
rect 228456 2382 228508 2388
rect 228468 2106 228496 2382
rect 228456 2100 228508 2106
rect 228456 2042 228508 2048
rect 228364 2032 228416 2038
rect 228364 1974 228416 1980
rect 228548 1760 228600 1766
rect 228548 1702 228600 1708
rect 228560 1358 228588 1702
rect 228548 1352 228600 1358
rect 228652 1329 228680 5170
rect 228744 3641 228772 9998
rect 229020 9654 229048 10066
rect 229008 9648 229060 9654
rect 229008 9590 229060 9596
rect 229006 9480 229062 9489
rect 229006 9415 229008 9424
rect 229060 9415 229062 9424
rect 229008 9386 229060 9392
rect 228824 8968 228876 8974
rect 229112 8956 229140 10084
rect 229192 10066 229244 10072
rect 229652 9920 229704 9926
rect 229652 9862 229704 9868
rect 229664 8974 229692 9862
rect 230676 9586 230704 10814
rect 233608 10804 233660 10810
rect 233608 10746 233660 10752
rect 233620 10538 233648 10746
rect 234712 10736 234764 10742
rect 234712 10678 234764 10684
rect 236644 10736 236696 10742
rect 236644 10678 236696 10684
rect 232780 10532 232832 10538
rect 232780 10474 232832 10480
rect 233608 10532 233660 10538
rect 233608 10474 233660 10480
rect 231860 10328 231912 10334
rect 231860 10270 231912 10276
rect 231952 10328 232004 10334
rect 231952 10270 232004 10276
rect 231872 10198 231900 10270
rect 231860 10192 231912 10198
rect 231860 10134 231912 10140
rect 230940 9920 230992 9926
rect 230940 9862 230992 9868
rect 231032 9920 231084 9926
rect 231032 9862 231084 9868
rect 230020 9580 230072 9586
rect 230020 9522 230072 9528
rect 230664 9580 230716 9586
rect 230664 9522 230716 9528
rect 230848 9580 230900 9586
rect 230848 9522 230900 9528
rect 229834 9480 229890 9489
rect 229834 9415 229836 9424
rect 229888 9415 229890 9424
rect 229836 9386 229888 9392
rect 230032 8974 230060 9522
rect 230296 9512 230348 9518
rect 230296 9454 230348 9460
rect 230308 9382 230336 9454
rect 230296 9376 230348 9382
rect 230296 9318 230348 9324
rect 230572 9104 230624 9110
rect 230572 9046 230624 9052
rect 228876 8928 229140 8956
rect 228824 8910 228876 8916
rect 229008 8832 229060 8838
rect 229008 8774 229060 8780
rect 229020 8498 229048 8774
rect 229008 8492 229060 8498
rect 229008 8434 229060 8440
rect 229112 8430 229140 8928
rect 229652 8968 229704 8974
rect 229652 8910 229704 8916
rect 230020 8968 230072 8974
rect 230020 8910 230072 8916
rect 230112 8968 230164 8974
rect 230112 8910 230164 8916
rect 229190 8664 229246 8673
rect 229190 8599 229192 8608
rect 229244 8599 229246 8608
rect 229192 8570 229244 8576
rect 230124 8498 230152 8910
rect 230204 8900 230256 8906
rect 230204 8842 230256 8848
rect 230216 8566 230244 8842
rect 230204 8560 230256 8566
rect 230204 8502 230256 8508
rect 230112 8492 230164 8498
rect 230112 8434 230164 8440
rect 228916 8424 228968 8430
rect 228916 8366 228968 8372
rect 229100 8424 229152 8430
rect 229100 8366 229152 8372
rect 229652 8424 229704 8430
rect 229652 8366 229704 8372
rect 228730 3632 228786 3641
rect 228730 3567 228786 3576
rect 228928 1970 228956 8366
rect 229006 5536 229062 5545
rect 229006 5471 229062 5480
rect 229020 4185 229048 5471
rect 229006 4176 229062 4185
rect 229006 4111 229062 4120
rect 229664 2774 229692 8366
rect 230584 8362 230612 9046
rect 230676 8906 230704 9522
rect 230860 8974 230888 9522
rect 230952 9178 230980 9862
rect 230940 9172 230992 9178
rect 230940 9114 230992 9120
rect 230848 8968 230900 8974
rect 230848 8910 230900 8916
rect 230664 8900 230716 8906
rect 230664 8842 230716 8848
rect 230952 8786 230980 9114
rect 230676 8758 230980 8786
rect 230572 8356 230624 8362
rect 230572 8298 230624 8304
rect 229744 7472 229796 7478
rect 229744 7414 229796 7420
rect 229756 7002 229784 7414
rect 229744 6996 229796 7002
rect 229744 6938 229796 6944
rect 229742 6488 229798 6497
rect 229742 6423 229798 6432
rect 229756 6225 229784 6423
rect 229742 6216 229798 6225
rect 229742 6151 229798 6160
rect 229836 4072 229888 4078
rect 229836 4014 229888 4020
rect 229744 3936 229796 3942
rect 229744 3878 229796 3884
rect 229756 3670 229784 3878
rect 229848 3670 229876 4014
rect 229744 3664 229796 3670
rect 229744 3606 229796 3612
rect 229836 3664 229888 3670
rect 229836 3606 229888 3612
rect 229926 3632 229982 3641
rect 229926 3567 229982 3576
rect 229744 3392 229796 3398
rect 229744 3334 229796 3340
rect 229756 2922 229784 3334
rect 229940 3233 229968 3567
rect 229926 3224 229982 3233
rect 229926 3159 229982 3168
rect 229744 2916 229796 2922
rect 229744 2858 229796 2864
rect 229664 2746 229784 2774
rect 229756 1970 229784 2746
rect 230572 2576 230624 2582
rect 230572 2518 230624 2524
rect 229928 2372 229980 2378
rect 229928 2314 229980 2320
rect 229836 2032 229888 2038
rect 229836 1974 229888 1980
rect 228916 1964 228968 1970
rect 228916 1906 228968 1912
rect 229744 1964 229796 1970
rect 229744 1906 229796 1912
rect 229848 1494 229876 1974
rect 229940 1970 229968 2314
rect 230020 2304 230072 2310
rect 230020 2246 230072 2252
rect 229928 1964 229980 1970
rect 229928 1906 229980 1912
rect 229836 1488 229888 1494
rect 229836 1430 229888 1436
rect 228548 1294 228600 1300
rect 228638 1320 228694 1329
rect 228638 1255 228694 1264
rect 228732 1216 228784 1222
rect 228732 1158 228784 1164
rect 229468 1216 229520 1222
rect 230032 1193 230060 2246
rect 230112 1760 230164 1766
rect 230112 1702 230164 1708
rect 230386 1728 230442 1737
rect 230124 1358 230152 1702
rect 230386 1663 230442 1672
rect 230296 1420 230348 1426
rect 230296 1362 230348 1368
rect 230112 1352 230164 1358
rect 230112 1294 230164 1300
rect 229468 1158 229520 1164
rect 230018 1184 230074 1193
rect 228744 649 228772 1158
rect 229480 649 229508 1158
rect 230018 1119 230074 1128
rect 228730 640 228786 649
rect 228730 575 228786 584
rect 229466 640 229522 649
rect 229466 575 229522 584
rect 230202 504 230258 513
rect 230202 439 230258 448
rect 228180 332 228232 338
rect 228180 274 228232 280
rect 213920 264 213972 270
rect 213920 206 213972 212
rect 218612 264 218664 270
rect 218612 206 218664 212
rect 223028 264 223080 270
rect 223028 206 223080 212
rect 224960 264 225012 270
rect 230216 241 230244 439
rect 230308 377 230336 1362
rect 230400 513 230428 1663
rect 230386 504 230442 513
rect 230386 439 230442 448
rect 230294 368 230350 377
rect 230584 338 230612 2518
rect 230676 1970 230704 8758
rect 230938 8664 230994 8673
rect 230848 8628 230900 8634
rect 230938 8599 230940 8608
rect 230848 8570 230900 8576
rect 230992 8599 230994 8608
rect 230940 8570 230992 8576
rect 230860 8514 230888 8570
rect 231044 8514 231072 9862
rect 231492 9376 231544 9382
rect 231492 9318 231544 9324
rect 231308 8832 231360 8838
rect 231308 8774 231360 8780
rect 230860 8486 231072 8514
rect 230756 2576 230808 2582
rect 230756 2518 230808 2524
rect 230768 1970 230796 2518
rect 230860 1970 230888 8486
rect 230940 2440 230992 2446
rect 230940 2382 230992 2388
rect 230952 2106 230980 2382
rect 230940 2100 230992 2106
rect 230940 2042 230992 2048
rect 230664 1964 230716 1970
rect 230664 1906 230716 1912
rect 230756 1964 230808 1970
rect 230756 1906 230808 1912
rect 230848 1964 230900 1970
rect 230848 1906 230900 1912
rect 231320 1426 231348 8774
rect 231504 8498 231532 9318
rect 231872 8974 231900 10134
rect 231964 10130 231992 10270
rect 231952 10124 232004 10130
rect 231952 10066 232004 10072
rect 232320 9580 232372 9586
rect 232320 9522 232372 9528
rect 231950 9480 232006 9489
rect 231950 9415 231952 9424
rect 232004 9415 232006 9424
rect 231952 9386 232004 9392
rect 232332 8974 232360 9522
rect 232792 9081 232820 10474
rect 233516 10124 233568 10130
rect 233516 10066 233568 10072
rect 233422 9480 233478 9489
rect 233422 9415 233424 9424
rect 233476 9415 233478 9424
rect 233424 9386 233476 9392
rect 232778 9072 232834 9081
rect 233528 9058 233556 10066
rect 232778 9007 232780 9016
rect 232832 9007 232834 9016
rect 233436 9030 233556 9058
rect 232780 8978 232832 8984
rect 231860 8968 231912 8974
rect 231860 8910 231912 8916
rect 232044 8968 232096 8974
rect 232044 8910 232096 8916
rect 232320 8968 232372 8974
rect 232320 8910 232372 8916
rect 231674 8664 231730 8673
rect 231674 8599 231676 8608
rect 231728 8599 231730 8608
rect 231768 8628 231820 8634
rect 231676 8570 231728 8576
rect 231768 8570 231820 8576
rect 231492 8492 231544 8498
rect 231492 8434 231544 8440
rect 231400 6384 231452 6390
rect 231400 6326 231452 6332
rect 231308 1420 231360 1426
rect 231308 1362 231360 1368
rect 230294 303 230350 312
rect 230572 332 230624 338
rect 230572 274 230624 280
rect 224960 206 225012 212
rect 230202 232 230258 241
rect 230202 167 230258 176
rect 231412 105 231440 6326
rect 231780 2774 231808 8570
rect 231858 3632 231914 3641
rect 231858 3567 231860 3576
rect 231912 3567 231914 3576
rect 231860 3538 231912 3544
rect 231688 2746 231808 2774
rect 231584 2304 231636 2310
rect 231584 2246 231636 2252
rect 231492 2032 231544 2038
rect 231492 1974 231544 1980
rect 231504 1358 231532 1974
rect 231492 1352 231544 1358
rect 231492 1294 231544 1300
rect 231596 1193 231624 2246
rect 231688 1902 231716 2746
rect 231768 2440 231820 2446
rect 231768 2382 231820 2388
rect 231780 2106 231808 2382
rect 231768 2100 231820 2106
rect 231768 2042 231820 2048
rect 232056 1970 232084 8910
rect 232412 8832 232464 8838
rect 232412 8774 232464 8780
rect 232502 8800 232558 8809
rect 232320 8560 232372 8566
rect 232320 8502 232372 8508
rect 232332 8401 232360 8502
rect 232424 8498 232452 8774
rect 232502 8735 232558 8744
rect 232516 8634 232544 8735
rect 232594 8664 232650 8673
rect 232504 8628 232556 8634
rect 232594 8599 232596 8608
rect 232504 8570 232556 8576
rect 232648 8599 232650 8608
rect 232596 8570 232648 8576
rect 232412 8492 232464 8498
rect 232412 8434 232464 8440
rect 232318 8392 232374 8401
rect 232318 8327 232374 8336
rect 232504 8288 232556 8294
rect 232688 8288 232740 8294
rect 232556 8236 232688 8242
rect 232504 8230 232740 8236
rect 232516 8214 232728 8230
rect 232596 2440 232648 2446
rect 232596 2382 232648 2388
rect 232412 2304 232464 2310
rect 232412 2246 232464 2252
rect 232044 1964 232096 1970
rect 232044 1906 232096 1912
rect 231676 1896 231728 1902
rect 231676 1838 231728 1844
rect 231860 1216 231912 1222
rect 231582 1184 231638 1193
rect 232424 1193 232452 2246
rect 232608 2106 232636 2382
rect 232596 2100 232648 2106
rect 232596 2042 232648 2048
rect 232792 1970 232820 8978
rect 233436 8430 233464 9030
rect 233620 8974 233648 10474
rect 233976 9580 234028 9586
rect 233976 9522 234028 9528
rect 233988 9178 234016 9522
rect 234724 9178 234752 10678
rect 236000 10260 236052 10266
rect 236000 10202 236052 10208
rect 236012 9602 236040 10202
rect 236656 9926 236684 10678
rect 257632 10538 257660 10814
rect 264704 10804 264756 10810
rect 264704 10746 264756 10752
rect 263784 10736 263836 10742
rect 263784 10678 263836 10684
rect 258540 10668 258592 10674
rect 258540 10610 258592 10616
rect 257620 10532 257672 10538
rect 257620 10474 257672 10480
rect 251272 10464 251324 10470
rect 246210 10432 246266 10441
rect 244096 10396 244148 10402
rect 251272 10406 251324 10412
rect 253846 10432 253902 10441
rect 246210 10367 246266 10376
rect 244096 10338 244148 10344
rect 239312 10328 239364 10334
rect 239312 10270 239364 10276
rect 239954 10296 240010 10305
rect 236644 9920 236696 9926
rect 236644 9862 236696 9868
rect 236736 9920 236788 9926
rect 236736 9862 236788 9868
rect 234804 9580 234856 9586
rect 234804 9522 234856 9528
rect 235828 9574 236132 9602
rect 233976 9172 234028 9178
rect 233976 9114 234028 9120
rect 234712 9172 234764 9178
rect 234712 9114 234764 9120
rect 233608 8968 233660 8974
rect 233528 8928 233608 8956
rect 233424 8424 233476 8430
rect 233424 8366 233476 8372
rect 233056 6724 233108 6730
rect 233056 6666 233108 6672
rect 233068 2582 233096 6666
rect 233056 2576 233108 2582
rect 233056 2518 233108 2524
rect 232964 2440 233016 2446
rect 232964 2382 233016 2388
rect 232976 2106 233004 2382
rect 233148 2304 233200 2310
rect 233148 2246 233200 2252
rect 232964 2100 233016 2106
rect 232964 2042 233016 2048
rect 232780 1964 232832 1970
rect 232780 1906 232832 1912
rect 233160 1193 233188 2246
rect 233436 1884 233464 8366
rect 233528 2774 233556 8928
rect 233608 8910 233660 8916
rect 234528 8968 234580 8974
rect 234724 8956 234752 9114
rect 234816 8974 234844 9522
rect 235632 9172 235684 9178
rect 235632 9114 235684 9120
rect 234632 8928 234752 8956
rect 234804 8968 234856 8974
rect 234632 8922 234660 8928
rect 234580 8916 234660 8922
rect 234528 8910 234660 8916
rect 234804 8910 234856 8916
rect 233700 8900 233752 8906
rect 234540 8894 234660 8910
rect 233700 8842 233752 8848
rect 233712 8498 233740 8842
rect 234712 8832 234764 8838
rect 234712 8774 234764 8780
rect 234434 8664 234490 8673
rect 234434 8599 234436 8608
rect 234488 8599 234490 8608
rect 234436 8570 234488 8576
rect 233700 8492 233752 8498
rect 233700 8434 233752 8440
rect 234436 8492 234488 8498
rect 234436 8434 234488 8440
rect 234448 8401 234476 8434
rect 234434 8392 234490 8401
rect 234434 8327 234490 8336
rect 234724 7886 234752 8774
rect 234894 8392 234950 8401
rect 234894 8327 234950 8336
rect 234528 7880 234580 7886
rect 234528 7822 234580 7828
rect 234712 7880 234764 7886
rect 234712 7822 234764 7828
rect 234804 7880 234856 7886
rect 234804 7822 234856 7828
rect 234436 7812 234488 7818
rect 234436 7754 234488 7760
rect 234448 7410 234476 7754
rect 234540 7750 234568 7822
rect 234816 7750 234844 7822
rect 234908 7750 234936 8327
rect 234528 7744 234580 7750
rect 234528 7686 234580 7692
rect 234804 7744 234856 7750
rect 234804 7686 234856 7692
rect 234896 7744 234948 7750
rect 234896 7686 234948 7692
rect 234436 7404 234488 7410
rect 234436 7346 234488 7352
rect 233528 2746 233648 2774
rect 233620 1970 233648 2746
rect 234988 2440 235040 2446
rect 234988 2382 235040 2388
rect 235000 2106 235028 2382
rect 235172 2304 235224 2310
rect 235172 2246 235224 2252
rect 234988 2100 235040 2106
rect 234988 2042 235040 2048
rect 233608 1964 233660 1970
rect 233608 1906 233660 1912
rect 233516 1896 233568 1902
rect 233436 1856 233516 1884
rect 233516 1838 233568 1844
rect 233700 1760 233752 1766
rect 233700 1702 233752 1708
rect 233712 1358 233740 1702
rect 233700 1352 233752 1358
rect 233700 1294 233752 1300
rect 233884 1216 233936 1222
rect 231860 1158 231912 1164
rect 232410 1184 232466 1193
rect 231582 1119 231638 1128
rect 231872 649 231900 1158
rect 232410 1119 232466 1128
rect 233146 1184 233202 1193
rect 233884 1158 233936 1164
rect 234620 1216 234672 1222
rect 235184 1193 235212 2246
rect 235644 1970 235672 9114
rect 235828 8974 235856 9574
rect 235908 9512 235960 9518
rect 235908 9454 235960 9460
rect 235998 9480 236054 9489
rect 235816 8968 235868 8974
rect 235816 8910 235868 8916
rect 235816 8424 235868 8430
rect 235816 8366 235868 8372
rect 235828 7750 235856 8366
rect 235816 7744 235868 7750
rect 235816 7686 235868 7692
rect 235816 2984 235868 2990
rect 235816 2926 235868 2932
rect 235828 2446 235856 2926
rect 235816 2440 235868 2446
rect 235816 2382 235868 2388
rect 235632 1964 235684 1970
rect 235632 1906 235684 1912
rect 235264 1760 235316 1766
rect 235264 1702 235316 1708
rect 235276 1358 235304 1702
rect 235920 1426 235948 9454
rect 235998 9415 236000 9424
rect 236052 9415 236054 9424
rect 236000 9386 236052 9392
rect 235998 8800 236054 8809
rect 235998 8735 236054 8744
rect 236012 8430 236040 8735
rect 236000 8424 236052 8430
rect 236000 8366 236052 8372
rect 236104 1970 236132 9574
rect 236460 9172 236512 9178
rect 236460 9114 236512 9120
rect 236274 8664 236330 8673
rect 236274 8599 236276 8608
rect 236328 8599 236330 8608
rect 236276 8570 236328 8576
rect 236472 8362 236500 9114
rect 236748 9081 236776 9862
rect 237288 9512 237340 9518
rect 237288 9454 237340 9460
rect 236826 9208 236882 9217
rect 236826 9143 236828 9152
rect 236880 9143 236882 9152
rect 236828 9114 236880 9120
rect 236734 9072 236790 9081
rect 236734 9007 236790 9016
rect 236460 8356 236512 8362
rect 236460 8298 236512 8304
rect 236644 7812 236696 7818
rect 236644 7754 236696 7760
rect 236656 7410 236684 7754
rect 237196 7744 237248 7750
rect 237196 7686 237248 7692
rect 237208 7585 237236 7686
rect 237194 7576 237250 7585
rect 237194 7511 237250 7520
rect 236644 7404 236696 7410
rect 236644 7346 236696 7352
rect 236460 6928 236512 6934
rect 236460 6870 236512 6876
rect 236472 5846 236500 6870
rect 236460 5840 236512 5846
rect 236460 5782 236512 5788
rect 237300 5273 237328 9454
rect 238852 9376 238904 9382
rect 238852 9318 238904 9324
rect 237539 9276 237847 9285
rect 237539 9274 237545 9276
rect 237601 9274 237625 9276
rect 237681 9274 237705 9276
rect 237761 9274 237785 9276
rect 237841 9274 237847 9276
rect 237601 9222 237603 9274
rect 237783 9222 237785 9274
rect 237539 9220 237545 9222
rect 237601 9220 237625 9222
rect 237681 9220 237705 9222
rect 237761 9220 237785 9222
rect 237841 9220 237847 9222
rect 237539 9211 237847 9220
rect 238864 8906 238892 9318
rect 238852 8900 238904 8906
rect 238852 8842 238904 8848
rect 239324 8566 239352 10270
rect 239954 10231 240010 10240
rect 240966 10296 241022 10305
rect 240966 10231 241022 10240
rect 241242 10296 241298 10305
rect 241242 10231 241298 10240
rect 242346 10296 242402 10305
rect 242346 10231 242402 10240
rect 242898 10296 242954 10305
rect 242898 10231 242954 10240
rect 243450 10296 243506 10305
rect 243450 10231 243506 10240
rect 239968 9586 239996 10231
rect 240980 9586 241008 10231
rect 239956 9580 240008 9586
rect 239956 9522 240008 9528
rect 240968 9580 241020 9586
rect 240968 9522 241020 9528
rect 240140 9444 240192 9450
rect 240140 9386 240192 9392
rect 239312 8560 239364 8566
rect 239312 8502 239364 8508
rect 237539 8188 237847 8197
rect 237539 8186 237545 8188
rect 237601 8186 237625 8188
rect 237681 8186 237705 8188
rect 237761 8186 237785 8188
rect 237841 8186 237847 8188
rect 237601 8134 237603 8186
rect 237783 8134 237785 8186
rect 237539 8132 237545 8134
rect 237601 8132 237625 8134
rect 237681 8132 237705 8134
rect 237761 8132 237785 8134
rect 237841 8132 237847 8134
rect 237378 8120 237434 8129
rect 237539 8123 237847 8132
rect 237378 8055 237434 8064
rect 237392 7585 237420 8055
rect 240152 7750 240180 9386
rect 241256 8974 241284 10231
rect 242360 9586 242388 10231
rect 242912 9586 242940 10231
rect 242348 9580 242400 9586
rect 242348 9522 242400 9528
rect 242900 9580 242952 9586
rect 242900 9522 242952 9528
rect 243464 9518 243492 10231
rect 242532 9512 242584 9518
rect 242532 9454 242584 9460
rect 243452 9512 243504 9518
rect 243452 9454 243504 9460
rect 241244 8968 241296 8974
rect 241244 8910 241296 8916
rect 241612 8968 241664 8974
rect 241612 8910 241664 8916
rect 240140 7744 240192 7750
rect 240140 7686 240192 7692
rect 237378 7576 237434 7585
rect 237378 7511 237434 7520
rect 237539 7100 237847 7109
rect 237539 7098 237545 7100
rect 237601 7098 237625 7100
rect 237681 7098 237705 7100
rect 237761 7098 237785 7100
rect 237841 7098 237847 7100
rect 237601 7046 237603 7098
rect 237783 7046 237785 7098
rect 237539 7044 237545 7046
rect 237601 7044 237625 7046
rect 237681 7044 237705 7046
rect 237761 7044 237785 7046
rect 237841 7044 237847 7046
rect 237539 7035 237847 7044
rect 241518 7032 241574 7041
rect 241518 6967 241574 6976
rect 241244 6860 241296 6866
rect 241244 6802 241296 6808
rect 241256 6746 241284 6802
rect 241336 6792 241388 6798
rect 241256 6740 241336 6746
rect 241256 6734 241388 6740
rect 239036 6724 239088 6730
rect 241256 6718 241376 6734
rect 239036 6666 239088 6672
rect 237539 6012 237847 6021
rect 237539 6010 237545 6012
rect 237601 6010 237625 6012
rect 237681 6010 237705 6012
rect 237761 6010 237785 6012
rect 237841 6010 237847 6012
rect 237601 5958 237603 6010
rect 237783 5958 237785 6010
rect 237539 5956 237545 5958
rect 237601 5956 237625 5958
rect 237681 5956 237705 5958
rect 237761 5956 237785 5958
rect 237841 5956 237847 5958
rect 237539 5947 237847 5956
rect 239048 5778 239076 6666
rect 239402 6488 239458 6497
rect 239402 6423 239458 6432
rect 239416 6225 239444 6423
rect 241532 6254 241560 6967
rect 241624 6633 241652 8910
rect 242544 7585 242572 9454
rect 244004 9376 244056 9382
rect 244004 9318 244056 9324
rect 242530 7576 242586 7585
rect 242530 7511 242586 7520
rect 241610 6624 241666 6633
rect 241610 6559 241666 6568
rect 241794 6624 241850 6633
rect 241794 6559 241850 6568
rect 241520 6248 241572 6254
rect 239402 6216 239458 6225
rect 241520 6190 241572 6196
rect 239402 6151 239458 6160
rect 239496 6112 239548 6118
rect 239496 6054 239548 6060
rect 239036 5772 239088 5778
rect 239036 5714 239088 5720
rect 238760 5568 238812 5574
rect 238760 5510 238812 5516
rect 237286 5264 237342 5273
rect 237286 5199 237342 5208
rect 237288 5160 237340 5166
rect 237288 5102 237340 5108
rect 237300 4321 237328 5102
rect 237539 4924 237847 4933
rect 237539 4922 237545 4924
rect 237601 4922 237625 4924
rect 237681 4922 237705 4924
rect 237761 4922 237785 4924
rect 237841 4922 237847 4924
rect 237601 4870 237603 4922
rect 237783 4870 237785 4922
rect 237539 4868 237545 4870
rect 237601 4868 237625 4870
rect 237681 4868 237705 4870
rect 237761 4868 237785 4870
rect 237841 4868 237847 4870
rect 237539 4859 237847 4868
rect 237286 4312 237342 4321
rect 237286 4247 237342 4256
rect 237539 3836 237847 3845
rect 237539 3834 237545 3836
rect 237601 3834 237625 3836
rect 237681 3834 237705 3836
rect 237761 3834 237785 3836
rect 237841 3834 237847 3836
rect 237601 3782 237603 3834
rect 237783 3782 237785 3834
rect 237539 3780 237545 3782
rect 237601 3780 237625 3782
rect 237681 3780 237705 3782
rect 237761 3780 237785 3782
rect 237841 3780 237847 3782
rect 237539 3771 237847 3780
rect 238772 3602 238800 5510
rect 239402 3768 239458 3777
rect 239402 3703 239458 3712
rect 238760 3596 238812 3602
rect 238760 3538 238812 3544
rect 236276 3528 236328 3534
rect 236276 3470 236328 3476
rect 236184 2304 236236 2310
rect 236184 2246 236236 2252
rect 236196 2038 236224 2246
rect 236184 2032 236236 2038
rect 236184 1974 236236 1980
rect 236000 1964 236052 1970
rect 236000 1906 236052 1912
rect 236092 1964 236144 1970
rect 236092 1906 236144 1912
rect 235908 1420 235960 1426
rect 235908 1362 235960 1368
rect 236012 1358 236040 1906
rect 235264 1352 235316 1358
rect 235264 1294 235316 1300
rect 236000 1352 236052 1358
rect 236000 1294 236052 1300
rect 235816 1216 235868 1222
rect 234620 1158 234672 1164
rect 235170 1184 235226 1193
rect 233146 1119 233202 1128
rect 233896 649 233924 1158
rect 234632 649 234660 1158
rect 235816 1158 235868 1164
rect 235170 1119 235226 1128
rect 235828 649 235856 1158
rect 231858 640 231914 649
rect 231858 575 231914 584
rect 233882 640 233938 649
rect 233882 575 233938 584
rect 234618 640 234674 649
rect 234618 575 234674 584
rect 235814 640 235870 649
rect 235814 575 235870 584
rect 236288 241 236316 3470
rect 239416 3233 239444 3703
rect 239402 3224 239458 3233
rect 239402 3159 239458 3168
rect 237010 3088 237066 3097
rect 237010 3023 237066 3032
rect 236920 2440 236972 2446
rect 236920 2382 236972 2388
rect 236828 2304 236880 2310
rect 236828 2246 236880 2252
rect 236840 1193 236868 2246
rect 236932 2106 236960 2382
rect 237024 2106 237052 3023
rect 237539 2748 237847 2757
rect 237539 2746 237545 2748
rect 237601 2746 237625 2748
rect 237681 2746 237705 2748
rect 237761 2746 237785 2748
rect 237841 2746 237847 2748
rect 237601 2694 237603 2746
rect 237783 2694 237785 2746
rect 237539 2692 237545 2694
rect 237601 2692 237625 2694
rect 237681 2692 237705 2694
rect 237761 2692 237785 2694
rect 237841 2692 237847 2694
rect 237539 2683 237847 2692
rect 239508 2106 239536 6054
rect 241808 3670 241836 6559
rect 242900 6112 242952 6118
rect 242900 6054 242952 6060
rect 242912 5409 242940 6054
rect 243084 5636 243136 5642
rect 243084 5578 243136 5584
rect 242992 5568 243044 5574
rect 242992 5510 243044 5516
rect 242898 5400 242954 5409
rect 242898 5335 242954 5344
rect 243004 5302 243032 5510
rect 242992 5296 243044 5302
rect 242992 5238 243044 5244
rect 242992 4276 243044 4282
rect 242992 4218 243044 4224
rect 242900 4072 242952 4078
rect 242900 4014 242952 4020
rect 241796 3664 241848 3670
rect 241796 3606 241848 3612
rect 242912 3233 242940 4014
rect 242898 3224 242954 3233
rect 242898 3159 242954 3168
rect 240048 2508 240100 2514
rect 240048 2450 240100 2456
rect 242900 2508 242952 2514
rect 242900 2450 242952 2456
rect 236920 2100 236972 2106
rect 236920 2042 236972 2048
rect 237012 2100 237064 2106
rect 237012 2042 237064 2048
rect 239496 2100 239548 2106
rect 239496 2042 239548 2048
rect 237380 1760 237432 1766
rect 237380 1702 237432 1708
rect 237392 1601 237420 1702
rect 237539 1660 237847 1669
rect 237539 1658 237545 1660
rect 237601 1658 237625 1660
rect 237681 1658 237705 1660
rect 237761 1658 237785 1660
rect 237841 1658 237847 1660
rect 237601 1606 237603 1658
rect 237783 1606 237785 1658
rect 237539 1604 237545 1606
rect 237601 1604 237625 1606
rect 237681 1604 237705 1606
rect 237761 1604 237785 1606
rect 237841 1604 237847 1606
rect 237378 1592 237434 1601
rect 237539 1595 237847 1604
rect 237378 1527 237434 1536
rect 239956 1420 240008 1426
rect 239956 1362 240008 1368
rect 236826 1184 236882 1193
rect 236826 1119 236882 1128
rect 239968 649 239996 1362
rect 240060 1018 240088 2450
rect 241244 1896 241296 1902
rect 241244 1838 241296 1844
rect 242808 1896 242860 1902
rect 242808 1838 242860 1844
rect 240968 1352 241020 1358
rect 240968 1294 241020 1300
rect 241060 1352 241112 1358
rect 241060 1294 241112 1300
rect 240048 1012 240100 1018
rect 240048 954 240100 960
rect 240980 649 241008 1294
rect 239954 640 240010 649
rect 239954 575 240010 584
rect 240966 640 241022 649
rect 240966 575 241022 584
rect 241072 406 241100 1294
rect 241256 649 241284 1838
rect 242820 1465 242848 1838
rect 242806 1456 242862 1465
rect 242806 1391 242862 1400
rect 241980 1352 242032 1358
rect 241980 1294 242032 1300
rect 241992 649 242020 1294
rect 242912 921 242940 2450
rect 242898 912 242954 921
rect 242898 847 242954 856
rect 241242 640 241298 649
rect 241242 575 241298 584
rect 241978 640 242034 649
rect 241978 575 242034 584
rect 243004 406 243032 4218
rect 243096 4185 243124 5578
rect 243082 4176 243138 4185
rect 243082 4111 243138 4120
rect 243636 3732 243688 3738
rect 243636 3674 243688 3680
rect 243360 3052 243412 3058
rect 243360 2994 243412 3000
rect 243372 746 243400 2994
rect 243452 2440 243504 2446
rect 243452 2382 243504 2388
rect 243360 740 243412 746
rect 243360 682 243412 688
rect 243464 649 243492 2382
rect 243648 2310 243676 3674
rect 244016 3602 244044 9318
rect 244108 7177 244136 10338
rect 244186 10296 244242 10305
rect 244186 10231 244242 10240
rect 245014 10296 245070 10305
rect 245014 10231 245070 10240
rect 244200 9518 244228 10231
rect 244188 9512 244240 9518
rect 244188 9454 244240 9460
rect 244924 9172 244976 9178
rect 244924 9114 244976 9120
rect 244094 7168 244150 7177
rect 244094 7103 244150 7112
rect 244648 6316 244700 6322
rect 244648 6258 244700 6264
rect 244200 4010 244504 4026
rect 244188 4004 244516 4010
rect 244240 3998 244464 4004
rect 244188 3946 244240 3952
rect 244464 3946 244516 3952
rect 244280 3936 244332 3942
rect 244332 3884 244504 3890
rect 244280 3878 244504 3884
rect 244292 3862 244504 3878
rect 244372 3664 244424 3670
rect 244372 3606 244424 3612
rect 244004 3596 244056 3602
rect 244004 3538 244056 3544
rect 244004 3460 244056 3466
rect 244004 3402 244056 3408
rect 244280 3460 244332 3466
rect 244280 3402 244332 3408
rect 244016 3126 244044 3402
rect 244004 3120 244056 3126
rect 244004 3062 244056 3068
rect 244292 3058 244320 3402
rect 244384 3194 244412 3606
rect 244372 3188 244424 3194
rect 244372 3130 244424 3136
rect 244280 3052 244332 3058
rect 244280 2994 244332 3000
rect 244372 2984 244424 2990
rect 244372 2926 244424 2932
rect 243912 2644 243964 2650
rect 243912 2586 243964 2592
rect 243728 2440 243780 2446
rect 243728 2382 243780 2388
rect 243636 2304 243688 2310
rect 243636 2246 243688 2252
rect 243636 2100 243688 2106
rect 243636 2042 243688 2048
rect 243544 1556 243596 1562
rect 243544 1498 243596 1504
rect 243556 1329 243584 1498
rect 243542 1320 243598 1329
rect 243542 1255 243598 1264
rect 243648 1057 243676 2042
rect 243634 1048 243690 1057
rect 243634 983 243690 992
rect 243542 912 243598 921
rect 243542 847 243598 856
rect 243556 678 243584 847
rect 243544 672 243596 678
rect 243450 640 243506 649
rect 243544 614 243596 620
rect 243450 575 243506 584
rect 241060 400 241112 406
rect 241060 342 241112 348
rect 242992 400 243044 406
rect 242992 342 243044 348
rect 236274 232 236330 241
rect 243740 202 243768 2382
rect 243820 1352 243872 1358
rect 243820 1294 243872 1300
rect 243832 542 243860 1294
rect 243924 678 243952 2586
rect 244188 2440 244240 2446
rect 244188 2382 244240 2388
rect 243912 672 243964 678
rect 244200 649 244228 2382
rect 244384 1290 244412 2926
rect 244476 2802 244504 3862
rect 244556 3596 244608 3602
rect 244556 3538 244608 3544
rect 244568 2922 244596 3538
rect 244660 3398 244688 6258
rect 244936 5030 244964 9114
rect 245028 8974 245056 10231
rect 245200 9376 245252 9382
rect 245200 9318 245252 9324
rect 245568 9376 245620 9382
rect 245568 9318 245620 9324
rect 245016 8968 245068 8974
rect 245016 8910 245068 8916
rect 245108 8832 245160 8838
rect 245108 8774 245160 8780
rect 245120 6390 245148 8774
rect 245212 8129 245240 9318
rect 245198 8120 245254 8129
rect 245198 8055 245254 8064
rect 245108 6384 245160 6390
rect 245108 6326 245160 6332
rect 245580 5914 245608 9318
rect 246224 8974 246252 10367
rect 246394 10296 246450 10305
rect 246394 10231 246450 10240
rect 247130 10296 247186 10305
rect 247130 10231 247186 10240
rect 247958 10296 248014 10305
rect 247958 10231 248014 10240
rect 248694 10296 248750 10305
rect 248694 10231 248750 10240
rect 249338 10296 249394 10305
rect 249338 10231 249394 10240
rect 250166 10296 250222 10305
rect 250166 10231 250222 10240
rect 251178 10296 251234 10305
rect 251178 10231 251234 10240
rect 246408 9586 246436 10231
rect 246396 9580 246448 9586
rect 246396 9522 246448 9528
rect 246672 9512 246724 9518
rect 246672 9454 246724 9460
rect 246212 8968 246264 8974
rect 246212 8910 246264 8916
rect 246304 8832 246356 8838
rect 246304 8774 246356 8780
rect 245568 5908 245620 5914
rect 245568 5850 245620 5856
rect 245568 5772 245620 5778
rect 245568 5714 245620 5720
rect 245016 5296 245068 5302
rect 245016 5238 245068 5244
rect 244924 5024 244976 5030
rect 244924 4966 244976 4972
rect 244924 4616 244976 4622
rect 244924 4558 244976 4564
rect 244648 3392 244700 3398
rect 244648 3334 244700 3340
rect 244832 3392 244884 3398
rect 244832 3334 244884 3340
rect 244844 3126 244872 3334
rect 244936 3194 244964 4558
rect 245028 4146 245056 5238
rect 245108 5024 245160 5030
rect 245108 4966 245160 4972
rect 245016 4140 245068 4146
rect 245016 4082 245068 4088
rect 245016 3460 245068 3466
rect 245016 3402 245068 3408
rect 245028 3194 245056 3402
rect 244924 3188 244976 3194
rect 244924 3130 244976 3136
rect 245016 3188 245068 3194
rect 245016 3130 245068 3136
rect 245120 3126 245148 4966
rect 245580 4826 245608 5714
rect 246212 5364 246264 5370
rect 246212 5306 246264 5312
rect 246224 5273 246252 5306
rect 246210 5264 246266 5273
rect 246210 5199 246266 5208
rect 246316 5137 246344 8774
rect 246684 7721 246712 9454
rect 247144 8974 247172 10231
rect 247972 9586 248000 10231
rect 247960 9580 248012 9586
rect 247960 9522 248012 9528
rect 248708 8974 248736 10231
rect 249352 9586 249380 10231
rect 249340 9580 249392 9586
rect 249340 9522 249392 9528
rect 249616 9512 249668 9518
rect 249616 9454 249668 9460
rect 249708 9512 249760 9518
rect 249708 9454 249760 9460
rect 247132 8968 247184 8974
rect 247132 8910 247184 8916
rect 247408 8968 247460 8974
rect 247408 8910 247460 8916
rect 248696 8968 248748 8974
rect 248696 8910 248748 8916
rect 246948 8900 247000 8906
rect 246948 8842 247000 8848
rect 246960 8129 246988 8842
rect 247040 8832 247092 8838
rect 247040 8774 247092 8780
rect 246946 8120 247002 8129
rect 246946 8055 247002 8064
rect 246670 7712 246726 7721
rect 246670 7647 246726 7656
rect 247052 5778 247080 8774
rect 247420 6118 247448 8910
rect 249064 8900 249116 8906
rect 249064 8842 249116 8848
rect 248880 8628 248932 8634
rect 248880 8570 248932 8576
rect 248972 8628 249024 8634
rect 248972 8570 249024 8576
rect 248892 7750 248920 8570
rect 248880 7744 248932 7750
rect 248880 7686 248932 7692
rect 248420 7200 248472 7206
rect 248420 7142 248472 7148
rect 248432 6798 248460 7142
rect 248984 7041 249012 8570
rect 249076 8294 249104 8842
rect 249064 8288 249116 8294
rect 249064 8230 249116 8236
rect 249628 7478 249656 9454
rect 249720 9178 249748 9454
rect 249708 9172 249760 9178
rect 249708 9114 249760 9120
rect 249800 9172 249852 9178
rect 249800 9114 249852 9120
rect 249812 8090 249840 9114
rect 250180 8974 250208 10231
rect 251192 8974 251220 10231
rect 250168 8968 250220 8974
rect 250168 8910 250220 8916
rect 251180 8968 251232 8974
rect 251180 8910 251232 8916
rect 250260 8832 250312 8838
rect 250260 8774 250312 8780
rect 250352 8832 250404 8838
rect 250352 8774 250404 8780
rect 250272 8498 250300 8774
rect 250260 8492 250312 8498
rect 250260 8434 250312 8440
rect 249800 8084 249852 8090
rect 249800 8026 249852 8032
rect 250166 7984 250222 7993
rect 250166 7919 250222 7928
rect 249800 7744 249852 7750
rect 249800 7686 249852 7692
rect 249616 7472 249668 7478
rect 249616 7414 249668 7420
rect 248970 7032 249026 7041
rect 248970 6967 249026 6976
rect 248420 6792 248472 6798
rect 248420 6734 248472 6740
rect 248512 6792 248564 6798
rect 248512 6734 248564 6740
rect 249340 6792 249392 6798
rect 249812 6769 249840 7686
rect 249984 7336 250036 7342
rect 249984 7278 250036 7284
rect 249996 7002 250024 7278
rect 249984 6996 250036 7002
rect 249984 6938 250036 6944
rect 250076 6860 250128 6866
rect 250076 6802 250128 6808
rect 249340 6734 249392 6740
rect 249798 6760 249854 6769
rect 248326 6488 248382 6497
rect 248326 6423 248328 6432
rect 248380 6423 248382 6432
rect 248328 6394 248380 6400
rect 248236 6316 248288 6322
rect 248236 6258 248288 6264
rect 248328 6316 248380 6322
rect 248328 6258 248380 6264
rect 248144 6180 248196 6186
rect 248144 6122 248196 6128
rect 247408 6112 247460 6118
rect 247408 6054 247460 6060
rect 248052 5908 248104 5914
rect 248052 5850 248104 5856
rect 247684 5840 247736 5846
rect 247684 5782 247736 5788
rect 247040 5772 247092 5778
rect 247040 5714 247092 5720
rect 246856 5704 246908 5710
rect 246856 5646 246908 5652
rect 247406 5672 247462 5681
rect 246580 5296 246632 5302
rect 246580 5238 246632 5244
rect 246302 5128 246358 5137
rect 246302 5063 246358 5072
rect 245568 4820 245620 4826
rect 245568 4762 245620 4768
rect 246488 4820 246540 4826
rect 246488 4762 246540 4768
rect 245934 4720 245990 4729
rect 245934 4655 245990 4664
rect 245568 4616 245620 4622
rect 245568 4558 245620 4564
rect 245384 4480 245436 4486
rect 245384 4422 245436 4428
rect 244832 3120 244884 3126
rect 244832 3062 244884 3068
rect 245108 3120 245160 3126
rect 245108 3062 245160 3068
rect 244556 2916 244608 2922
rect 244556 2858 244608 2864
rect 244648 2916 244700 2922
rect 244648 2858 244700 2864
rect 244660 2802 244688 2858
rect 244476 2774 244688 2802
rect 245016 2440 245068 2446
rect 245016 2382 245068 2388
rect 245028 2281 245056 2382
rect 245014 2272 245070 2281
rect 245014 2207 245070 2216
rect 245396 2038 245424 4422
rect 245580 3398 245608 4558
rect 245660 3732 245712 3738
rect 245660 3674 245712 3680
rect 245568 3392 245620 3398
rect 245474 3360 245530 3369
rect 245568 3334 245620 3340
rect 245474 3295 245530 3304
rect 245488 2650 245516 3295
rect 245672 2854 245700 3674
rect 245660 2848 245712 2854
rect 245660 2790 245712 2796
rect 245476 2644 245528 2650
rect 245476 2586 245528 2592
rect 245384 2032 245436 2038
rect 245384 1974 245436 1980
rect 245948 1902 245976 4655
rect 246304 4548 246356 4554
rect 246304 4490 246356 4496
rect 246316 2854 246344 4490
rect 246500 3738 246528 4762
rect 246592 4554 246620 5238
rect 246672 5228 246724 5234
rect 246672 5170 246724 5176
rect 246580 4548 246632 4554
rect 246580 4490 246632 4496
rect 246488 3732 246540 3738
rect 246488 3674 246540 3680
rect 246304 2848 246356 2854
rect 246304 2790 246356 2796
rect 246500 2774 246528 3674
rect 246592 3466 246620 4490
rect 246684 3738 246712 5170
rect 246868 5166 246896 5646
rect 247040 5636 247092 5642
rect 247406 5607 247462 5616
rect 247040 5578 247092 5584
rect 247052 5386 247080 5578
rect 246960 5358 247080 5386
rect 246960 5302 246988 5358
rect 246948 5296 247000 5302
rect 246948 5238 247000 5244
rect 247040 5228 247092 5234
rect 247224 5228 247276 5234
rect 247092 5188 247172 5216
rect 247040 5170 247092 5176
rect 246856 5160 246908 5166
rect 246856 5102 246908 5108
rect 246868 4622 246896 5102
rect 247040 5092 247092 5098
rect 247040 5034 247092 5040
rect 246948 5024 247000 5030
rect 246948 4966 247000 4972
rect 246960 4826 246988 4966
rect 246948 4820 247000 4826
rect 246948 4762 247000 4768
rect 246856 4616 246908 4622
rect 246856 4558 246908 4564
rect 246948 4616 247000 4622
rect 246948 4558 247000 4564
rect 246868 4214 246896 4558
rect 246856 4208 246908 4214
rect 246856 4150 246908 4156
rect 246672 3732 246724 3738
rect 246672 3674 246724 3680
rect 246868 3602 246896 4150
rect 246960 3618 246988 4558
rect 247052 4282 247080 5034
rect 247144 4622 247172 5188
rect 247224 5170 247276 5176
rect 247132 4616 247184 4622
rect 247132 4558 247184 4564
rect 247132 4480 247184 4486
rect 247132 4422 247184 4428
rect 247040 4276 247092 4282
rect 247040 4218 247092 4224
rect 247144 4146 247172 4422
rect 247236 4146 247264 5170
rect 247316 4548 247368 4554
rect 247316 4490 247368 4496
rect 247132 4140 247184 4146
rect 247132 4082 247184 4088
rect 247224 4140 247276 4146
rect 247224 4082 247276 4088
rect 246856 3596 246908 3602
rect 246856 3538 246908 3544
rect 246960 3590 247172 3618
rect 247328 3602 247356 4490
rect 246960 3534 246988 3590
rect 246948 3528 247000 3534
rect 246948 3470 247000 3476
rect 247040 3528 247092 3534
rect 247040 3470 247092 3476
rect 246580 3460 246632 3466
rect 246580 3402 246632 3408
rect 246856 2984 246908 2990
rect 246854 2952 246856 2961
rect 246908 2952 246910 2961
rect 246854 2887 246910 2896
rect 246500 2746 246620 2774
rect 246304 2372 246356 2378
rect 246304 2314 246356 2320
rect 244832 1896 244884 1902
rect 244832 1838 244884 1844
rect 245936 1896 245988 1902
rect 245936 1838 245988 1844
rect 244372 1284 244424 1290
rect 244372 1226 244424 1232
rect 243912 614 243964 620
rect 244186 640 244242 649
rect 244186 575 244242 584
rect 243820 536 243872 542
rect 243820 478 243872 484
rect 244844 270 244872 1838
rect 245752 1828 245804 1834
rect 245752 1770 245804 1776
rect 245764 1465 245792 1770
rect 245750 1456 245806 1465
rect 245750 1391 245806 1400
rect 246028 1352 246080 1358
rect 246080 1300 246252 1306
rect 246028 1294 246252 1300
rect 246040 1290 246252 1294
rect 244924 1284 244976 1290
rect 246040 1284 246264 1290
rect 246040 1278 246212 1284
rect 244924 1226 244976 1232
rect 246212 1226 246264 1232
rect 244936 649 244964 1226
rect 246316 1222 246344 2314
rect 246592 1562 246620 2746
rect 246856 2576 246908 2582
rect 246856 2518 246908 2524
rect 246672 1896 246724 1902
rect 246672 1838 246724 1844
rect 246684 1737 246712 1838
rect 246670 1728 246726 1737
rect 246670 1663 246726 1672
rect 246580 1556 246632 1562
rect 246580 1498 246632 1504
rect 246396 1352 246448 1358
rect 246396 1294 246448 1300
rect 246304 1216 246356 1222
rect 246304 1158 246356 1164
rect 246408 950 246436 1294
rect 246396 944 246448 950
rect 246396 886 246448 892
rect 244922 640 244978 649
rect 244922 575 244978 584
rect 246868 542 246896 2518
rect 246946 1592 247002 1601
rect 246946 1527 247002 1536
rect 246960 1057 246988 1527
rect 246946 1048 247002 1057
rect 246946 983 247002 992
rect 247052 649 247080 3470
rect 247144 1170 247172 3590
rect 247316 3596 247368 3602
rect 247316 3538 247368 3544
rect 247224 3460 247276 3466
rect 247224 3402 247276 3408
rect 247236 1358 247264 3402
rect 247420 2990 247448 5607
rect 247696 5302 247724 5782
rect 247960 5772 248012 5778
rect 247960 5714 248012 5720
rect 247776 5636 247828 5642
rect 247776 5578 247828 5584
rect 247684 5296 247736 5302
rect 247684 5238 247736 5244
rect 247500 4752 247552 4758
rect 247500 4694 247552 4700
rect 247408 2984 247460 2990
rect 247408 2926 247460 2932
rect 247406 2272 247462 2281
rect 247406 2207 247462 2216
rect 247420 1970 247448 2207
rect 247408 1964 247460 1970
rect 247408 1906 247460 1912
rect 247512 1902 247540 4694
rect 247696 4690 247724 5238
rect 247684 4684 247736 4690
rect 247684 4626 247736 4632
rect 247788 4622 247816 5578
rect 247868 5228 247920 5234
rect 247972 5216 248000 5714
rect 247920 5188 248000 5216
rect 247868 5170 247920 5176
rect 248064 4826 248092 5850
rect 248156 5370 248184 6122
rect 248248 5914 248276 6258
rect 248236 5908 248288 5914
rect 248236 5850 248288 5856
rect 248340 5778 248368 6258
rect 248524 5846 248552 6734
rect 248880 6656 248932 6662
rect 248880 6598 248932 6604
rect 249248 6656 249300 6662
rect 249248 6598 249300 6604
rect 248696 6248 248748 6254
rect 248696 6190 248748 6196
rect 248604 6112 248656 6118
rect 248604 6054 248656 6060
rect 248420 5840 248472 5846
rect 248420 5782 248472 5788
rect 248512 5840 248564 5846
rect 248512 5782 248564 5788
rect 248328 5772 248380 5778
rect 248328 5714 248380 5720
rect 248432 5710 248460 5782
rect 248236 5704 248288 5710
rect 248236 5646 248288 5652
rect 248420 5704 248472 5710
rect 248420 5646 248472 5652
rect 248144 5364 248196 5370
rect 248144 5306 248196 5312
rect 248052 4820 248104 4826
rect 248052 4762 248104 4768
rect 248248 4758 248276 5646
rect 248512 5568 248564 5574
rect 248512 5510 248564 5516
rect 248326 5264 248382 5273
rect 248326 5199 248382 5208
rect 248340 5098 248368 5199
rect 248328 5092 248380 5098
rect 248328 5034 248380 5040
rect 248236 4752 248288 4758
rect 248236 4694 248288 4700
rect 247776 4616 247828 4622
rect 247776 4558 247828 4564
rect 248248 4554 248276 4694
rect 248236 4548 248288 4554
rect 248236 4490 248288 4496
rect 247592 4140 247644 4146
rect 247592 4082 247644 4088
rect 247604 3738 247632 4082
rect 248420 4072 248472 4078
rect 248420 4014 248472 4020
rect 247592 3732 247644 3738
rect 247644 3692 247724 3720
rect 247592 3674 247644 3680
rect 247500 1896 247552 1902
rect 247500 1838 247552 1844
rect 247696 1426 247724 3692
rect 248142 3496 248198 3505
rect 248142 3431 248144 3440
rect 248196 3431 248198 3440
rect 248144 3402 248196 3408
rect 248432 3398 248460 4014
rect 248420 3392 248472 3398
rect 248420 3334 248472 3340
rect 248420 3052 248472 3058
rect 248420 2994 248472 3000
rect 248432 2417 248460 2994
rect 248524 2774 248552 5510
rect 248616 3126 248644 6054
rect 248708 5234 248736 6190
rect 248788 6112 248840 6118
rect 248788 6054 248840 6060
rect 248800 5914 248828 6054
rect 248788 5908 248840 5914
rect 248788 5850 248840 5856
rect 248696 5228 248748 5234
rect 248696 5170 248748 5176
rect 248800 5030 248828 5850
rect 248892 5302 248920 6598
rect 249156 6316 249208 6322
rect 249156 6258 249208 6264
rect 249064 6112 249116 6118
rect 249064 6054 249116 6060
rect 248880 5296 248932 5302
rect 248880 5238 248932 5244
rect 248788 5024 248840 5030
rect 248788 4966 248840 4972
rect 249076 4690 249104 6054
rect 249168 5710 249196 6258
rect 249156 5704 249208 5710
rect 249156 5646 249208 5652
rect 249168 5166 249196 5646
rect 249156 5160 249208 5166
rect 249156 5102 249208 5108
rect 249064 4684 249116 4690
rect 249064 4626 249116 4632
rect 248880 4616 248932 4622
rect 248880 4558 248932 4564
rect 248892 4321 248920 4558
rect 248878 4312 248934 4321
rect 248878 4247 248934 4256
rect 249062 4312 249118 4321
rect 249062 4247 249118 4256
rect 248786 4176 248842 4185
rect 248786 4111 248842 4120
rect 248696 4072 248748 4078
rect 248696 4014 248748 4020
rect 248708 3913 248736 4014
rect 248694 3904 248750 3913
rect 248694 3839 248750 3848
rect 248604 3120 248656 3126
rect 248604 3062 248656 3068
rect 248696 3052 248748 3058
rect 248800 3040 248828 4111
rect 249076 3097 249104 4247
rect 249260 3602 249288 6598
rect 249352 6458 249380 6734
rect 249798 6695 249854 6704
rect 249340 6452 249392 6458
rect 249340 6394 249392 6400
rect 249340 6248 249392 6254
rect 249340 6190 249392 6196
rect 249352 5642 249380 6190
rect 249892 6112 249944 6118
rect 249812 6072 249892 6100
rect 249432 5840 249484 5846
rect 249432 5782 249484 5788
rect 249340 5636 249392 5642
rect 249340 5578 249392 5584
rect 249444 4078 249472 5782
rect 249812 5778 249840 6072
rect 249892 6054 249944 6060
rect 249800 5772 249852 5778
rect 249800 5714 249852 5720
rect 249984 5772 250036 5778
rect 249984 5714 250036 5720
rect 249996 5574 250024 5714
rect 249984 5568 250036 5574
rect 249984 5510 250036 5516
rect 249708 4480 249760 4486
rect 249708 4422 249760 4428
rect 249432 4072 249484 4078
rect 249432 4014 249484 4020
rect 249248 3596 249300 3602
rect 249248 3538 249300 3544
rect 249616 3392 249668 3398
rect 249616 3334 249668 3340
rect 248748 3012 248828 3040
rect 249062 3088 249118 3097
rect 249062 3023 249118 3032
rect 248696 2994 248748 3000
rect 249628 2825 249656 3334
rect 249614 2816 249670 2825
rect 248524 2746 248644 2774
rect 249614 2751 249670 2760
rect 248512 2576 248564 2582
rect 248512 2518 248564 2524
rect 248418 2408 248474 2417
rect 248418 2343 248474 2352
rect 247684 1420 247736 1426
rect 247684 1362 247736 1368
rect 247224 1352 247276 1358
rect 247592 1352 247644 1358
rect 247224 1294 247276 1300
rect 247328 1312 247592 1340
rect 247328 1170 247356 1312
rect 247592 1294 247644 1300
rect 247144 1142 247356 1170
rect 248052 1216 248104 1222
rect 248052 1158 248104 1164
rect 248420 1216 248472 1222
rect 248420 1158 248472 1164
rect 247038 640 247094 649
rect 247038 575 247094 584
rect 246856 536 246908 542
rect 246856 478 246908 484
rect 248064 338 248092 1158
rect 248432 649 248460 1158
rect 248524 785 248552 2518
rect 248616 2514 248644 2746
rect 248880 2644 248932 2650
rect 248880 2586 248932 2592
rect 248604 2508 248656 2514
rect 248604 2450 248656 2456
rect 248788 2440 248840 2446
rect 248788 2382 248840 2388
rect 248800 882 248828 2382
rect 248892 2106 248920 2586
rect 249720 2553 249748 4422
rect 250088 3058 250116 6802
rect 250180 4321 250208 7919
rect 250364 5545 250392 8774
rect 251284 8294 251312 10406
rect 253846 10367 253902 10376
rect 251546 10296 251602 10305
rect 251546 10231 251602 10240
rect 252282 10296 252338 10305
rect 252282 10231 252338 10240
rect 253754 10296 253810 10305
rect 253754 10231 253810 10240
rect 251560 9586 251588 10231
rect 251548 9580 251600 9586
rect 251548 9522 251600 9528
rect 252296 8974 252324 10231
rect 253768 8974 253796 10231
rect 253860 9586 253888 10367
rect 255042 10296 255098 10305
rect 255042 10231 255098 10240
rect 255318 10296 255374 10305
rect 255318 10231 255374 10240
rect 256422 10296 256478 10305
rect 256422 10231 256478 10240
rect 256698 10296 256754 10305
rect 256698 10231 256754 10240
rect 257710 10296 257766 10305
rect 257710 10231 257766 10240
rect 258262 10296 258318 10305
rect 258262 10231 258318 10240
rect 253848 9580 253900 9586
rect 253848 9522 253900 9528
rect 254124 9512 254176 9518
rect 254124 9454 254176 9460
rect 252284 8968 252336 8974
rect 252284 8910 252336 8916
rect 253756 8968 253808 8974
rect 253756 8910 253808 8916
rect 251548 8832 251600 8838
rect 251548 8774 251600 8780
rect 251560 8634 251588 8774
rect 251548 8628 251600 8634
rect 251548 8570 251600 8576
rect 251272 8288 251324 8294
rect 251272 8230 251324 8236
rect 254136 7993 254164 9454
rect 254676 9172 254728 9178
rect 254676 9114 254728 9120
rect 254688 9042 254716 9114
rect 254768 9104 254820 9110
rect 254952 9104 255004 9110
rect 254820 9052 254952 9058
rect 254768 9046 255004 9052
rect 254676 9036 254728 9042
rect 254780 9030 254992 9046
rect 255056 9042 255084 10231
rect 255228 9648 255280 9654
rect 255228 9590 255280 9596
rect 255044 9036 255096 9042
rect 254676 8978 254728 8984
rect 255044 8978 255096 8984
rect 254122 7984 254178 7993
rect 254122 7919 254178 7928
rect 253112 7880 253164 7886
rect 253112 7822 253164 7828
rect 253124 7478 253152 7822
rect 252100 7472 252152 7478
rect 252098 7440 252100 7449
rect 253112 7472 253164 7478
rect 252152 7440 252154 7449
rect 251456 7404 251508 7410
rect 253112 7414 253164 7420
rect 252098 7375 252154 7384
rect 252836 7404 252888 7410
rect 251456 7346 251508 7352
rect 252836 7346 252888 7352
rect 253204 7404 253256 7410
rect 253204 7346 253256 7352
rect 251180 7336 251232 7342
rect 251178 7304 251180 7313
rect 251232 7304 251234 7313
rect 251178 7239 251234 7248
rect 251468 6798 251496 7346
rect 251640 7268 251692 7274
rect 251640 7210 251692 7216
rect 251652 6866 251680 7210
rect 252848 7206 252876 7346
rect 252836 7200 252888 7206
rect 252836 7142 252888 7148
rect 251640 6860 251692 6866
rect 251640 6802 251692 6808
rect 253216 6798 253244 7346
rect 251364 6792 251416 6798
rect 251364 6734 251416 6740
rect 251456 6792 251508 6798
rect 251456 6734 251508 6740
rect 253020 6792 253072 6798
rect 253020 6734 253072 6740
rect 253204 6792 253256 6798
rect 253204 6734 253256 6740
rect 251376 6322 251404 6734
rect 251640 6656 251692 6662
rect 251640 6598 251692 6604
rect 251732 6656 251784 6662
rect 251732 6598 251784 6604
rect 251652 6361 251680 6598
rect 251638 6352 251694 6361
rect 251364 6316 251416 6322
rect 251638 6287 251694 6296
rect 251364 6258 251416 6264
rect 251456 6112 251508 6118
rect 251456 6054 251508 6060
rect 250628 5840 250680 5846
rect 250628 5782 250680 5788
rect 250996 5840 251048 5846
rect 250996 5782 251048 5788
rect 250536 5704 250588 5710
rect 250640 5692 250668 5782
rect 250588 5664 250668 5692
rect 250720 5704 250772 5710
rect 250536 5646 250588 5652
rect 250720 5646 250772 5652
rect 250444 5568 250496 5574
rect 250350 5536 250406 5545
rect 250732 5556 250760 5646
rect 250496 5528 250760 5556
rect 250444 5510 250496 5516
rect 250350 5471 250406 5480
rect 250166 4312 250222 4321
rect 250166 4247 250222 4256
rect 251008 4146 251036 5782
rect 251272 5636 251324 5642
rect 251272 5578 251324 5584
rect 251284 5098 251312 5578
rect 251272 5092 251324 5098
rect 251272 5034 251324 5040
rect 251180 5024 251232 5030
rect 251180 4966 251232 4972
rect 251086 4856 251142 4865
rect 251192 4826 251220 4966
rect 251086 4791 251142 4800
rect 251180 4820 251232 4826
rect 250996 4140 251048 4146
rect 250996 4082 251048 4088
rect 250812 4072 250864 4078
rect 250812 4014 250864 4020
rect 250076 3052 250128 3058
rect 250076 2994 250128 3000
rect 250536 2984 250588 2990
rect 250534 2952 250536 2961
rect 250588 2952 250590 2961
rect 250534 2887 250590 2896
rect 249706 2544 249762 2553
rect 249706 2479 249762 2488
rect 248880 2100 248932 2106
rect 248880 2042 248932 2048
rect 250824 2009 250852 4014
rect 250996 3528 251048 3534
rect 250996 3470 251048 3476
rect 251008 3097 251036 3470
rect 250994 3088 251050 3097
rect 250994 3023 251050 3032
rect 251100 2689 251128 4791
rect 251180 4762 251232 4768
rect 251272 4548 251324 4554
rect 251272 4490 251324 4496
rect 251364 4548 251416 4554
rect 251364 4490 251416 4496
rect 251284 4214 251312 4490
rect 251272 4208 251324 4214
rect 251272 4150 251324 4156
rect 251376 4078 251404 4490
rect 251364 4072 251416 4078
rect 251364 4014 251416 4020
rect 251376 3534 251404 4014
rect 251364 3528 251416 3534
rect 251364 3470 251416 3476
rect 251180 2984 251232 2990
rect 251180 2926 251232 2932
rect 251086 2680 251142 2689
rect 251086 2615 251142 2624
rect 250810 2000 250866 2009
rect 250810 1935 250866 1944
rect 250536 1896 250588 1902
rect 250536 1838 250588 1844
rect 249800 1828 249852 1834
rect 249800 1770 249852 1776
rect 249812 1465 249840 1770
rect 250548 1494 250576 1838
rect 250536 1488 250588 1494
rect 249798 1456 249854 1465
rect 250536 1430 250588 1436
rect 249798 1391 249854 1400
rect 248972 1284 249024 1290
rect 248972 1226 249024 1232
rect 248984 950 249012 1226
rect 251192 1222 251220 2926
rect 251468 2514 251496 6054
rect 251744 5914 251772 6598
rect 251732 5908 251784 5914
rect 251732 5850 251784 5856
rect 251744 5302 251772 5850
rect 251732 5296 251784 5302
rect 251732 5238 251784 5244
rect 252652 5160 252704 5166
rect 252652 5102 252704 5108
rect 251732 5024 251784 5030
rect 251732 4966 251784 4972
rect 251640 4684 251692 4690
rect 251640 4626 251692 4632
rect 251652 3738 251680 4626
rect 251640 3732 251692 3738
rect 251640 3674 251692 3680
rect 251652 3602 251680 3674
rect 251640 3596 251692 3602
rect 251640 3538 251692 3544
rect 251456 2508 251508 2514
rect 251456 2450 251508 2456
rect 251272 1896 251324 1902
rect 251270 1864 251272 1873
rect 251364 1896 251416 1902
rect 251324 1864 251326 1873
rect 251364 1838 251416 1844
rect 251270 1799 251326 1808
rect 251376 1601 251404 1838
rect 251362 1592 251418 1601
rect 251362 1527 251418 1536
rect 251548 1352 251600 1358
rect 251548 1294 251600 1300
rect 251180 1216 251232 1222
rect 251180 1158 251232 1164
rect 249064 1012 249116 1018
rect 249064 954 249116 960
rect 250076 1012 250128 1018
rect 250076 954 250128 960
rect 248972 944 249024 950
rect 248972 886 249024 892
rect 248788 876 248840 882
rect 248788 818 248840 824
rect 248510 776 248566 785
rect 248510 711 248566 720
rect 249076 678 249104 954
rect 249064 672 249116 678
rect 248418 640 248474 649
rect 250088 649 250116 954
rect 249064 614 249116 620
rect 250074 640 250130 649
rect 248418 575 248474 584
rect 250074 575 250130 584
rect 251560 474 251588 1294
rect 251744 950 251772 4966
rect 252468 4820 252520 4826
rect 252468 4762 252520 4768
rect 252480 4026 252508 4762
rect 252560 4548 252612 4554
rect 252560 4490 252612 4496
rect 252572 4214 252600 4490
rect 252664 4321 252692 5102
rect 253032 4826 253060 6734
rect 253112 6724 253164 6730
rect 253112 6666 253164 6672
rect 253124 6458 253152 6666
rect 253112 6452 253164 6458
rect 253112 6394 253164 6400
rect 253216 6322 253244 6734
rect 253848 6656 253900 6662
rect 253848 6598 253900 6604
rect 253204 6316 253256 6322
rect 253204 6258 253256 6264
rect 253216 4826 253244 6258
rect 253478 6216 253534 6225
rect 253478 6151 253534 6160
rect 253296 5772 253348 5778
rect 253296 5714 253348 5720
rect 253020 4820 253072 4826
rect 253020 4762 253072 4768
rect 253204 4820 253256 4826
rect 253204 4762 253256 4768
rect 253112 4752 253164 4758
rect 253112 4694 253164 4700
rect 253020 4684 253072 4690
rect 253020 4626 253072 4632
rect 252836 4616 252888 4622
rect 252836 4558 252888 4564
rect 252744 4480 252796 4486
rect 252744 4422 252796 4428
rect 252650 4312 252706 4321
rect 252650 4247 252706 4256
rect 252560 4208 252612 4214
rect 252560 4150 252612 4156
rect 252652 4140 252704 4146
rect 252652 4082 252704 4088
rect 252480 3998 252600 4026
rect 252572 3738 252600 3998
rect 252560 3732 252612 3738
rect 252560 3674 252612 3680
rect 252664 3466 252692 4082
rect 252652 3460 252704 3466
rect 252652 3402 252704 3408
rect 252652 2440 252704 2446
rect 252652 2382 252704 2388
rect 252376 2372 252428 2378
rect 252376 2314 252428 2320
rect 252388 2038 252416 2314
rect 252376 2032 252428 2038
rect 252376 1974 252428 1980
rect 252560 1760 252612 1766
rect 252560 1702 252612 1708
rect 252572 1601 252600 1702
rect 252558 1592 252614 1601
rect 252558 1527 252614 1536
rect 252664 1465 252692 2382
rect 252650 1456 252706 1465
rect 252650 1391 252706 1400
rect 252756 1358 252784 4422
rect 252848 3942 252876 4558
rect 252928 4548 252980 4554
rect 252928 4490 252980 4496
rect 252940 4146 252968 4490
rect 252928 4140 252980 4146
rect 252928 4082 252980 4088
rect 253032 4078 253060 4626
rect 253020 4072 253072 4078
rect 253020 4014 253072 4020
rect 252836 3936 252888 3942
rect 252836 3878 252888 3884
rect 252848 3738 252876 3878
rect 252836 3732 252888 3738
rect 252836 3674 252888 3680
rect 253124 2774 253152 4694
rect 253308 3670 253336 5714
rect 253296 3664 253348 3670
rect 253296 3606 253348 3612
rect 252940 2746 253152 2774
rect 252744 1352 252796 1358
rect 252744 1294 252796 1300
rect 252836 1352 252888 1358
rect 252836 1294 252888 1300
rect 252848 1018 252876 1294
rect 252940 1018 252968 2746
rect 253492 2514 253520 6151
rect 253860 5710 253888 6598
rect 255240 6390 255268 9590
rect 255332 9586 255360 10231
rect 255320 9580 255372 9586
rect 255320 9522 255372 9528
rect 256436 9042 256464 10231
rect 256424 9036 256476 9042
rect 256424 8978 256476 8984
rect 255320 8968 255372 8974
rect 255320 8910 255372 8916
rect 255332 7954 255360 8910
rect 256712 8498 256740 10231
rect 256884 9512 256936 9518
rect 256884 9454 256936 9460
rect 256792 8968 256844 8974
rect 256792 8910 256844 8916
rect 256700 8492 256752 8498
rect 256700 8434 256752 8440
rect 255320 7948 255372 7954
rect 255320 7890 255372 7896
rect 256804 7546 256832 8910
rect 256896 8022 256924 9454
rect 257724 9042 257752 10231
rect 257896 9580 257948 9586
rect 257896 9522 257948 9528
rect 257988 9580 258040 9586
rect 257988 9522 258040 9528
rect 257908 9042 257936 9522
rect 257712 9036 257764 9042
rect 257712 8978 257764 8984
rect 257896 9036 257948 9042
rect 257896 8978 257948 8984
rect 256976 8424 257028 8430
rect 256976 8366 257028 8372
rect 256884 8016 256936 8022
rect 256884 7958 256936 7964
rect 256988 7818 257016 8366
rect 256976 7812 257028 7818
rect 256976 7754 257028 7760
rect 256792 7540 256844 7546
rect 256792 7482 256844 7488
rect 256700 6792 256752 6798
rect 256700 6734 256752 6740
rect 255596 6656 255648 6662
rect 255596 6598 255648 6604
rect 255780 6656 255832 6662
rect 255780 6598 255832 6604
rect 256608 6656 256660 6662
rect 256608 6598 256660 6604
rect 255608 6458 255636 6598
rect 255320 6452 255372 6458
rect 255320 6394 255372 6400
rect 255596 6452 255648 6458
rect 255596 6394 255648 6400
rect 255228 6384 255280 6390
rect 255228 6326 255280 6332
rect 254032 6316 254084 6322
rect 254032 6258 254084 6264
rect 253848 5704 253900 5710
rect 253848 5646 253900 5652
rect 253848 5160 253900 5166
rect 253848 5102 253900 5108
rect 253860 4214 253888 5102
rect 253940 5024 253992 5030
rect 253940 4966 253992 4972
rect 253848 4208 253900 4214
rect 253676 4156 253848 4162
rect 253676 4150 253900 4156
rect 253676 4146 253888 4150
rect 253664 4140 253888 4146
rect 253716 4134 253888 4140
rect 253664 4082 253716 4088
rect 253952 3466 253980 4966
rect 254044 3942 254072 6258
rect 254584 6248 254636 6254
rect 254584 6190 254636 6196
rect 254400 6112 254452 6118
rect 254400 6054 254452 6060
rect 254412 5642 254440 6054
rect 254596 5846 254624 6190
rect 254584 5840 254636 5846
rect 254584 5782 254636 5788
rect 254676 5840 254728 5846
rect 254676 5782 254728 5788
rect 254308 5636 254360 5642
rect 254308 5578 254360 5584
rect 254400 5636 254452 5642
rect 254400 5578 254452 5584
rect 254216 5568 254268 5574
rect 254320 5545 254348 5578
rect 254216 5510 254268 5516
rect 254306 5536 254362 5545
rect 254228 5386 254256 5510
rect 254306 5471 254362 5480
rect 254228 5358 254348 5386
rect 254124 5296 254176 5302
rect 254124 5238 254176 5244
rect 254136 4146 254164 5238
rect 254124 4140 254176 4146
rect 254124 4082 254176 4088
rect 254032 3936 254084 3942
rect 254032 3878 254084 3884
rect 254124 3936 254176 3942
rect 254124 3878 254176 3884
rect 254136 3738 254164 3878
rect 254124 3732 254176 3738
rect 254124 3674 254176 3680
rect 254030 3632 254086 3641
rect 254030 3567 254032 3576
rect 254084 3567 254086 3576
rect 254032 3538 254084 3544
rect 254320 3466 254348 5358
rect 254492 5364 254544 5370
rect 254492 5306 254544 5312
rect 254504 5030 254532 5306
rect 254596 5166 254624 5782
rect 254688 5234 254716 5782
rect 255134 5400 255190 5409
rect 255134 5335 255190 5344
rect 255148 5234 255176 5335
rect 255332 5302 255360 6394
rect 255412 6316 255464 6322
rect 255412 6258 255464 6264
rect 255424 5710 255452 6258
rect 255792 6118 255820 6598
rect 256332 6384 256384 6390
rect 256332 6326 256384 6332
rect 255780 6112 255832 6118
rect 255780 6054 255832 6060
rect 256344 5914 256372 6326
rect 256424 6112 256476 6118
rect 256424 6054 256476 6060
rect 256516 6112 256568 6118
rect 256516 6054 256568 6060
rect 256332 5908 256384 5914
rect 256332 5850 256384 5856
rect 256344 5710 256372 5850
rect 255412 5704 255464 5710
rect 255412 5646 255464 5652
rect 256332 5704 256384 5710
rect 256332 5646 256384 5652
rect 255424 5302 255452 5646
rect 255688 5568 255740 5574
rect 255688 5510 255740 5516
rect 255320 5296 255372 5302
rect 255320 5238 255372 5244
rect 255412 5296 255464 5302
rect 255412 5238 255464 5244
rect 254676 5228 254728 5234
rect 254676 5170 254728 5176
rect 255136 5228 255188 5234
rect 255136 5170 255188 5176
rect 255424 5166 255452 5238
rect 254584 5160 254636 5166
rect 254584 5102 254636 5108
rect 255412 5160 255464 5166
rect 255412 5102 255464 5108
rect 254492 5024 254544 5030
rect 254492 4966 254544 4972
rect 254504 4758 254532 4966
rect 254492 4752 254544 4758
rect 254492 4694 254544 4700
rect 254596 4078 254624 5102
rect 255134 4584 255190 4593
rect 255134 4519 255190 4528
rect 254584 4072 254636 4078
rect 254584 4014 254636 4020
rect 255148 3602 255176 4519
rect 255136 3596 255188 3602
rect 255136 3538 255188 3544
rect 253940 3460 253992 3466
rect 253940 3402 253992 3408
rect 254308 3460 254360 3466
rect 254308 3402 254360 3408
rect 254124 3392 254176 3398
rect 254124 3334 254176 3340
rect 253848 2984 253900 2990
rect 253848 2926 253900 2932
rect 253480 2508 253532 2514
rect 253480 2450 253532 2456
rect 253112 2372 253164 2378
rect 253112 2314 253164 2320
rect 253124 1562 253152 2314
rect 253112 1556 253164 1562
rect 253112 1498 253164 1504
rect 252836 1012 252888 1018
rect 252836 954 252888 960
rect 252928 1012 252980 1018
rect 252928 954 252980 960
rect 251732 944 251784 950
rect 251732 886 251784 892
rect 253860 513 253888 2926
rect 254136 2281 254164 3334
rect 254860 2440 254912 2446
rect 254860 2382 254912 2388
rect 254122 2272 254178 2281
rect 254122 2207 254178 2216
rect 254124 1352 254176 1358
rect 254124 1294 254176 1300
rect 254136 610 254164 1294
rect 254872 649 254900 2382
rect 255700 2038 255728 5510
rect 256436 5370 256464 6054
rect 256424 5364 256476 5370
rect 256424 5306 256476 5312
rect 256436 5030 256464 5306
rect 255872 5024 255924 5030
rect 255872 4966 255924 4972
rect 256424 5024 256476 5030
rect 256424 4966 256476 4972
rect 255884 4622 255912 4966
rect 255872 4616 255924 4622
rect 255872 4558 255924 4564
rect 256424 4616 256476 4622
rect 256424 4558 256476 4564
rect 256436 4457 256464 4558
rect 256422 4448 256478 4457
rect 256422 4383 256478 4392
rect 256528 3210 256556 6054
rect 256620 4690 256648 6598
rect 256712 6458 256740 6734
rect 256700 6452 256752 6458
rect 256700 6394 256752 6400
rect 256792 6316 256844 6322
rect 256792 6258 256844 6264
rect 256700 6248 256752 6254
rect 256700 6190 256752 6196
rect 256712 5166 256740 6190
rect 256804 5846 256832 6258
rect 256792 5840 256844 5846
rect 256792 5782 256844 5788
rect 256804 5710 256832 5782
rect 256792 5704 256844 5710
rect 256792 5646 256844 5652
rect 257620 5704 257672 5710
rect 257620 5646 257672 5652
rect 257632 5234 257660 5646
rect 257804 5568 257856 5574
rect 257804 5510 257856 5516
rect 257344 5228 257396 5234
rect 257344 5170 257396 5176
rect 257620 5228 257672 5234
rect 257620 5170 257672 5176
rect 256700 5160 256752 5166
rect 256700 5102 256752 5108
rect 257356 4690 257384 5170
rect 257528 5160 257580 5166
rect 257448 5120 257528 5148
rect 256608 4684 256660 4690
rect 256608 4626 256660 4632
rect 257344 4684 257396 4690
rect 257344 4626 257396 4632
rect 257356 4146 257384 4626
rect 257448 4146 257476 5120
rect 257528 5102 257580 5108
rect 257632 4146 257660 5170
rect 257344 4140 257396 4146
rect 257344 4082 257396 4088
rect 257436 4140 257488 4146
rect 257436 4082 257488 4088
rect 257620 4140 257672 4146
rect 257620 4082 257672 4088
rect 257068 4072 257120 4078
rect 257120 4020 257476 4026
rect 257068 4014 257476 4020
rect 257080 3998 257476 4014
rect 257448 3942 257476 3998
rect 257344 3936 257396 3942
rect 257344 3878 257396 3884
rect 257436 3936 257488 3942
rect 257436 3878 257488 3884
rect 257356 3738 257384 3878
rect 257344 3732 257396 3738
rect 257344 3674 257396 3680
rect 256436 3182 256556 3210
rect 256436 2774 256464 3182
rect 256516 3052 256568 3058
rect 256516 2994 256568 3000
rect 256528 2961 256556 2994
rect 256514 2952 256570 2961
rect 256514 2887 256570 2896
rect 256436 2746 256556 2774
rect 256528 2582 256556 2746
rect 256516 2576 256568 2582
rect 256516 2518 256568 2524
rect 256424 2440 256476 2446
rect 256424 2382 256476 2388
rect 255228 2032 255280 2038
rect 255228 1974 255280 1980
rect 255688 2032 255740 2038
rect 255688 1974 255740 1980
rect 255240 1465 255268 1974
rect 255688 1760 255740 1766
rect 255688 1702 255740 1708
rect 255226 1456 255282 1465
rect 255226 1391 255282 1400
rect 255596 1352 255648 1358
rect 255596 1294 255648 1300
rect 255320 1284 255372 1290
rect 255320 1226 255372 1232
rect 255332 814 255360 1226
rect 255608 1034 255636 1294
rect 255700 1193 255728 1702
rect 255964 1352 256016 1358
rect 255964 1294 256016 1300
rect 255872 1284 255924 1290
rect 255792 1244 255872 1272
rect 255686 1184 255742 1193
rect 255686 1119 255742 1128
rect 255792 1034 255820 1244
rect 255872 1226 255924 1232
rect 255608 1006 255820 1034
rect 255320 808 255372 814
rect 255320 750 255372 756
rect 254858 640 254914 649
rect 254124 604 254176 610
rect 254858 575 254914 584
rect 254124 546 254176 552
rect 253846 504 253902 513
rect 251548 468 251600 474
rect 253846 439 253902 448
rect 251548 410 251600 416
rect 255976 377 256004 1294
rect 256436 406 256464 2382
rect 257528 2372 257580 2378
rect 257528 2314 257580 2320
rect 257540 1465 257568 2314
rect 257712 1760 257764 1766
rect 257712 1702 257764 1708
rect 257526 1456 257582 1465
rect 257724 1426 257752 1702
rect 257526 1391 257582 1400
rect 257712 1420 257764 1426
rect 257712 1362 257764 1368
rect 256700 1352 256752 1358
rect 256700 1294 256752 1300
rect 256792 1352 256844 1358
rect 256792 1294 256844 1300
rect 256712 542 256740 1294
rect 256804 649 256832 1294
rect 257816 1193 257844 5510
rect 257896 4208 257948 4214
rect 257896 4150 257948 4156
rect 257908 4010 257936 4150
rect 257896 4004 257948 4010
rect 257896 3946 257948 3952
rect 258000 1766 258028 9522
rect 258080 9376 258132 9382
rect 258080 9318 258132 9324
rect 258092 8498 258120 9318
rect 258276 8634 258304 10231
rect 258552 10130 258580 10610
rect 258632 10532 258684 10538
rect 258632 10474 258684 10480
rect 258540 10124 258592 10130
rect 258540 10066 258592 10072
rect 258644 9450 258672 10474
rect 259552 10464 259604 10470
rect 259552 10406 259604 10412
rect 261758 10432 261814 10441
rect 259182 10296 259238 10305
rect 259182 10231 259238 10240
rect 258908 10124 258960 10130
rect 258736 10084 258908 10112
rect 258736 9926 258764 10084
rect 258908 10066 258960 10072
rect 258724 9920 258776 9926
rect 258724 9862 258776 9868
rect 258816 9920 258868 9926
rect 258816 9862 258868 9868
rect 258828 9722 258856 9862
rect 259196 9722 259224 10231
rect 258816 9716 258868 9722
rect 258816 9658 258868 9664
rect 259184 9716 259236 9722
rect 259184 9658 259236 9664
rect 259368 9580 259420 9586
rect 259368 9522 259420 9528
rect 259184 9512 259236 9518
rect 259184 9454 259236 9460
rect 258632 9444 258684 9450
rect 258632 9386 258684 9392
rect 258724 9444 258776 9450
rect 258724 9386 258776 9392
rect 258736 9178 258764 9386
rect 258724 9172 258776 9178
rect 258724 9114 258776 9120
rect 259196 8974 259224 9454
rect 259380 9178 259408 9522
rect 259368 9172 259420 9178
rect 259368 9114 259420 9120
rect 259092 8968 259144 8974
rect 259092 8910 259144 8916
rect 259184 8968 259236 8974
rect 259184 8910 259236 8916
rect 258264 8628 258316 8634
rect 258264 8570 258316 8576
rect 258080 8492 258132 8498
rect 258080 8434 258132 8440
rect 258264 8492 258316 8498
rect 258264 8434 258316 8440
rect 258170 6760 258226 6769
rect 258170 6695 258226 6704
rect 258184 2990 258212 6695
rect 258276 6089 258304 8434
rect 258724 8288 258776 8294
rect 258724 8230 258776 8236
rect 258736 8022 258764 8230
rect 258724 8016 258776 8022
rect 258724 7958 258776 7964
rect 258908 6316 258960 6322
rect 258908 6258 258960 6264
rect 258816 6180 258868 6186
rect 258816 6122 258868 6128
rect 258262 6080 258318 6089
rect 258262 6015 258318 6024
rect 258262 5808 258318 5817
rect 258262 5743 258318 5752
rect 258276 4842 258304 5743
rect 258724 5160 258776 5166
rect 258724 5102 258776 5108
rect 258632 5092 258684 5098
rect 258632 5034 258684 5040
rect 258276 4814 258396 4842
rect 258644 4826 258672 5034
rect 258264 4548 258316 4554
rect 258264 4490 258316 4496
rect 258276 4282 258304 4490
rect 258264 4276 258316 4282
rect 258264 4218 258316 4224
rect 258172 2984 258224 2990
rect 258172 2926 258224 2932
rect 258264 2848 258316 2854
rect 258264 2790 258316 2796
rect 258172 1896 258224 1902
rect 258172 1838 258224 1844
rect 257988 1760 258040 1766
rect 257988 1702 258040 1708
rect 258000 1358 258028 1702
rect 258184 1601 258212 1838
rect 258170 1592 258226 1601
rect 258170 1527 258226 1536
rect 258276 1442 258304 2790
rect 258368 2378 258396 4814
rect 258632 4820 258684 4826
rect 258632 4762 258684 4768
rect 258540 4208 258592 4214
rect 258540 4150 258592 4156
rect 258446 3496 258502 3505
rect 258446 3431 258502 3440
rect 258356 2372 258408 2378
rect 258356 2314 258408 2320
rect 258460 1970 258488 3431
rect 258552 1970 258580 4150
rect 258644 3738 258672 4762
rect 258736 4690 258764 5102
rect 258828 5030 258856 6122
rect 258816 5024 258868 5030
rect 258816 4966 258868 4972
rect 258724 4684 258776 4690
rect 258724 4626 258776 4632
rect 258632 3732 258684 3738
rect 258632 3674 258684 3680
rect 258736 3602 258764 4626
rect 258816 3936 258868 3942
rect 258816 3878 258868 3884
rect 258724 3596 258776 3602
rect 258724 3538 258776 3544
rect 258828 2922 258856 3878
rect 258920 3398 258948 6258
rect 259000 3732 259052 3738
rect 259000 3674 259052 3680
rect 258908 3392 258960 3398
rect 258908 3334 258960 3340
rect 259012 3233 259040 3674
rect 258998 3224 259054 3233
rect 258998 3159 259054 3168
rect 258816 2916 258868 2922
rect 258816 2858 258868 2864
rect 259104 2854 259132 8910
rect 259196 8634 259224 8910
rect 259184 8628 259236 8634
rect 259184 8570 259236 8576
rect 259564 8090 259592 10406
rect 260196 10396 260248 10402
rect 261758 10367 261814 10376
rect 260196 10338 260248 10344
rect 259918 10296 259974 10305
rect 259644 10260 259696 10266
rect 259918 10231 259974 10240
rect 259644 10202 259696 10208
rect 259552 8084 259604 8090
rect 259552 8026 259604 8032
rect 259550 7032 259606 7041
rect 259550 6967 259606 6976
rect 259564 5846 259592 6967
rect 259656 6390 259684 10202
rect 259828 8968 259880 8974
rect 259828 8910 259880 8916
rect 259736 8832 259788 8838
rect 259736 8774 259788 8780
rect 259748 8498 259776 8774
rect 259736 8492 259788 8498
rect 259736 8434 259788 8440
rect 259736 8084 259788 8090
rect 259736 8026 259788 8032
rect 259748 7002 259776 8026
rect 259736 6996 259788 7002
rect 259736 6938 259788 6944
rect 259644 6384 259696 6390
rect 259644 6326 259696 6332
rect 259552 5840 259604 5846
rect 259552 5782 259604 5788
rect 259184 5704 259236 5710
rect 259564 5658 259592 5782
rect 259656 5710 259684 6326
rect 259840 5930 259868 8910
rect 259932 8634 259960 10231
rect 260208 9586 260236 10338
rect 260470 10296 260526 10305
rect 260470 10231 260526 10240
rect 260196 9580 260248 9586
rect 260196 9522 260248 9528
rect 260288 8832 260340 8838
rect 260288 8774 260340 8780
rect 259920 8628 259972 8634
rect 259920 8570 259972 8576
rect 260300 8498 260328 8774
rect 260484 8634 260512 10231
rect 261576 10056 261628 10062
rect 261576 9998 261628 10004
rect 261588 9518 261616 9998
rect 261392 9512 261444 9518
rect 261392 9454 261444 9460
rect 261576 9512 261628 9518
rect 261628 9472 261708 9500
rect 261576 9454 261628 9460
rect 260840 9444 260892 9450
rect 260840 9386 260892 9392
rect 260748 9036 260800 9042
rect 260748 8978 260800 8984
rect 260564 8968 260616 8974
rect 260564 8910 260616 8916
rect 260472 8628 260524 8634
rect 260472 8570 260524 8576
rect 260288 8492 260340 8498
rect 260288 8434 260340 8440
rect 260380 8492 260432 8498
rect 260380 8434 260432 8440
rect 260392 8362 260420 8434
rect 260380 8356 260432 8362
rect 260380 8298 260432 8304
rect 260380 6112 260432 6118
rect 260380 6054 260432 6060
rect 259840 5902 259960 5930
rect 259184 5646 259236 5652
rect 259196 4826 259224 5646
rect 259472 5642 259592 5658
rect 259644 5704 259696 5710
rect 259644 5646 259696 5652
rect 259460 5636 259592 5642
rect 259512 5630 259592 5636
rect 259460 5578 259512 5584
rect 259828 5568 259880 5574
rect 259828 5510 259880 5516
rect 259368 5228 259420 5234
rect 259368 5170 259420 5176
rect 259184 4820 259236 4826
rect 259184 4762 259236 4768
rect 259380 4622 259408 5170
rect 259840 4622 259868 5510
rect 259368 4616 259420 4622
rect 259368 4558 259420 4564
rect 259828 4616 259880 4622
rect 259828 4558 259880 4564
rect 259184 4548 259236 4554
rect 259184 4490 259236 4496
rect 259196 3618 259224 4490
rect 259276 4072 259328 4078
rect 259276 4014 259328 4020
rect 259288 3942 259316 4014
rect 259276 3936 259328 3942
rect 259276 3878 259328 3884
rect 259288 3777 259316 3878
rect 259274 3768 259330 3777
rect 259274 3703 259330 3712
rect 259196 3590 259316 3618
rect 259288 3466 259316 3590
rect 259380 3534 259408 4558
rect 259828 4480 259880 4486
rect 259828 4422 259880 4428
rect 259840 4214 259868 4422
rect 259828 4208 259880 4214
rect 259828 4150 259880 4156
rect 259368 3528 259420 3534
rect 259368 3470 259420 3476
rect 259276 3460 259328 3466
rect 259276 3402 259328 3408
rect 259736 3460 259788 3466
rect 259736 3402 259788 3408
rect 259748 3369 259776 3402
rect 259734 3360 259790 3369
rect 259734 3295 259790 3304
rect 259092 2848 259144 2854
rect 259092 2790 259144 2796
rect 259748 2582 259776 3295
rect 259828 2848 259880 2854
rect 259826 2816 259828 2825
rect 259880 2816 259882 2825
rect 259826 2751 259882 2760
rect 259736 2576 259788 2582
rect 259736 2518 259788 2524
rect 259932 2310 259960 5902
rect 260392 5710 260420 6054
rect 260380 5704 260432 5710
rect 260380 5646 260432 5652
rect 260288 5296 260340 5302
rect 260288 5238 260340 5244
rect 260104 5160 260156 5166
rect 260104 5102 260156 5108
rect 260010 4448 260066 4457
rect 260010 4383 260066 4392
rect 260024 3058 260052 4383
rect 260012 3052 260064 3058
rect 260012 2994 260064 3000
rect 260116 2378 260144 5102
rect 260300 4826 260328 5238
rect 260288 4820 260340 4826
rect 260288 4762 260340 4768
rect 260472 3392 260524 3398
rect 260472 3334 260524 3340
rect 260484 3058 260512 3334
rect 260472 3052 260524 3058
rect 260472 2994 260524 3000
rect 260576 2990 260604 8910
rect 260760 5642 260788 8978
rect 260852 8129 260880 9386
rect 261404 8430 261432 9454
rect 261484 9376 261536 9382
rect 261484 9318 261536 9324
rect 261576 9376 261628 9382
rect 261576 9318 261628 9324
rect 261496 8498 261524 9318
rect 261484 8492 261536 8498
rect 261484 8434 261536 8440
rect 260932 8424 260984 8430
rect 260932 8366 260984 8372
rect 261392 8424 261444 8430
rect 261392 8366 261444 8372
rect 260838 8120 260894 8129
rect 260838 8055 260894 8064
rect 260944 7177 260972 8366
rect 261404 7426 261432 8366
rect 261588 7886 261616 9318
rect 261680 9178 261708 9472
rect 261668 9172 261720 9178
rect 261668 9114 261720 9120
rect 261576 7880 261628 7886
rect 261576 7822 261628 7828
rect 261680 7834 261708 9114
rect 261772 8090 261800 10367
rect 261850 10296 261906 10305
rect 261850 10231 261906 10240
rect 262494 10296 262550 10305
rect 262494 10231 262550 10240
rect 263322 10296 263378 10305
rect 263322 10231 263378 10240
rect 261864 8634 261892 10231
rect 262128 9988 262180 9994
rect 262128 9930 262180 9936
rect 262140 9518 262168 9930
rect 262128 9512 262180 9518
rect 262128 9454 262180 9460
rect 262140 9178 262168 9454
rect 262312 9376 262364 9382
rect 262312 9318 262364 9324
rect 262128 9172 262180 9178
rect 262128 9114 262180 9120
rect 262036 8900 262088 8906
rect 262036 8842 262088 8848
rect 261852 8628 261904 8634
rect 261852 8570 261904 8576
rect 261760 8084 261812 8090
rect 261760 8026 261812 8032
rect 261680 7806 261892 7834
rect 261666 7440 261722 7449
rect 261404 7398 261524 7426
rect 260930 7168 260986 7177
rect 260986 7126 261064 7154
rect 260930 7103 260986 7112
rect 260840 6724 260892 6730
rect 260840 6666 260892 6672
rect 260852 6089 260880 6666
rect 260930 6624 260986 6633
rect 260930 6559 260986 6568
rect 260838 6080 260894 6089
rect 260838 6015 260894 6024
rect 260852 5914 260880 6015
rect 260840 5908 260892 5914
rect 260840 5850 260892 5856
rect 260944 5778 260972 6559
rect 260932 5772 260984 5778
rect 260932 5714 260984 5720
rect 261036 5642 261064 7126
rect 260748 5636 260800 5642
rect 260748 5578 260800 5584
rect 261024 5636 261076 5642
rect 261024 5578 261076 5584
rect 261022 5264 261078 5273
rect 261022 5199 261024 5208
rect 261076 5199 261078 5208
rect 261024 5170 261076 5176
rect 261392 5160 261444 5166
rect 261392 5102 261444 5108
rect 260840 4548 260892 4554
rect 260840 4490 260892 4496
rect 260852 4185 260880 4490
rect 260838 4176 260894 4185
rect 260838 4111 260894 4120
rect 260748 4072 260800 4078
rect 260748 4014 260800 4020
rect 260656 3528 260708 3534
rect 260656 3470 260708 3476
rect 260288 2984 260340 2990
rect 260288 2926 260340 2932
rect 260564 2984 260616 2990
rect 260564 2926 260616 2932
rect 260104 2372 260156 2378
rect 260104 2314 260156 2320
rect 259920 2304 259972 2310
rect 259920 2246 259972 2252
rect 258722 2000 258778 2009
rect 258448 1964 258500 1970
rect 258448 1906 258500 1912
rect 258540 1964 258592 1970
rect 258722 1935 258778 1944
rect 258540 1906 258592 1912
rect 258736 1465 258764 1935
rect 258722 1456 258778 1465
rect 258276 1426 258396 1442
rect 258276 1420 258408 1426
rect 258276 1414 258356 1420
rect 257988 1352 258040 1358
rect 257988 1294 258040 1300
rect 258172 1352 258224 1358
rect 258172 1294 258224 1300
rect 258184 1222 258212 1294
rect 258080 1216 258132 1222
rect 257802 1184 257858 1193
rect 258080 1158 258132 1164
rect 258172 1216 258224 1222
rect 258172 1158 258224 1164
rect 257802 1119 257858 1128
rect 258092 649 258120 1158
rect 258276 746 258304 1414
rect 258722 1391 258778 1400
rect 258356 1362 258408 1368
rect 259276 1352 259328 1358
rect 259276 1294 259328 1300
rect 259288 882 259316 1294
rect 259276 876 259328 882
rect 259276 818 259328 824
rect 260116 785 260144 2314
rect 260196 2304 260248 2310
rect 260196 2246 260248 2252
rect 260208 1902 260236 2246
rect 260300 2145 260328 2926
rect 260472 2916 260524 2922
rect 260472 2858 260524 2864
rect 260484 2825 260512 2858
rect 260470 2816 260526 2825
rect 260470 2751 260526 2760
rect 260286 2136 260342 2145
rect 260286 2071 260288 2080
rect 260340 2071 260342 2080
rect 260288 2042 260340 2048
rect 260472 1964 260524 1970
rect 260472 1906 260524 1912
rect 260196 1896 260248 1902
rect 260196 1838 260248 1844
rect 260102 776 260158 785
rect 258264 740 258316 746
rect 260102 711 260158 720
rect 258264 682 258316 688
rect 260208 678 260236 1838
rect 260484 921 260512 1906
rect 260668 1358 260696 3470
rect 260656 1352 260708 1358
rect 260656 1294 260708 1300
rect 260760 1018 260788 4014
rect 261024 3052 261076 3058
rect 261024 2994 261076 3000
rect 261116 3052 261168 3058
rect 261116 2994 261168 3000
rect 261036 2446 261064 2994
rect 261024 2440 261076 2446
rect 261024 2382 261076 2388
rect 261128 2106 261156 2994
rect 261116 2100 261168 2106
rect 261116 2042 261168 2048
rect 261404 1970 261432 5102
rect 261496 2774 261524 7398
rect 261576 7404 261628 7410
rect 261666 7375 261668 7384
rect 261576 7346 261628 7352
rect 261720 7375 261722 7384
rect 261668 7346 261720 7352
rect 261588 7002 261616 7346
rect 261576 6996 261628 7002
rect 261576 6938 261628 6944
rect 261758 6488 261814 6497
rect 261758 6423 261814 6432
rect 261772 6390 261800 6423
rect 261760 6384 261812 6390
rect 261760 6326 261812 6332
rect 261576 6316 261628 6322
rect 261576 6258 261628 6264
rect 261588 5778 261616 6258
rect 261760 6180 261812 6186
rect 261760 6122 261812 6128
rect 261668 6112 261720 6118
rect 261668 6054 261720 6060
rect 261576 5772 261628 5778
rect 261576 5714 261628 5720
rect 261588 5370 261616 5714
rect 261680 5710 261708 6054
rect 261668 5704 261720 5710
rect 261668 5646 261720 5652
rect 261576 5364 261628 5370
rect 261576 5306 261628 5312
rect 261588 4486 261616 5306
rect 261576 4480 261628 4486
rect 261576 4422 261628 4428
rect 261772 4146 261800 6122
rect 261760 4140 261812 4146
rect 261760 4082 261812 4088
rect 261760 3936 261812 3942
rect 261760 3878 261812 3884
rect 261496 2746 261616 2774
rect 261588 2514 261616 2746
rect 261576 2508 261628 2514
rect 261576 2450 261628 2456
rect 261484 2440 261536 2446
rect 261484 2382 261536 2388
rect 261496 1970 261524 2382
rect 261772 1970 261800 3878
rect 261392 1964 261444 1970
rect 261392 1906 261444 1912
rect 261484 1964 261536 1970
rect 261484 1906 261536 1912
rect 261760 1964 261812 1970
rect 261760 1906 261812 1912
rect 261496 1290 261524 1906
rect 261864 1426 261892 7806
rect 261944 6792 261996 6798
rect 261944 6734 261996 6740
rect 261956 6458 261984 6734
rect 262048 6497 262076 8842
rect 262034 6488 262090 6497
rect 261944 6452 261996 6458
rect 262034 6423 262090 6432
rect 261944 6394 261996 6400
rect 262140 6338 262168 9114
rect 262218 7984 262274 7993
rect 262218 7919 262274 7928
rect 262232 7750 262260 7919
rect 262324 7886 262352 9318
rect 262404 8424 262456 8430
rect 262404 8366 262456 8372
rect 262312 7880 262364 7886
rect 262312 7822 262364 7828
rect 262220 7744 262272 7750
rect 262220 7686 262272 7692
rect 262416 7546 262444 8366
rect 262508 8090 262536 10231
rect 262680 10056 262732 10062
rect 262680 9998 262732 10004
rect 262588 8628 262640 8634
rect 262588 8570 262640 8576
rect 262600 8265 262628 8570
rect 262586 8256 262642 8265
rect 262586 8191 262642 8200
rect 262496 8084 262548 8090
rect 262496 8026 262548 8032
rect 262404 7540 262456 7546
rect 262404 7482 262456 7488
rect 262312 7404 262364 7410
rect 262312 7346 262364 7352
rect 262324 7313 262352 7346
rect 262310 7304 262366 7313
rect 262310 7239 262366 7248
rect 262692 6769 262720 9998
rect 263232 9512 263284 9518
rect 263232 9454 263284 9460
rect 263244 9110 263272 9454
rect 263232 9104 263284 9110
rect 263232 9046 263284 9052
rect 262956 8968 263008 8974
rect 262956 8910 263008 8916
rect 262968 8294 262996 8910
rect 263140 8832 263192 8838
rect 263140 8774 263192 8780
rect 263048 8492 263100 8498
rect 263048 8434 263100 8440
rect 262956 8288 263008 8294
rect 262956 8230 263008 8236
rect 262772 7744 262824 7750
rect 262772 7686 262824 7692
rect 262784 7546 262812 7686
rect 262772 7540 262824 7546
rect 262772 7482 262824 7488
rect 262678 6760 262734 6769
rect 262678 6695 262734 6704
rect 262048 6310 262168 6338
rect 262496 6316 262548 6322
rect 262048 3942 262076 6310
rect 262496 6258 262548 6264
rect 262128 6248 262180 6254
rect 262128 6190 262180 6196
rect 262036 3936 262088 3942
rect 262036 3878 262088 3884
rect 262140 3398 262168 6190
rect 262508 5370 262536 6258
rect 262312 5364 262364 5370
rect 262312 5306 262364 5312
rect 262496 5364 262548 5370
rect 262496 5306 262548 5312
rect 262324 5234 262352 5306
rect 262312 5228 262364 5234
rect 262312 5170 262364 5176
rect 262588 5160 262640 5166
rect 262588 5102 262640 5108
rect 262128 3392 262180 3398
rect 262128 3334 262180 3340
rect 262600 2825 262628 5102
rect 262126 2816 262182 2825
rect 262586 2816 262642 2825
rect 262182 2760 262260 2774
rect 262126 2751 262260 2760
rect 262968 2774 262996 8230
rect 263060 7698 263088 8434
rect 263152 7886 263180 8774
rect 263232 8288 263284 8294
rect 263232 8230 263284 8236
rect 263244 8022 263272 8230
rect 263336 8090 263364 10231
rect 263600 9580 263652 9586
rect 263600 9522 263652 9528
rect 263612 8974 263640 9522
rect 263796 9450 263824 10678
rect 264428 10600 264480 10606
rect 264428 10542 264480 10548
rect 264334 10296 264390 10305
rect 264334 10231 264390 10240
rect 264244 9920 264296 9926
rect 264244 9862 264296 9868
rect 263968 9512 264020 9518
rect 263968 9454 264020 9460
rect 263692 9444 263744 9450
rect 263692 9386 263744 9392
rect 263784 9444 263836 9450
rect 263784 9386 263836 9392
rect 263704 9110 263732 9386
rect 263692 9104 263744 9110
rect 263692 9046 263744 9052
rect 263600 8968 263652 8974
rect 263600 8910 263652 8916
rect 263324 8084 263376 8090
rect 263324 8026 263376 8032
rect 263232 8016 263284 8022
rect 263232 7958 263284 7964
rect 263140 7880 263192 7886
rect 263796 7868 263824 9386
rect 263876 8968 263928 8974
rect 263876 8910 263928 8916
rect 263888 8566 263916 8910
rect 263876 8560 263928 8566
rect 263876 8502 263928 8508
rect 263874 8392 263930 8401
rect 263980 8362 264008 9454
rect 264152 9376 264204 9382
rect 264152 9318 264204 9324
rect 264060 9036 264112 9042
rect 264060 8978 264112 8984
rect 263874 8327 263876 8336
rect 263928 8327 263930 8336
rect 263968 8356 264020 8362
rect 263876 8298 263928 8304
rect 263968 8298 264020 8304
rect 264072 8294 264100 8978
rect 264060 8288 264112 8294
rect 263966 8256 264022 8265
rect 264060 8230 264112 8236
rect 263966 8191 264022 8200
rect 263876 7880 263928 7886
rect 263796 7840 263876 7868
rect 263140 7822 263192 7828
rect 263876 7822 263928 7828
rect 263060 7670 263180 7698
rect 263048 6656 263100 6662
rect 263152 6644 263180 7670
rect 263416 7540 263468 7546
rect 263416 7482 263468 7488
rect 263230 7168 263286 7177
rect 263230 7103 263286 7112
rect 263244 6798 263272 7103
rect 263232 6792 263284 6798
rect 263232 6734 263284 6740
rect 263152 6616 263272 6644
rect 263048 6598 263100 6604
rect 263060 6186 263088 6598
rect 263140 6316 263192 6322
rect 263140 6258 263192 6264
rect 263048 6180 263100 6186
rect 263048 6122 263100 6128
rect 263152 5914 263180 6258
rect 263244 6254 263272 6616
rect 263232 6248 263284 6254
rect 263232 6190 263284 6196
rect 263140 5908 263192 5914
rect 263140 5850 263192 5856
rect 263244 4865 263272 6190
rect 263428 5681 263456 7482
rect 263692 6792 263744 6798
rect 263692 6734 263744 6740
rect 263414 5672 263470 5681
rect 263414 5607 263470 5616
rect 263704 5370 263732 6734
rect 263784 6656 263836 6662
rect 263784 6598 263836 6604
rect 263796 6390 263824 6598
rect 263784 6384 263836 6390
rect 263784 6326 263836 6332
rect 263692 5364 263744 5370
rect 263692 5306 263744 5312
rect 263600 5228 263652 5234
rect 263600 5170 263652 5176
rect 263230 4856 263286 4865
rect 263230 4791 263286 4800
rect 263612 4554 263640 5170
rect 263600 4548 263652 4554
rect 263600 4490 263652 4496
rect 262586 2751 262642 2760
rect 262140 2746 262260 2751
rect 262232 2582 262260 2746
rect 262876 2746 262996 2774
rect 263888 2774 263916 7822
rect 263980 6866 264008 8191
rect 264164 7410 264192 9318
rect 264256 8566 264284 9862
rect 264244 8560 264296 8566
rect 264244 8502 264296 8508
rect 264244 8356 264296 8362
rect 264244 8298 264296 8304
rect 264060 7404 264112 7410
rect 264060 7346 264112 7352
rect 264152 7404 264204 7410
rect 264152 7346 264204 7352
rect 264072 6866 264100 7346
rect 264256 7290 264284 8298
rect 264348 7546 264376 10231
rect 264440 9586 264468 10542
rect 264428 9580 264480 9586
rect 264428 9522 264480 9528
rect 264336 7540 264388 7546
rect 264336 7482 264388 7488
rect 264336 7404 264388 7410
rect 264336 7346 264388 7352
rect 264164 7262 264284 7290
rect 263968 6860 264020 6866
rect 263968 6802 264020 6808
rect 264060 6860 264112 6866
rect 264060 6802 264112 6808
rect 264164 2774 264192 7262
rect 264348 4622 264376 7346
rect 264440 5710 264468 9522
rect 264716 9518 264744 10746
rect 266266 10432 266322 10441
rect 266266 10367 266322 10376
rect 266174 10296 266230 10305
rect 266174 10231 266230 10240
rect 265624 10192 265676 10198
rect 265624 10134 265676 10140
rect 264796 9988 264848 9994
rect 264796 9930 264848 9936
rect 264704 9512 264756 9518
rect 264704 9454 264756 9460
rect 264520 8560 264572 8566
rect 264520 8502 264572 8508
rect 264532 6254 264560 8502
rect 264612 6996 264664 7002
rect 264612 6938 264664 6944
rect 264520 6248 264572 6254
rect 264520 6190 264572 6196
rect 264428 5704 264480 5710
rect 264428 5646 264480 5652
rect 264624 5234 264652 6938
rect 264612 5228 264664 5234
rect 264612 5170 264664 5176
rect 264336 4616 264388 4622
rect 264336 4558 264388 4564
rect 264244 3188 264296 3194
rect 264244 3130 264296 3136
rect 263888 2746 264008 2774
rect 262220 2576 262272 2582
rect 262220 2518 262272 2524
rect 262876 1970 262904 2746
rect 263980 2514 264008 2746
rect 264072 2746 264192 2774
rect 263968 2508 264020 2514
rect 263968 2450 264020 2456
rect 263140 2440 263192 2446
rect 263140 2382 263192 2388
rect 263152 2106 263180 2382
rect 263968 2372 264020 2378
rect 263968 2314 264020 2320
rect 263324 2304 263376 2310
rect 263324 2246 263376 2252
rect 263140 2100 263192 2106
rect 263140 2042 263192 2048
rect 262864 1964 262916 1970
rect 262864 1906 262916 1912
rect 263140 1760 263192 1766
rect 263140 1702 263192 1708
rect 261852 1420 261904 1426
rect 261852 1362 261904 1368
rect 263152 1358 263180 1702
rect 263140 1352 263192 1358
rect 263140 1294 263192 1300
rect 261484 1284 261536 1290
rect 261484 1226 261536 1232
rect 261116 1216 261168 1222
rect 261116 1158 261168 1164
rect 262864 1216 262916 1222
rect 262864 1158 262916 1164
rect 260748 1012 260800 1018
rect 260748 954 260800 960
rect 260470 912 260526 921
rect 260470 847 260526 856
rect 260196 672 260248 678
rect 256790 640 256846 649
rect 256790 575 256846 584
rect 258078 640 258134 649
rect 261128 649 261156 1158
rect 262876 649 262904 1158
rect 263336 649 263364 2246
rect 263980 2038 264008 2314
rect 263968 2032 264020 2038
rect 263968 1974 264020 1980
rect 264072 1970 264100 2746
rect 264256 2378 264284 3130
rect 264716 2774 264744 9454
rect 264808 7410 264836 9930
rect 265440 9920 265492 9926
rect 265440 9862 265492 9868
rect 264980 9648 265032 9654
rect 264980 9590 265032 9596
rect 264886 8120 264942 8129
rect 264886 8055 264888 8064
rect 264940 8055 264942 8064
rect 264888 8026 264940 8032
rect 264886 7848 264942 7857
rect 264886 7783 264888 7792
rect 264940 7783 264942 7792
rect 264888 7754 264940 7760
rect 264796 7404 264848 7410
rect 264796 7346 264848 7352
rect 264992 6882 265020 9590
rect 265256 9580 265308 9586
rect 265256 9522 265308 9528
rect 265072 9172 265124 9178
rect 265072 9114 265124 9120
rect 264900 6854 265020 6882
rect 264900 6730 264928 6854
rect 264888 6724 264940 6730
rect 264888 6666 264940 6672
rect 264796 6452 264848 6458
rect 264796 6394 264848 6400
rect 264808 5953 264836 6394
rect 264794 5944 264850 5953
rect 264900 5914 264928 6666
rect 264794 5879 264850 5888
rect 264888 5908 264940 5914
rect 264888 5850 264940 5856
rect 264980 5772 265032 5778
rect 264980 5714 265032 5720
rect 264888 5704 264940 5710
rect 264888 5646 264940 5652
rect 264900 5250 264928 5646
rect 264992 5370 265020 5714
rect 264980 5364 265032 5370
rect 264980 5306 265032 5312
rect 264900 5222 265020 5250
rect 264992 5030 265020 5222
rect 264980 5024 265032 5030
rect 264980 4966 265032 4972
rect 265084 4622 265112 9114
rect 265268 8974 265296 9522
rect 265256 8968 265308 8974
rect 265256 8910 265308 8916
rect 265164 8288 265216 8294
rect 265164 8230 265216 8236
rect 265176 4826 265204 8230
rect 265256 8084 265308 8090
rect 265256 8026 265308 8032
rect 265268 7410 265296 8026
rect 265346 7712 265402 7721
rect 265346 7647 265402 7656
rect 265360 7546 265388 7647
rect 265348 7540 265400 7546
rect 265348 7482 265400 7488
rect 265256 7404 265308 7410
rect 265256 7346 265308 7352
rect 265256 6316 265308 6322
rect 265256 6258 265308 6264
rect 265268 5914 265296 6258
rect 265452 5914 265480 9862
rect 265532 9376 265584 9382
rect 265532 9318 265584 9324
rect 265256 5908 265308 5914
rect 265256 5850 265308 5856
rect 265440 5908 265492 5914
rect 265440 5850 265492 5856
rect 265256 5772 265308 5778
rect 265256 5714 265308 5720
rect 265268 5234 265296 5714
rect 265256 5228 265308 5234
rect 265256 5170 265308 5176
rect 265348 5092 265400 5098
rect 265348 5034 265400 5040
rect 265360 4826 265388 5034
rect 265164 4820 265216 4826
rect 265164 4762 265216 4768
rect 265348 4820 265400 4826
rect 265348 4762 265400 4768
rect 265072 4616 265124 4622
rect 265072 4558 265124 4564
rect 265544 4146 265572 9318
rect 265636 8634 265664 10134
rect 265624 8628 265676 8634
rect 265624 8570 265676 8576
rect 265636 7886 265664 8570
rect 265900 8560 265952 8566
rect 265900 8502 265952 8508
rect 265716 8492 265768 8498
rect 265716 8434 265768 8440
rect 265808 8492 265860 8498
rect 265808 8434 265860 8440
rect 265624 7880 265676 7886
rect 265624 7822 265676 7828
rect 265532 4140 265584 4146
rect 265532 4082 265584 4088
rect 264796 3936 264848 3942
rect 264796 3878 264848 3884
rect 264808 3738 264836 3878
rect 264796 3732 264848 3738
rect 264796 3674 264848 3680
rect 264440 2746 264744 2774
rect 265636 2774 265664 7822
rect 265728 6254 265756 8434
rect 265716 6248 265768 6254
rect 265716 6190 265768 6196
rect 265716 5704 265768 5710
rect 265716 5646 265768 5652
rect 265728 5574 265756 5646
rect 265716 5568 265768 5574
rect 265716 5510 265768 5516
rect 265716 5024 265768 5030
rect 265716 4966 265768 4972
rect 265728 4826 265756 4966
rect 265716 4820 265768 4826
rect 265716 4762 265768 4768
rect 265820 3942 265848 8434
rect 265912 6798 265940 8502
rect 265992 7744 266044 7750
rect 265992 7686 266044 7692
rect 266004 7410 266032 7686
rect 266188 7546 266216 10231
rect 266280 9722 266308 10367
rect 266544 10124 266596 10130
rect 266544 10066 266596 10072
rect 266268 9716 266320 9722
rect 266268 9658 266320 9664
rect 266360 9376 266412 9382
rect 266360 9318 266412 9324
rect 266268 8628 266320 8634
rect 266268 8570 266320 8576
rect 266176 7540 266228 7546
rect 266176 7482 266228 7488
rect 265992 7404 266044 7410
rect 265992 7346 266044 7352
rect 266280 7206 266308 8570
rect 266372 8090 266400 9318
rect 266452 8968 266504 8974
rect 266452 8910 266504 8916
rect 266464 8838 266492 8910
rect 266556 8838 266584 10066
rect 266924 9518 266952 10814
rect 267556 10668 267608 10674
rect 267556 10610 267608 10616
rect 267004 10532 267056 10538
rect 267004 10474 267056 10480
rect 267016 9722 267044 10474
rect 267096 10260 267148 10266
rect 267096 10202 267148 10208
rect 267004 9716 267056 9722
rect 267004 9658 267056 9664
rect 266912 9512 266964 9518
rect 266912 9454 266964 9460
rect 266728 8900 266780 8906
rect 266728 8842 266780 8848
rect 266452 8832 266504 8838
rect 266452 8774 266504 8780
rect 266544 8832 266596 8838
rect 266544 8774 266596 8780
rect 266360 8084 266412 8090
rect 266360 8026 266412 8032
rect 266268 7200 266320 7206
rect 266268 7142 266320 7148
rect 266358 6896 266414 6905
rect 266358 6831 266414 6840
rect 265900 6792 265952 6798
rect 265900 6734 265952 6740
rect 265990 6760 266046 6769
rect 265990 6695 266046 6704
rect 266004 6662 266032 6695
rect 266372 6662 266400 6831
rect 265992 6656 266044 6662
rect 265992 6598 266044 6604
rect 266360 6656 266412 6662
rect 266360 6598 266412 6604
rect 265900 5908 265952 5914
rect 265900 5850 265952 5856
rect 266176 5908 266228 5914
rect 266176 5850 266228 5856
rect 265808 3936 265860 3942
rect 265808 3878 265860 3884
rect 265912 3602 265940 5850
rect 265992 5568 266044 5574
rect 265992 5510 266044 5516
rect 266004 5302 266032 5510
rect 265992 5296 266044 5302
rect 265992 5238 266044 5244
rect 266188 4622 266216 5850
rect 266358 5808 266414 5817
rect 266464 5794 266492 8774
rect 266556 8430 266584 8774
rect 266740 8498 266768 8842
rect 266728 8492 266780 8498
rect 266728 8434 266780 8440
rect 266544 8424 266596 8430
rect 266544 8366 266596 8372
rect 266556 7528 266584 8366
rect 267016 8022 267044 9658
rect 267108 8634 267136 10202
rect 267568 9518 267596 10610
rect 269028 10464 269080 10470
rect 269028 10406 269080 10412
rect 268292 10396 268344 10402
rect 268292 10338 268344 10344
rect 268108 10328 268160 10334
rect 268108 10270 268160 10276
rect 267740 9920 267792 9926
rect 267740 9862 267792 9868
rect 268120 9874 268148 10270
rect 268198 10024 268254 10033
rect 268198 9959 268200 9968
rect 268252 9959 268254 9968
rect 268200 9930 268252 9936
rect 267648 9580 267700 9586
rect 267648 9522 267700 9528
rect 267464 9512 267516 9518
rect 267556 9512 267608 9518
rect 267464 9454 267516 9460
rect 267554 9480 267556 9489
rect 267608 9480 267610 9489
rect 267188 9036 267240 9042
rect 267188 8978 267240 8984
rect 267280 9036 267332 9042
rect 267280 8978 267332 8984
rect 267200 8906 267228 8978
rect 267188 8900 267240 8906
rect 267188 8842 267240 8848
rect 267096 8628 267148 8634
rect 267096 8570 267148 8576
rect 267004 8016 267056 8022
rect 266924 7976 267004 8004
rect 266556 7500 266768 7528
rect 266636 6656 266688 6662
rect 266636 6598 266688 6604
rect 266648 6322 266676 6598
rect 266544 6316 266596 6322
rect 266544 6258 266596 6264
rect 266636 6316 266688 6322
rect 266636 6258 266688 6264
rect 266414 5766 266492 5794
rect 266358 5743 266414 5752
rect 266372 5642 266400 5743
rect 266360 5636 266412 5642
rect 266360 5578 266412 5584
rect 266556 5370 266584 6258
rect 266544 5364 266596 5370
rect 266544 5306 266596 5312
rect 266452 5228 266504 5234
rect 266452 5170 266504 5176
rect 266544 5228 266596 5234
rect 266544 5170 266596 5176
rect 266176 4616 266228 4622
rect 266176 4558 266228 4564
rect 266464 4282 266492 5170
rect 266268 4276 266320 4282
rect 266268 4218 266320 4224
rect 266452 4276 266504 4282
rect 266452 4218 266504 4224
rect 266280 4049 266308 4218
rect 266266 4040 266322 4049
rect 266266 3975 266322 3984
rect 266556 3602 266584 5170
rect 265900 3596 265952 3602
rect 265900 3538 265952 3544
rect 266544 3596 266596 3602
rect 266544 3538 266596 3544
rect 266740 2774 266768 7500
rect 266924 7290 266952 7976
rect 267004 7958 267056 7964
rect 267096 7336 267148 7342
rect 266924 7262 267044 7290
rect 267096 7278 267148 7284
rect 266912 7200 266964 7206
rect 266912 7142 266964 7148
rect 266820 6792 266872 6798
rect 266820 6734 266872 6740
rect 266832 6458 266860 6734
rect 266820 6452 266872 6458
rect 266820 6394 266872 6400
rect 266924 5710 266952 7142
rect 266912 5704 266964 5710
rect 266912 5646 266964 5652
rect 266912 5296 266964 5302
rect 266910 5264 266912 5273
rect 266964 5264 266966 5273
rect 266910 5199 266966 5208
rect 267016 4978 267044 7262
rect 267108 5574 267136 7278
rect 267200 6322 267228 8842
rect 267292 8430 267320 8978
rect 267372 8900 267424 8906
rect 267372 8842 267424 8848
rect 267280 8424 267332 8430
rect 267278 8392 267280 8401
rect 267332 8392 267334 8401
rect 267278 8327 267334 8336
rect 267280 7404 267332 7410
rect 267280 7346 267332 7352
rect 267292 6798 267320 7346
rect 267280 6792 267332 6798
rect 267280 6734 267332 6740
rect 267188 6316 267240 6322
rect 267188 6258 267240 6264
rect 267096 5568 267148 5574
rect 267096 5510 267148 5516
rect 267292 5234 267320 6734
rect 267280 5228 267332 5234
rect 267280 5170 267332 5176
rect 267384 5114 267412 8842
rect 267476 8838 267504 9454
rect 267554 9415 267610 9424
rect 267464 8832 267516 8838
rect 267464 8774 267516 8780
rect 267200 5086 267412 5114
rect 266832 4950 267044 4978
rect 267096 5024 267148 5030
rect 267096 4966 267148 4972
rect 266832 2922 266860 4950
rect 266912 4820 266964 4826
rect 266912 4762 266964 4768
rect 266924 4146 266952 4762
rect 267108 4146 267136 4966
rect 267200 4554 267228 5086
rect 267476 4978 267504 8774
rect 267660 8498 267688 9522
rect 267752 9489 267780 9862
rect 268120 9846 268240 9874
rect 268106 9752 268162 9761
rect 268106 9687 268162 9696
rect 267738 9480 267794 9489
rect 267738 9415 267794 9424
rect 268014 9344 268070 9353
rect 268014 9279 268070 9288
rect 267924 9104 267976 9110
rect 267924 9046 267976 9052
rect 267936 8974 267964 9046
rect 267924 8968 267976 8974
rect 267924 8910 267976 8916
rect 268028 8906 268056 9279
rect 268016 8900 268068 8906
rect 268016 8842 268068 8848
rect 268016 8560 268068 8566
rect 268016 8502 268068 8508
rect 267648 8492 267700 8498
rect 267648 8434 267700 8440
rect 267556 7880 267608 7886
rect 267660 7868 267688 8434
rect 268028 8401 268056 8502
rect 268014 8392 268070 8401
rect 268014 8327 268070 8336
rect 268016 8016 268068 8022
rect 267738 7984 267794 7993
rect 267738 7919 267740 7928
rect 267792 7919 267794 7928
rect 268014 7984 268016 7993
rect 268068 7984 268070 7993
rect 268014 7919 268070 7928
rect 267740 7890 267792 7896
rect 267608 7840 267688 7868
rect 267556 7822 267608 7828
rect 267568 6798 267596 7822
rect 268016 7744 268068 7750
rect 267922 7712 267978 7721
rect 267752 7670 267922 7698
rect 267752 7154 267780 7670
rect 268016 7686 268068 7692
rect 267922 7647 267978 7656
rect 267924 7472 267976 7478
rect 267924 7414 267976 7420
rect 267660 7126 267780 7154
rect 267832 7200 267884 7206
rect 267832 7142 267884 7148
rect 267660 7002 267688 7126
rect 267738 7032 267794 7041
rect 267648 6996 267700 7002
rect 267738 6967 267740 6976
rect 267648 6938 267700 6944
rect 267792 6967 267794 6976
rect 267740 6938 267792 6944
rect 267556 6792 267608 6798
rect 267556 6734 267608 6740
rect 267646 6760 267702 6769
rect 267646 6695 267702 6704
rect 267740 6724 267792 6730
rect 267660 6662 267688 6695
rect 267740 6666 267792 6672
rect 267648 6656 267700 6662
rect 267648 6598 267700 6604
rect 267648 6112 267700 6118
rect 267648 6054 267700 6060
rect 267660 5545 267688 6054
rect 267646 5536 267702 5545
rect 267646 5471 267702 5480
rect 267752 5370 267780 6666
rect 267844 6322 267872 7142
rect 267936 7041 267964 7414
rect 267922 7032 267978 7041
rect 267922 6967 267978 6976
rect 267922 6896 267978 6905
rect 267922 6831 267924 6840
rect 267976 6831 267978 6840
rect 267924 6802 267976 6808
rect 268028 6798 268056 7686
rect 268120 7290 268148 9687
rect 268212 8378 268240 9846
rect 268304 8537 268332 10338
rect 268384 10056 268436 10062
rect 268384 9998 268436 10004
rect 268290 8528 268346 8537
rect 268396 8498 268424 9998
rect 268842 9752 268898 9761
rect 268842 9687 268898 9696
rect 268856 9518 268884 9687
rect 268936 9580 268988 9586
rect 268936 9522 268988 9528
rect 268476 9512 268528 9518
rect 268476 9454 268528 9460
rect 268568 9512 268620 9518
rect 268568 9454 268620 9460
rect 268844 9512 268896 9518
rect 268844 9454 268896 9460
rect 268488 9110 268516 9454
rect 268476 9104 268528 9110
rect 268476 9046 268528 9052
rect 268290 8463 268346 8472
rect 268384 8492 268436 8498
rect 268384 8434 268436 8440
rect 268212 8350 268516 8378
rect 268488 8294 268516 8350
rect 268384 8288 268436 8294
rect 268384 8230 268436 8236
rect 268476 8288 268528 8294
rect 268476 8230 268528 8236
rect 268290 8120 268346 8129
rect 268290 8055 268346 8064
rect 268200 7880 268252 7886
rect 268200 7822 268252 7828
rect 268212 7410 268240 7822
rect 268200 7404 268252 7410
rect 268200 7346 268252 7352
rect 268120 7262 268240 7290
rect 268212 6882 268240 7262
rect 268304 6934 268332 8055
rect 268396 7970 268424 8230
rect 268396 7942 268516 7970
rect 268488 7886 268516 7942
rect 268384 7880 268436 7886
rect 268384 7822 268436 7828
rect 268476 7880 268528 7886
rect 268476 7822 268528 7828
rect 268120 6854 268240 6882
rect 268292 6928 268344 6934
rect 268292 6870 268344 6876
rect 268016 6792 268068 6798
rect 268016 6734 268068 6740
rect 268120 6610 268148 6854
rect 268396 6780 268424 7822
rect 268476 7540 268528 7546
rect 268476 7482 268528 7488
rect 268028 6582 268148 6610
rect 268212 6752 268424 6780
rect 267832 6316 267884 6322
rect 267832 6258 267884 6264
rect 268028 5642 268056 6582
rect 268106 6488 268162 6497
rect 268106 6423 268162 6432
rect 268016 5636 268068 5642
rect 268016 5578 268068 5584
rect 267740 5364 267792 5370
rect 267740 5306 267792 5312
rect 267556 5228 267608 5234
rect 267556 5170 267608 5176
rect 267568 5030 267596 5170
rect 267832 5160 267884 5166
rect 267832 5102 267884 5108
rect 267384 4950 267504 4978
rect 267556 5024 267608 5030
rect 267556 4966 267608 4972
rect 267738 4992 267794 5001
rect 267188 4548 267240 4554
rect 267188 4490 267240 4496
rect 267280 4548 267332 4554
rect 267280 4490 267332 4496
rect 267292 4457 267320 4490
rect 267278 4448 267334 4457
rect 267278 4383 267334 4392
rect 266912 4140 266964 4146
rect 266912 4082 266964 4088
rect 267004 4140 267056 4146
rect 267004 4082 267056 4088
rect 267096 4140 267148 4146
rect 267096 4082 267148 4088
rect 266820 2916 266872 2922
rect 266820 2858 266872 2864
rect 265636 2746 265848 2774
rect 264336 2440 264388 2446
rect 264336 2382 264388 2388
rect 264244 2372 264296 2378
rect 264244 2314 264296 2320
rect 264348 1970 264376 2382
rect 264440 1970 264468 2746
rect 265164 2440 265216 2446
rect 265164 2382 265216 2388
rect 264888 2304 264940 2310
rect 264888 2246 264940 2252
rect 264060 1964 264112 1970
rect 264060 1906 264112 1912
rect 264336 1964 264388 1970
rect 264336 1906 264388 1912
rect 264428 1964 264480 1970
rect 264428 1906 264480 1912
rect 264152 1760 264204 1766
rect 264152 1702 264204 1708
rect 264164 1358 264192 1702
rect 264900 1358 264928 2246
rect 265176 1970 265204 2382
rect 265820 1970 265848 2746
rect 266556 2746 266768 2774
rect 266556 1970 266584 2746
rect 267016 2650 267044 4082
rect 267280 4072 267332 4078
rect 267280 4014 267332 4020
rect 267292 3194 267320 4014
rect 267280 3188 267332 3194
rect 267280 3130 267332 3136
rect 267004 2644 267056 2650
rect 267004 2586 267056 2592
rect 267004 2440 267056 2446
rect 267004 2382 267056 2388
rect 266912 2304 266964 2310
rect 266912 2246 266964 2252
rect 265164 1964 265216 1970
rect 265164 1906 265216 1912
rect 265808 1964 265860 1970
rect 265808 1906 265860 1912
rect 266544 1964 266596 1970
rect 266544 1906 266596 1912
rect 265624 1760 265676 1766
rect 265624 1702 265676 1708
rect 266728 1760 266780 1766
rect 266728 1702 266780 1708
rect 265636 1358 265664 1702
rect 266740 1358 266768 1702
rect 264152 1352 264204 1358
rect 264152 1294 264204 1300
rect 264888 1352 264940 1358
rect 264888 1294 264940 1300
rect 265624 1352 265676 1358
rect 265624 1294 265676 1300
rect 266728 1352 266780 1358
rect 266728 1294 266780 1300
rect 264336 1216 264388 1222
rect 264336 1158 264388 1164
rect 264980 1216 265032 1222
rect 264980 1158 265032 1164
rect 265808 1216 265860 1222
rect 265808 1158 265860 1164
rect 266360 1216 266412 1222
rect 266360 1158 266412 1164
rect 264348 649 264376 1158
rect 264992 649 265020 1158
rect 265820 649 265848 1158
rect 266372 649 266400 1158
rect 266924 649 266952 2246
rect 267016 1970 267044 2382
rect 267384 1970 267412 4950
rect 267738 4927 267794 4936
rect 267752 4706 267780 4927
rect 267476 4678 267780 4706
rect 267476 3534 267504 4678
rect 267648 4616 267700 4622
rect 267648 4558 267700 4564
rect 267738 4584 267794 4593
rect 267556 4548 267608 4554
rect 267556 4490 267608 4496
rect 267464 3528 267516 3534
rect 267568 3505 267596 4490
rect 267660 4026 267688 4558
rect 267738 4519 267794 4528
rect 267752 4214 267780 4519
rect 267740 4208 267792 4214
rect 267740 4150 267792 4156
rect 267660 3998 267780 4026
rect 267752 3942 267780 3998
rect 267740 3936 267792 3942
rect 267740 3878 267792 3884
rect 267738 3768 267794 3777
rect 267738 3703 267740 3712
rect 267792 3703 267794 3712
rect 267740 3674 267792 3680
rect 267464 3470 267516 3476
rect 267554 3496 267610 3505
rect 267554 3431 267610 3440
rect 267740 3392 267792 3398
rect 267740 3334 267792 3340
rect 267752 3058 267780 3334
rect 267844 3194 267872 5102
rect 268014 3768 268070 3777
rect 268014 3703 268070 3712
rect 268028 3670 268056 3703
rect 268016 3664 268068 3670
rect 268016 3606 268068 3612
rect 268120 3534 268148 6423
rect 268212 5658 268240 6752
rect 268488 6089 268516 7482
rect 268474 6080 268530 6089
rect 268474 6015 268530 6024
rect 268384 5840 268436 5846
rect 268290 5808 268346 5817
rect 268384 5782 268436 5788
rect 268290 5743 268292 5752
rect 268344 5743 268346 5752
rect 268292 5714 268344 5720
rect 268212 5630 268332 5658
rect 268304 5234 268332 5630
rect 268396 5370 268424 5782
rect 268474 5672 268530 5681
rect 268474 5607 268530 5616
rect 268384 5364 268436 5370
rect 268384 5306 268436 5312
rect 268488 5234 268516 5607
rect 268292 5228 268344 5234
rect 268292 5170 268344 5176
rect 268476 5228 268528 5234
rect 268476 5170 268528 5176
rect 268200 5160 268252 5166
rect 268200 5102 268252 5108
rect 268474 5128 268530 5137
rect 268212 3738 268240 5102
rect 268474 5063 268530 5072
rect 268290 4720 268346 4729
rect 268488 4690 268516 5063
rect 268290 4655 268346 4664
rect 268476 4684 268528 4690
rect 268200 3732 268252 3738
rect 268200 3674 268252 3680
rect 268108 3528 268160 3534
rect 268014 3496 268070 3505
rect 267924 3460 267976 3466
rect 268108 3470 268160 3476
rect 268014 3431 268070 3440
rect 267924 3402 267976 3408
rect 267832 3188 267884 3194
rect 267832 3130 267884 3136
rect 267936 3097 267964 3402
rect 268028 3126 268056 3431
rect 268016 3120 268068 3126
rect 267922 3088 267978 3097
rect 267740 3052 267792 3058
rect 268016 3062 268068 3068
rect 267922 3023 267978 3032
rect 267740 2994 267792 3000
rect 267556 2916 267608 2922
rect 267556 2858 267608 2864
rect 267568 2514 267596 2858
rect 267648 2848 267700 2854
rect 267924 2848 267976 2854
rect 267648 2790 267700 2796
rect 267922 2816 267924 2825
rect 267976 2816 267978 2825
rect 267556 2508 267608 2514
rect 267556 2450 267608 2456
rect 267004 1964 267056 1970
rect 267004 1906 267056 1912
rect 267372 1964 267424 1970
rect 267372 1906 267424 1912
rect 267660 1306 267688 2790
rect 267922 2751 267978 2760
rect 267922 2680 267978 2689
rect 267922 2615 267978 2624
rect 267936 2582 267964 2615
rect 267924 2576 267976 2582
rect 267924 2518 267976 2524
rect 268304 2446 268332 4655
rect 268476 4626 268528 4632
rect 268474 4448 268530 4457
rect 268474 4383 268530 4392
rect 268382 2544 268438 2553
rect 268382 2479 268438 2488
rect 268292 2440 268344 2446
rect 268292 2382 268344 2388
rect 268396 2378 268424 2479
rect 268488 2446 268516 4383
rect 268580 4282 268608 9454
rect 268752 9444 268804 9450
rect 268752 9386 268804 9392
rect 268764 9217 268792 9386
rect 268750 9208 268806 9217
rect 268660 9172 268712 9178
rect 268750 9143 268806 9152
rect 268660 9114 268712 9120
rect 268672 9081 268700 9114
rect 268658 9072 268714 9081
rect 268658 9007 268714 9016
rect 268752 8492 268804 8498
rect 268752 8434 268804 8440
rect 268658 7712 268714 7721
rect 268658 7647 268714 7656
rect 268672 5953 268700 7647
rect 268764 6866 268792 8434
rect 268844 8084 268896 8090
rect 268844 8026 268896 8032
rect 268856 7478 268884 8026
rect 268948 7886 268976 9522
rect 269040 8945 269068 10406
rect 272154 10024 272210 10033
rect 272154 9959 272210 9968
rect 271337 9820 271645 9829
rect 271337 9818 271343 9820
rect 271399 9818 271423 9820
rect 271479 9818 271503 9820
rect 271559 9818 271583 9820
rect 271639 9818 271645 9820
rect 271399 9766 271401 9818
rect 271581 9766 271583 9818
rect 271337 9764 271343 9766
rect 271399 9764 271423 9766
rect 271479 9764 271503 9766
rect 271559 9764 271583 9766
rect 271639 9764 271645 9766
rect 271337 9755 271645 9764
rect 270408 9716 270460 9722
rect 270408 9658 270460 9664
rect 269948 9648 270000 9654
rect 269948 9590 270000 9596
rect 269856 9512 269908 9518
rect 269856 9454 269908 9460
rect 269212 9376 269264 9382
rect 269212 9318 269264 9324
rect 269672 9376 269724 9382
rect 269672 9318 269724 9324
rect 269026 8936 269082 8945
rect 269026 8871 269082 8880
rect 269224 8838 269252 9318
rect 269684 9042 269712 9318
rect 269672 9036 269724 9042
rect 269672 8978 269724 8984
rect 269028 8832 269080 8838
rect 269028 8774 269080 8780
rect 269212 8832 269264 8838
rect 269212 8774 269264 8780
rect 268936 7880 268988 7886
rect 268936 7822 268988 7828
rect 268844 7472 268896 7478
rect 268844 7414 268896 7420
rect 268752 6860 268804 6866
rect 268752 6802 268804 6808
rect 268750 6352 268806 6361
rect 268750 6287 268806 6296
rect 268658 5944 268714 5953
rect 268658 5879 268714 5888
rect 268658 5536 268714 5545
rect 268658 5471 268714 5480
rect 268568 4276 268620 4282
rect 268568 4218 268620 4224
rect 268566 3360 268622 3369
rect 268566 3295 268622 3304
rect 268476 2440 268528 2446
rect 268476 2382 268528 2388
rect 268384 2372 268436 2378
rect 268384 2314 268436 2320
rect 267738 2136 267794 2145
rect 267738 2071 267794 2080
rect 267752 1970 267780 2071
rect 268580 2038 268608 3295
rect 268672 3126 268700 5471
rect 268764 3534 268792 6287
rect 268856 6186 268884 7414
rect 269040 6746 269068 8774
rect 269304 8424 269356 8430
rect 269304 8366 269356 8372
rect 269212 7744 269264 7750
rect 269212 7686 269264 7692
rect 269120 7200 269172 7206
rect 269120 7142 269172 7148
rect 268948 6718 269068 6746
rect 268948 6322 268976 6718
rect 269026 6624 269082 6633
rect 269132 6610 269160 7142
rect 269224 6798 269252 7686
rect 269212 6792 269264 6798
rect 269212 6734 269264 6740
rect 269082 6582 269160 6610
rect 269026 6559 269082 6568
rect 269120 6452 269172 6458
rect 269120 6394 269172 6400
rect 268936 6316 268988 6322
rect 268936 6258 268988 6264
rect 268934 6216 268990 6225
rect 268844 6180 268896 6186
rect 268934 6151 268990 6160
rect 268844 6122 268896 6128
rect 268842 6080 268898 6089
rect 268842 6015 268898 6024
rect 268856 3738 268884 6015
rect 268948 5846 268976 6151
rect 269026 5944 269082 5953
rect 269026 5879 269028 5888
rect 269080 5879 269082 5888
rect 269028 5850 269080 5856
rect 268936 5840 268988 5846
rect 268936 5782 268988 5788
rect 269026 5264 269082 5273
rect 269026 5199 269082 5208
rect 268934 4856 268990 4865
rect 269040 4826 269068 5199
rect 268934 4791 268990 4800
rect 269028 4820 269080 4826
rect 268844 3732 268896 3738
rect 268844 3674 268896 3680
rect 268842 3632 268898 3641
rect 268842 3567 268898 3576
rect 268752 3528 268804 3534
rect 268752 3470 268804 3476
rect 268660 3120 268712 3126
rect 268660 3062 268712 3068
rect 268660 2984 268712 2990
rect 268660 2926 268712 2932
rect 268672 2514 268700 2926
rect 268660 2508 268712 2514
rect 268660 2450 268712 2456
rect 268856 2106 268884 3567
rect 268948 3398 268976 4791
rect 269028 4762 269080 4768
rect 269028 4548 269080 4554
rect 269028 4490 269080 4496
rect 268936 3392 268988 3398
rect 268936 3334 268988 3340
rect 269040 3058 269068 4490
rect 269132 3738 269160 6394
rect 269212 4616 269264 4622
rect 269212 4558 269264 4564
rect 269120 3732 269172 3738
rect 269120 3674 269172 3680
rect 269028 3052 269080 3058
rect 269028 2994 269080 3000
rect 269120 2440 269172 2446
rect 269120 2382 269172 2388
rect 268844 2100 268896 2106
rect 268844 2042 268896 2048
rect 268568 2032 268620 2038
rect 268568 1974 268620 1980
rect 269132 1970 269160 2382
rect 269224 2310 269252 4558
rect 269316 4146 269344 8366
rect 269580 8084 269632 8090
rect 269580 8026 269632 8032
rect 269592 7410 269620 8026
rect 269580 7404 269632 7410
rect 269580 7346 269632 7352
rect 269396 6316 269448 6322
rect 269396 6258 269448 6264
rect 269408 5370 269436 6258
rect 269580 5704 269632 5710
rect 269486 5672 269542 5681
rect 269580 5646 269632 5652
rect 269486 5607 269542 5616
rect 269396 5364 269448 5370
rect 269396 5306 269448 5312
rect 269304 4140 269356 4146
rect 269304 4082 269356 4088
rect 269500 4010 269528 5607
rect 269488 4004 269540 4010
rect 269488 3946 269540 3952
rect 269592 3194 269620 5646
rect 269684 4298 269712 8978
rect 269764 8492 269816 8498
rect 269764 8434 269816 8440
rect 269776 7410 269804 8434
rect 269868 7886 269896 9454
rect 269856 7880 269908 7886
rect 269856 7822 269908 7828
rect 269764 7404 269816 7410
rect 269764 7346 269816 7352
rect 269776 4486 269804 7346
rect 269868 6798 269896 7822
rect 269856 6792 269908 6798
rect 269856 6734 269908 6740
rect 269960 5710 269988 9590
rect 270420 9178 270448 9658
rect 270498 9616 270554 9625
rect 270498 9551 270500 9560
rect 270552 9551 270554 9560
rect 270500 9522 270552 9528
rect 272168 9489 272196 9959
rect 271970 9480 272026 9489
rect 270592 9444 270644 9450
rect 271970 9415 272026 9424
rect 272154 9480 272210 9489
rect 272154 9415 272210 9424
rect 270592 9386 270644 9392
rect 270408 9172 270460 9178
rect 270408 9114 270460 9120
rect 270408 8832 270460 8838
rect 270408 8774 270460 8780
rect 270040 8288 270092 8294
rect 270040 8230 270092 8236
rect 270052 8090 270080 8230
rect 270040 8084 270092 8090
rect 270040 8026 270092 8032
rect 270316 8016 270368 8022
rect 270316 7958 270368 7964
rect 270132 7880 270184 7886
rect 270132 7822 270184 7828
rect 270040 7744 270092 7750
rect 270040 7686 270092 7692
rect 270052 6798 270080 7686
rect 270040 6792 270092 6798
rect 270040 6734 270092 6740
rect 270144 6662 270172 7822
rect 270224 7812 270276 7818
rect 270224 7754 270276 7760
rect 270236 6866 270264 7754
rect 270328 7546 270356 7958
rect 270316 7540 270368 7546
rect 270316 7482 270368 7488
rect 270420 7478 270448 8774
rect 270500 8356 270552 8362
rect 270500 8298 270552 8304
rect 270408 7472 270460 7478
rect 270408 7414 270460 7420
rect 270512 7154 270540 8298
rect 270420 7126 270540 7154
rect 270224 6860 270276 6866
rect 270224 6802 270276 6808
rect 270132 6656 270184 6662
rect 270132 6598 270184 6604
rect 270236 6390 270264 6802
rect 270224 6384 270276 6390
rect 270224 6326 270276 6332
rect 270420 6236 270448 7126
rect 270500 6996 270552 7002
rect 270500 6938 270552 6944
rect 270512 6390 270540 6938
rect 270500 6384 270552 6390
rect 270500 6326 270552 6332
rect 270500 6248 270552 6254
rect 270314 6216 270370 6225
rect 270420 6208 270500 6236
rect 270500 6190 270552 6196
rect 270314 6151 270370 6160
rect 269948 5704 270000 5710
rect 269948 5646 270000 5652
rect 269856 5636 269908 5642
rect 269856 5578 269908 5584
rect 269868 5166 269896 5578
rect 269856 5160 269908 5166
rect 269856 5102 269908 5108
rect 269868 4622 269896 5102
rect 270328 4826 270356 6151
rect 270512 5794 270540 6190
rect 270420 5766 270540 5794
rect 270316 4820 270368 4826
rect 270316 4762 270368 4768
rect 269856 4616 269908 4622
rect 269856 4558 269908 4564
rect 270420 4486 270448 5766
rect 270498 5672 270554 5681
rect 270498 5607 270554 5616
rect 269764 4480 269816 4486
rect 269764 4422 269816 4428
rect 270408 4480 270460 4486
rect 270408 4422 270460 4428
rect 269684 4270 269988 4298
rect 269580 3188 269632 3194
rect 269580 3130 269632 3136
rect 269856 3052 269908 3058
rect 269856 2994 269908 3000
rect 269868 2650 269896 2994
rect 269856 2644 269908 2650
rect 269856 2586 269908 2592
rect 269212 2304 269264 2310
rect 269212 2246 269264 2252
rect 269960 2038 269988 4270
rect 270512 4010 270540 5607
rect 270500 4004 270552 4010
rect 270500 3946 270552 3952
rect 270604 3534 270632 9386
rect 271984 8945 272012 9415
rect 271970 8936 272026 8945
rect 270868 8900 270920 8906
rect 271970 8871 272026 8880
rect 270868 8842 270920 8848
rect 270684 8492 270736 8498
rect 270684 8434 270736 8440
rect 270696 7546 270724 8434
rect 270684 7540 270736 7546
rect 270684 7482 270736 7488
rect 270776 7268 270828 7274
rect 270776 7210 270828 7216
rect 270682 6352 270738 6361
rect 270682 6287 270738 6296
rect 270696 3738 270724 6287
rect 270788 4282 270816 7210
rect 270880 6458 270908 8842
rect 271337 8732 271645 8741
rect 271337 8730 271343 8732
rect 271399 8730 271423 8732
rect 271479 8730 271503 8732
rect 271559 8730 271583 8732
rect 271639 8730 271645 8732
rect 271399 8678 271401 8730
rect 271581 8678 271583 8730
rect 271337 8676 271343 8678
rect 271399 8676 271423 8678
rect 271479 8676 271503 8678
rect 271559 8676 271583 8678
rect 271639 8676 271645 8678
rect 271337 8667 271645 8676
rect 271786 8256 271842 8265
rect 271786 8191 271842 8200
rect 271052 8084 271104 8090
rect 271052 8026 271104 8032
rect 271144 8084 271196 8090
rect 271800 8072 271828 8191
rect 272154 8120 272210 8129
rect 271800 8044 271920 8072
rect 272154 8055 272156 8064
rect 271144 8026 271196 8032
rect 270958 6760 271014 6769
rect 270958 6695 271014 6704
rect 270868 6452 270920 6458
rect 270868 6394 270920 6400
rect 270868 6112 270920 6118
rect 270868 6054 270920 6060
rect 270776 4276 270828 4282
rect 270776 4218 270828 4224
rect 270880 4146 270908 6054
rect 270868 4140 270920 4146
rect 270868 4082 270920 4088
rect 270774 4040 270830 4049
rect 270774 3975 270830 3984
rect 270684 3732 270736 3738
rect 270684 3674 270736 3680
rect 270788 3670 270816 3975
rect 270776 3664 270828 3670
rect 270776 3606 270828 3612
rect 270592 3528 270644 3534
rect 270592 3470 270644 3476
rect 270972 3058 271000 6695
rect 271064 4622 271092 8026
rect 271156 7721 271184 8026
rect 271786 7984 271842 7993
rect 271786 7919 271842 7928
rect 271800 7721 271828 7919
rect 271142 7712 271198 7721
rect 271142 7647 271198 7656
rect 271786 7712 271842 7721
rect 271337 7644 271645 7653
rect 271786 7647 271842 7656
rect 271337 7642 271343 7644
rect 271399 7642 271423 7644
rect 271479 7642 271503 7644
rect 271559 7642 271583 7644
rect 271639 7642 271645 7644
rect 271399 7590 271401 7642
rect 271581 7590 271583 7642
rect 271337 7588 271343 7590
rect 271399 7588 271423 7590
rect 271479 7588 271503 7590
rect 271559 7588 271583 7590
rect 271639 7588 271645 7590
rect 271142 7576 271198 7585
rect 271337 7579 271645 7588
rect 271142 7511 271144 7520
rect 271196 7511 271198 7520
rect 271144 7482 271196 7488
rect 271892 7426 271920 8044
rect 272208 8055 272210 8064
rect 272156 8026 272208 8032
rect 272154 7984 272210 7993
rect 272154 7919 272210 7928
rect 272168 7546 272196 7919
rect 272156 7540 272208 7546
rect 272156 7482 272208 7488
rect 271970 7440 272026 7449
rect 271892 7398 271970 7426
rect 271970 7375 272026 7384
rect 272062 6624 272118 6633
rect 271337 6556 271645 6565
rect 272062 6559 272118 6568
rect 271337 6554 271343 6556
rect 271399 6554 271423 6556
rect 271479 6554 271503 6556
rect 271559 6554 271583 6556
rect 271639 6554 271645 6556
rect 271399 6502 271401 6554
rect 271581 6502 271583 6554
rect 271337 6500 271343 6502
rect 271399 6500 271423 6502
rect 271479 6500 271503 6502
rect 271559 6500 271583 6502
rect 271639 6500 271645 6502
rect 271142 6488 271198 6497
rect 271337 6491 271645 6500
rect 271142 6423 271198 6432
rect 271878 6488 271934 6497
rect 271878 6423 271934 6432
rect 271156 5953 271184 6423
rect 271326 6352 271382 6361
rect 271326 6287 271382 6296
rect 271340 6089 271368 6287
rect 271326 6080 271382 6089
rect 271326 6015 271382 6024
rect 271694 6080 271750 6089
rect 271694 6015 271750 6024
rect 271142 5944 271198 5953
rect 271142 5879 271198 5888
rect 271236 5636 271288 5642
rect 271236 5578 271288 5584
rect 271144 5568 271196 5574
rect 271142 5536 271144 5545
rect 271196 5536 271198 5545
rect 271142 5471 271198 5480
rect 271052 4616 271104 4622
rect 271052 4558 271104 4564
rect 271144 4616 271196 4622
rect 271144 4558 271196 4564
rect 271052 4480 271104 4486
rect 271156 4457 271184 4558
rect 271052 4422 271104 4428
rect 271142 4448 271198 4457
rect 270960 3052 271012 3058
rect 270960 2994 271012 3000
rect 270684 2848 270736 2854
rect 270682 2816 270684 2825
rect 270736 2816 270738 2825
rect 270682 2751 270738 2760
rect 270040 2440 270092 2446
rect 270040 2382 270092 2388
rect 269948 2032 270000 2038
rect 269948 1974 270000 1980
rect 267740 1964 267792 1970
rect 267740 1906 267792 1912
rect 269120 1964 269172 1970
rect 269120 1906 269172 1912
rect 268842 1864 268898 1873
rect 268842 1799 268898 1808
rect 267832 1760 267884 1766
rect 267832 1702 267884 1708
rect 268200 1760 268252 1766
rect 268200 1702 268252 1708
rect 267844 1358 267872 1702
rect 268212 1358 268240 1702
rect 268856 1494 268884 1799
rect 268844 1488 268896 1494
rect 268844 1430 268896 1436
rect 269132 1358 269160 1906
rect 269764 1760 269816 1766
rect 269764 1702 269816 1708
rect 267832 1352 267884 1358
rect 267660 1278 267780 1306
rect 268200 1352 268252 1358
rect 267832 1294 267884 1300
rect 268014 1320 268070 1329
rect 267648 1216 267700 1222
rect 267648 1158 267700 1164
rect 267660 649 267688 1158
rect 267752 785 267780 1278
rect 268200 1294 268252 1300
rect 269120 1352 269172 1358
rect 269120 1294 269172 1300
rect 268014 1255 268070 1264
rect 267924 1012 267976 1018
rect 267924 954 267976 960
rect 267936 921 267964 954
rect 268028 950 268056 1255
rect 268384 1216 268436 1222
rect 268384 1158 268436 1164
rect 268016 944 268068 950
rect 267922 912 267978 921
rect 268016 886 268068 892
rect 267922 847 267978 856
rect 267738 776 267794 785
rect 267738 711 267794 720
rect 268396 649 268424 1158
rect 269776 649 269804 1702
rect 269854 1592 269910 1601
rect 269854 1527 269856 1536
rect 269908 1527 269910 1536
rect 269856 1498 269908 1504
rect 270052 1358 270080 2382
rect 270132 2304 270184 2310
rect 270132 2246 270184 2252
rect 270776 2304 270828 2310
rect 270776 2246 270828 2252
rect 270144 1358 270172 2246
rect 270040 1352 270092 1358
rect 270040 1294 270092 1300
rect 270132 1352 270184 1358
rect 270132 1294 270184 1300
rect 270316 1216 270368 1222
rect 270316 1158 270368 1164
rect 260196 614 260248 620
rect 261114 640 261170 649
rect 258078 575 258134 584
rect 261114 575 261170 584
rect 262862 640 262918 649
rect 262862 575 262918 584
rect 263322 640 263378 649
rect 263322 575 263378 584
rect 264334 640 264390 649
rect 264334 575 264390 584
rect 264978 640 265034 649
rect 264978 575 265034 584
rect 265806 640 265862 649
rect 265806 575 265862 584
rect 266358 640 266414 649
rect 266358 575 266414 584
rect 266910 640 266966 649
rect 266910 575 266966 584
rect 267646 640 267702 649
rect 267646 575 267702 584
rect 268382 640 268438 649
rect 268382 575 268438 584
rect 269762 640 269818 649
rect 269762 575 269818 584
rect 256700 536 256752 542
rect 256700 478 256752 484
rect 256424 400 256476 406
rect 255962 368 256018 377
rect 248052 332 248104 338
rect 270328 377 270356 1158
rect 270788 649 270816 2246
rect 271064 1426 271092 4422
rect 271142 4383 271198 4392
rect 271248 3466 271276 5578
rect 271337 5468 271645 5477
rect 271337 5466 271343 5468
rect 271399 5466 271423 5468
rect 271479 5466 271503 5468
rect 271559 5466 271583 5468
rect 271639 5466 271645 5468
rect 271399 5414 271401 5466
rect 271581 5414 271583 5466
rect 271337 5412 271343 5414
rect 271399 5412 271423 5414
rect 271479 5412 271503 5414
rect 271559 5412 271583 5414
rect 271639 5412 271645 5414
rect 271337 5403 271645 5412
rect 271708 4554 271736 6015
rect 271788 5568 271840 5574
rect 271786 5536 271788 5545
rect 271840 5536 271842 5545
rect 271786 5471 271842 5480
rect 271786 5400 271842 5409
rect 271786 5335 271842 5344
rect 271800 5001 271828 5335
rect 271786 4992 271842 5001
rect 271786 4927 271842 4936
rect 271696 4548 271748 4554
rect 271696 4490 271748 4496
rect 271337 4380 271645 4389
rect 271337 4378 271343 4380
rect 271399 4378 271423 4380
rect 271479 4378 271503 4380
rect 271559 4378 271583 4380
rect 271639 4378 271645 4380
rect 271399 4326 271401 4378
rect 271581 4326 271583 4378
rect 271337 4324 271343 4326
rect 271399 4324 271423 4326
rect 271479 4324 271503 4326
rect 271559 4324 271583 4326
rect 271639 4324 271645 4326
rect 271337 4315 271645 4324
rect 271786 4312 271842 4321
rect 271708 4270 271786 4298
rect 271708 4185 271736 4270
rect 271786 4247 271842 4256
rect 271694 4176 271750 4185
rect 271694 4111 271750 4120
rect 271788 3664 271840 3670
rect 271788 3606 271840 3612
rect 271236 3460 271288 3466
rect 271236 3402 271288 3408
rect 271144 3392 271196 3398
rect 271142 3360 271144 3369
rect 271196 3360 271198 3369
rect 271142 3295 271198 3304
rect 271337 3292 271645 3301
rect 271337 3290 271343 3292
rect 271399 3290 271423 3292
rect 271479 3290 271503 3292
rect 271559 3290 271583 3292
rect 271639 3290 271645 3292
rect 271399 3238 271401 3290
rect 271581 3238 271583 3290
rect 271337 3236 271343 3238
rect 271399 3236 271423 3238
rect 271479 3236 271503 3238
rect 271559 3236 271583 3238
rect 271639 3236 271645 3238
rect 271142 3224 271198 3233
rect 271337 3227 271645 3236
rect 271800 3233 271828 3606
rect 271892 3534 271920 6423
rect 271970 4992 272026 5001
rect 271970 4927 272026 4936
rect 271984 4622 272012 4927
rect 271972 4616 272024 4622
rect 271972 4558 272024 4564
rect 272076 4146 272104 6559
rect 272156 4752 272208 4758
rect 272156 4694 272208 4700
rect 272064 4140 272116 4146
rect 272064 4082 272116 4088
rect 272168 3913 272196 4694
rect 272154 3904 272210 3913
rect 272154 3839 272210 3848
rect 272154 3632 272210 3641
rect 272154 3567 272210 3576
rect 271880 3528 271932 3534
rect 271880 3470 271932 3476
rect 272168 3398 272196 3567
rect 272156 3392 272208 3398
rect 272156 3334 272208 3340
rect 271142 3159 271198 3168
rect 271786 3224 271842 3233
rect 271786 3159 271842 3168
rect 271156 2802 271184 3159
rect 271234 2816 271290 2825
rect 271156 2774 271234 2802
rect 271234 2751 271290 2760
rect 271142 2272 271198 2281
rect 271142 2207 271198 2216
rect 271156 1834 271184 2207
rect 271337 2204 271645 2213
rect 271337 2202 271343 2204
rect 271399 2202 271423 2204
rect 271479 2202 271503 2204
rect 271559 2202 271583 2204
rect 271639 2202 271645 2204
rect 271399 2150 271401 2202
rect 271581 2150 271583 2202
rect 271337 2148 271343 2150
rect 271399 2148 271423 2150
rect 271479 2148 271503 2150
rect 271559 2148 271583 2150
rect 271639 2148 271645 2150
rect 271337 2139 271645 2148
rect 271970 2136 272026 2145
rect 271970 2071 272026 2080
rect 271144 1828 271196 1834
rect 271144 1770 271196 1776
rect 271984 1601 272012 2071
rect 272062 2000 272118 2009
rect 272062 1935 272118 1944
rect 271970 1592 272026 1601
rect 271970 1527 272026 1536
rect 271052 1420 271104 1426
rect 271052 1362 271104 1368
rect 271970 1320 272026 1329
rect 271970 1255 272026 1264
rect 271337 1116 271645 1125
rect 271337 1114 271343 1116
rect 271399 1114 271423 1116
rect 271479 1114 271503 1116
rect 271559 1114 271583 1116
rect 271639 1114 271645 1116
rect 271399 1062 271401 1114
rect 271581 1062 271583 1114
rect 271337 1060 271343 1062
rect 271399 1060 271423 1062
rect 271479 1060 271503 1062
rect 271559 1060 271583 1062
rect 271639 1060 271645 1062
rect 271337 1051 271645 1060
rect 271984 921 272012 1255
rect 271970 912 272026 921
rect 271970 847 272026 856
rect 272076 814 272104 1935
rect 272156 1828 272208 1834
rect 272156 1770 272208 1776
rect 272168 1601 272196 1770
rect 272154 1592 272210 1601
rect 272154 1527 272210 1536
rect 272064 808 272116 814
rect 272064 750 272116 756
rect 270774 640 270830 649
rect 270774 575 270830 584
rect 256424 342 256476 348
rect 270314 368 270370 377
rect 255962 303 256018 312
rect 270314 303 270370 312
rect 248052 274 248104 280
rect 244832 264 244884 270
rect 244832 206 244884 212
rect 236274 167 236330 176
rect 243728 196 243780 202
rect 243728 138 243780 144
rect 213366 96 213422 105
rect 160006 31 160062 40
rect 181996 60 182048 66
rect 149336 2 149388 8
rect 213366 31 213422 40
rect 231398 96 231454 105
rect 231398 31 231454 40
rect 181996 2 182048 8
<< via2 >>
rect 53102 10512 53158 10568
rect 1674 10104 1730 10160
rect 2410 10104 2466 10160
rect 3238 10104 3294 10160
rect 4342 10104 4398 10160
rect 5078 10104 5134 10160
rect 5814 10104 5870 10160
rect 3146 9832 3202 9888
rect 1398 9172 1454 9208
rect 1398 9152 1400 9172
rect 1400 9152 1452 9172
rect 1452 9152 1454 9172
rect 6826 10104 6882 10160
rect 7562 10104 7618 10160
rect 8390 10104 8446 10160
rect 9586 10104 9642 10160
rect 10230 10104 10286 10160
rect 10966 10104 11022 10160
rect 11978 10104 12034 10160
rect 12714 10104 12770 10160
rect 13726 10104 13782 10160
rect 14646 10104 14702 10160
rect 15382 10104 15438 10160
rect 16118 10104 16174 10160
rect 17130 10104 17186 10160
rect 17866 10104 17922 10160
rect 18602 10104 18658 10160
rect 8206 9832 8262 9888
rect 13450 9832 13506 9888
rect 19246 6860 19302 6896
rect 19246 6840 19248 6860
rect 19248 6840 19300 6860
rect 19300 6840 19302 6860
rect 21362 8628 21418 8664
rect 22098 8880 22154 8936
rect 21362 8608 21364 8628
rect 21364 8608 21416 8628
rect 21416 8608 21418 8628
rect 21914 8336 21970 8392
rect 19338 5208 19394 5264
rect 846 2760 902 2816
rect 4802 2508 4858 2544
rect 4802 2488 4804 2508
rect 4804 2488 4856 2508
rect 4856 2488 4858 2508
rect 1674 992 1730 1048
rect 1950 584 2006 640
rect 4526 1264 4582 1320
rect 3790 992 3846 1048
rect 5170 992 5226 1048
rect 2962 720 3018 776
rect 5354 720 5410 776
rect 6734 1264 6790 1320
rect 15106 3440 15162 3496
rect 14370 3168 14426 3224
rect 8666 1964 8722 2000
rect 8666 1944 8668 1964
rect 8668 1944 8720 1964
rect 8720 1944 8722 1964
rect 7102 992 7158 1048
rect 7746 448 7802 504
rect 9678 992 9734 1048
rect 11978 992 12034 1048
rect 12714 992 12770 1048
rect 10322 720 10378 776
rect 11702 720 11758 776
rect 13450 584 13506 640
rect 14094 992 14150 1048
rect 14830 1264 14886 1320
rect 19246 2760 19302 2816
rect 23202 9832 23258 9888
rect 15474 992 15530 1048
rect 15658 720 15714 776
rect 22006 1708 22008 1728
rect 22008 1708 22060 1728
rect 22060 1708 22062 1728
rect 22006 1672 22062 1708
rect 20718 1556 20774 1592
rect 20718 1536 20720 1556
rect 20720 1536 20772 1556
rect 20772 1536 20774 1556
rect 22374 1400 22430 1456
rect 22926 8336 22982 8392
rect 22834 2760 22890 2816
rect 23110 2080 23166 2136
rect 23662 8336 23718 8392
rect 23938 9172 23994 9208
rect 23938 9152 23940 9172
rect 23940 9152 23992 9172
rect 23992 9152 23994 9172
rect 23754 1420 23810 1456
rect 23754 1400 23756 1420
rect 23756 1400 23808 1420
rect 23808 1400 23810 1420
rect 25870 9716 25926 9752
rect 25870 9696 25872 9716
rect 25872 9696 25924 9716
rect 25924 9696 25926 9716
rect 27342 9716 27398 9752
rect 27342 9696 27344 9716
rect 27344 9696 27396 9716
rect 27396 9696 27398 9716
rect 25042 2760 25098 2816
rect 25226 8336 25282 8392
rect 23570 1264 23626 1320
rect 23846 1264 23902 1320
rect 25778 1264 25834 1320
rect 27434 8628 27490 8664
rect 27434 8608 27436 8628
rect 27436 8608 27488 8628
rect 27488 8608 27490 8628
rect 29090 9716 29146 9752
rect 29090 9696 29092 9716
rect 29092 9696 29144 9716
rect 29144 9696 29146 9716
rect 27526 2760 27582 2816
rect 28170 8628 28226 8664
rect 28170 8608 28172 8628
rect 28172 8608 28224 8628
rect 28224 8608 28226 8628
rect 28906 8628 28962 8664
rect 28906 8608 28908 8628
rect 28908 8608 28960 8628
rect 28960 8608 28962 8628
rect 32494 10240 32550 10296
rect 35162 10240 35218 10296
rect 35622 10240 35678 10296
rect 36266 10240 36322 10296
rect 36910 10240 36966 10296
rect 38106 10240 38162 10296
rect 38842 10240 38898 10296
rect 39486 10240 39542 10296
rect 40314 10240 40370 10296
rect 40774 10240 40830 10296
rect 41418 10240 41474 10296
rect 42062 10240 42118 10296
rect 43258 10240 43314 10296
rect 43994 10240 44050 10296
rect 44638 10240 44694 10296
rect 45466 10240 45522 10296
rect 45926 10240 45982 10296
rect 46570 10240 46626 10296
rect 47214 10240 47270 10296
rect 48226 10240 48282 10296
rect 49146 10240 49202 10296
rect 49790 10240 49846 10296
rect 50618 10240 50674 10296
rect 51354 10240 51410 10296
rect 52090 10240 52146 10296
rect 30286 9716 30342 9752
rect 30286 9696 30288 9716
rect 30288 9696 30340 9716
rect 30340 9696 30342 9716
rect 26514 1264 26570 1320
rect 17866 992 17922 1048
rect 17038 720 17094 776
rect 34754 9274 34810 9276
rect 34834 9274 34890 9276
rect 34914 9274 34970 9276
rect 34994 9274 35050 9276
rect 34754 9222 34800 9274
rect 34800 9222 34810 9274
rect 34834 9222 34864 9274
rect 34864 9222 34876 9274
rect 34876 9222 34890 9274
rect 34914 9222 34928 9274
rect 34928 9222 34940 9274
rect 34940 9222 34970 9274
rect 34994 9222 35004 9274
rect 35004 9222 35050 9274
rect 34754 9220 34810 9222
rect 34834 9220 34890 9222
rect 34914 9220 34970 9222
rect 34994 9220 35050 9222
rect 33046 9172 33102 9208
rect 33046 9152 33048 9172
rect 33048 9152 33100 9172
rect 33100 9152 33102 9172
rect 31022 8628 31078 8664
rect 31022 8608 31024 8628
rect 31024 8608 31076 8628
rect 31076 8608 31078 8628
rect 34754 8186 34810 8188
rect 34834 8186 34890 8188
rect 34914 8186 34970 8188
rect 34994 8186 35050 8188
rect 34754 8134 34800 8186
rect 34800 8134 34810 8186
rect 34834 8134 34864 8186
rect 34864 8134 34876 8186
rect 34876 8134 34890 8186
rect 34914 8134 34928 8186
rect 34928 8134 34940 8186
rect 34940 8134 34970 8186
rect 34994 8134 35004 8186
rect 35004 8134 35050 8186
rect 34754 8132 34810 8134
rect 34834 8132 34890 8134
rect 34914 8132 34970 8134
rect 34994 8132 35050 8134
rect 34754 7098 34810 7100
rect 34834 7098 34890 7100
rect 34914 7098 34970 7100
rect 34994 7098 35050 7100
rect 34754 7046 34800 7098
rect 34800 7046 34810 7098
rect 34834 7046 34864 7098
rect 34864 7046 34876 7098
rect 34876 7046 34890 7098
rect 34914 7046 34928 7098
rect 34928 7046 34940 7098
rect 34940 7046 34970 7098
rect 34994 7046 35004 7098
rect 35004 7046 35050 7098
rect 34754 7044 34810 7046
rect 34834 7044 34890 7046
rect 34914 7044 34970 7046
rect 34994 7044 35050 7046
rect 34754 6010 34810 6012
rect 34834 6010 34890 6012
rect 34914 6010 34970 6012
rect 34994 6010 35050 6012
rect 34754 5958 34800 6010
rect 34800 5958 34810 6010
rect 34834 5958 34864 6010
rect 34864 5958 34876 6010
rect 34876 5958 34890 6010
rect 34914 5958 34928 6010
rect 34928 5958 34940 6010
rect 34940 5958 34970 6010
rect 34994 5958 35004 6010
rect 35004 5958 35050 6010
rect 34754 5956 34810 5958
rect 34834 5956 34890 5958
rect 34914 5956 34970 5958
rect 34994 5956 35050 5958
rect 34754 4922 34810 4924
rect 34834 4922 34890 4924
rect 34914 4922 34970 4924
rect 34994 4922 35050 4924
rect 34754 4870 34800 4922
rect 34800 4870 34810 4922
rect 34834 4870 34864 4922
rect 34864 4870 34876 4922
rect 34876 4870 34890 4922
rect 34914 4870 34928 4922
rect 34928 4870 34940 4922
rect 34940 4870 34970 4922
rect 34994 4870 35004 4922
rect 35004 4870 35050 4922
rect 34754 4868 34810 4870
rect 34834 4868 34890 4870
rect 34914 4868 34970 4870
rect 34994 4868 35050 4870
rect 34754 3834 34810 3836
rect 34834 3834 34890 3836
rect 34914 3834 34970 3836
rect 34994 3834 35050 3836
rect 34754 3782 34800 3834
rect 34800 3782 34810 3834
rect 34834 3782 34864 3834
rect 34864 3782 34876 3834
rect 34876 3782 34890 3834
rect 34914 3782 34928 3834
rect 34928 3782 34940 3834
rect 34940 3782 34970 3834
rect 34994 3782 35004 3834
rect 35004 3782 35050 3834
rect 34754 3780 34810 3782
rect 34834 3780 34890 3782
rect 34914 3780 34970 3782
rect 34994 3780 35050 3782
rect 32770 3032 32826 3088
rect 34754 2746 34810 2748
rect 34834 2746 34890 2748
rect 34914 2746 34970 2748
rect 34994 2746 35050 2748
rect 34754 2694 34800 2746
rect 34800 2694 34810 2746
rect 34834 2694 34864 2746
rect 34864 2694 34876 2746
rect 34876 2694 34890 2746
rect 34914 2694 34928 2746
rect 34928 2694 34940 2746
rect 34940 2694 34970 2746
rect 34994 2694 35004 2746
rect 35004 2694 35050 2746
rect 34754 2692 34810 2694
rect 34834 2692 34890 2694
rect 34914 2692 34970 2694
rect 34994 2692 35050 2694
rect 34754 1658 34810 1660
rect 34834 1658 34890 1660
rect 34914 1658 34970 1660
rect 34994 1658 35050 1660
rect 34754 1606 34800 1658
rect 34800 1606 34810 1658
rect 34834 1606 34864 1658
rect 34864 1606 34876 1658
rect 34876 1606 34890 1658
rect 34914 1606 34928 1658
rect 34928 1606 34940 1658
rect 34940 1606 34970 1658
rect 34994 1606 35004 1658
rect 35004 1606 35050 1658
rect 34754 1604 34810 1606
rect 34834 1604 34890 1606
rect 34914 1604 34970 1606
rect 34994 1604 35050 1606
rect 33138 1536 33194 1592
rect 21454 584 21510 640
rect 28170 584 28226 640
rect 8390 312 8446 368
rect 18602 312 18658 368
rect 28814 312 28870 368
rect 29918 1128 29974 1184
rect 36266 5244 36268 5264
rect 36268 5244 36320 5264
rect 36320 5244 36322 5264
rect 36266 5208 36322 5244
rect 36818 4972 36820 4992
rect 36820 4972 36872 4992
rect 36872 4972 36874 4992
rect 36818 4936 36874 4972
rect 30286 584 30342 640
rect 31206 584 31262 640
rect 32494 584 32550 640
rect 35162 584 35218 640
rect 35622 584 35678 640
rect 36266 584 36322 640
rect 36910 584 36966 640
rect 38934 4004 38990 4040
rect 38934 3984 38936 4004
rect 38936 3984 38988 4004
rect 38988 3984 38990 4004
rect 38750 2488 38806 2544
rect 38106 584 38162 640
rect 38566 584 38622 640
rect 39946 584 40002 640
rect 39854 448 39910 504
rect 42614 5072 42670 5128
rect 42798 5888 42854 5944
rect 40406 1708 40408 1728
rect 40408 1708 40460 1728
rect 40460 1708 40462 1728
rect 40406 1672 40462 1708
rect 40774 584 40830 640
rect 42614 4140 42670 4176
rect 42614 4120 42616 4140
rect 42616 4120 42668 4140
rect 42668 4120 42670 4140
rect 42062 2896 42118 2952
rect 43534 4528 43590 4584
rect 43350 1944 43406 2000
rect 53286 10240 53342 10296
rect 53838 10240 53894 10296
rect 54850 10240 54906 10296
rect 55678 10240 55734 10296
rect 56506 10240 56562 10296
rect 57334 10240 57390 10296
rect 57794 10240 57850 10296
rect 46662 5072 46718 5128
rect 47122 5092 47178 5128
rect 47122 5072 47124 5092
rect 47124 5072 47176 5092
rect 47176 5072 47178 5092
rect 45742 720 45798 776
rect 47122 4120 47178 4176
rect 47582 3304 47638 3360
rect 41418 584 41474 640
rect 42062 584 42118 640
rect 43258 584 43314 640
rect 43994 584 44050 640
rect 44638 584 44694 640
rect 45466 584 45522 640
rect 45926 584 45982 640
rect 46570 584 46626 640
rect 47214 584 47270 640
rect 48226 3304 48282 3360
rect 48778 3576 48834 3632
rect 49330 3440 49386 3496
rect 49054 3168 49110 3224
rect 49238 2916 49294 2952
rect 49238 2896 49240 2916
rect 49240 2896 49292 2916
rect 49292 2896 49294 2916
rect 51630 3596 51686 3632
rect 51630 3576 51632 3596
rect 51632 3576 51684 3596
rect 51684 3576 51686 3596
rect 48226 584 48282 640
rect 49146 584 49202 640
rect 49790 584 49846 640
rect 50618 584 50674 640
rect 51354 584 51410 640
rect 52182 7928 52238 7984
rect 51814 3440 51870 3496
rect 53746 6180 53802 6216
rect 53746 6160 53748 6180
rect 53748 6160 53800 6180
rect 53800 6160 53802 6180
rect 53286 5616 53342 5672
rect 52090 2760 52146 2816
rect 53286 2080 53342 2136
rect 54298 1420 54354 1456
rect 54298 1400 54300 1420
rect 54300 1400 54352 1420
rect 54352 1400 54354 1420
rect 52090 584 52146 640
rect 52918 584 52974 640
rect 38842 312 38898 368
rect 55126 2760 55182 2816
rect 58806 10240 58862 10296
rect 59266 10240 59322 10296
rect 60278 10240 60334 10296
rect 57978 1536 58034 1592
rect 54482 584 54538 640
rect 61014 10240 61070 10296
rect 61750 10240 61806 10296
rect 62486 10240 62542 10296
rect 59358 1536 59414 1592
rect 59542 1536 59598 1592
rect 63406 10240 63462 10296
rect 63958 10240 64014 10296
rect 64694 10240 64750 10296
rect 65522 10240 65578 10296
rect 65890 10240 65946 10296
rect 67178 10240 67234 10296
rect 68552 9818 68608 9820
rect 68632 9818 68688 9820
rect 68712 9818 68768 9820
rect 68792 9818 68848 9820
rect 68552 9766 68598 9818
rect 68598 9766 68608 9818
rect 68632 9766 68662 9818
rect 68662 9766 68674 9818
rect 68674 9766 68688 9818
rect 68712 9766 68726 9818
rect 68726 9766 68738 9818
rect 68738 9766 68768 9818
rect 68792 9766 68802 9818
rect 68802 9766 68848 9818
rect 68552 9764 68608 9766
rect 68632 9764 68688 9766
rect 68712 9764 68768 9766
rect 68792 9764 68848 9766
rect 69110 9580 69166 9616
rect 69110 9560 69112 9580
rect 69112 9560 69164 9580
rect 69164 9560 69166 9580
rect 81622 10512 81678 10568
rect 82634 10512 82690 10568
rect 86774 10512 86830 10568
rect 72054 10376 72110 10432
rect 71502 10104 71558 10160
rect 70030 9832 70086 9888
rect 70306 9580 70362 9616
rect 70306 9560 70308 9580
rect 70308 9560 70360 9580
rect 70360 9560 70362 9580
rect 72146 9580 72202 9616
rect 72146 9560 72148 9580
rect 72148 9560 72200 9580
rect 72200 9560 72202 9580
rect 74262 9560 74318 9616
rect 73434 9036 73490 9072
rect 73434 9016 73436 9036
rect 73436 9016 73488 9036
rect 73488 9016 73490 9036
rect 68552 8730 68608 8732
rect 68632 8730 68688 8732
rect 68712 8730 68768 8732
rect 68792 8730 68848 8732
rect 68552 8678 68598 8730
rect 68598 8678 68608 8730
rect 68632 8678 68662 8730
rect 68662 8678 68674 8730
rect 68674 8678 68688 8730
rect 68712 8678 68726 8730
rect 68726 8678 68738 8730
rect 68738 8678 68768 8730
rect 68792 8678 68802 8730
rect 68802 8678 68848 8730
rect 68552 8676 68608 8678
rect 68632 8676 68688 8678
rect 68712 8676 68768 8678
rect 68792 8676 68848 8678
rect 68552 7642 68608 7644
rect 68632 7642 68688 7644
rect 68712 7642 68768 7644
rect 68792 7642 68848 7644
rect 68552 7590 68598 7642
rect 68598 7590 68608 7642
rect 68632 7590 68662 7642
rect 68662 7590 68674 7642
rect 68674 7590 68688 7642
rect 68712 7590 68726 7642
rect 68726 7590 68738 7642
rect 68738 7590 68768 7642
rect 68792 7590 68802 7642
rect 68802 7590 68848 7642
rect 68552 7588 68608 7590
rect 68632 7588 68688 7590
rect 68712 7588 68768 7590
rect 68792 7588 68848 7590
rect 65062 2352 65118 2408
rect 55678 448 55734 504
rect 56414 448 56470 504
rect 57150 448 57206 504
rect 58254 448 58310 504
rect 60002 448 60058 504
rect 60922 448 60978 504
rect 61474 448 61530 504
rect 62394 448 62450 504
rect 63130 448 63186 504
rect 65890 448 65946 504
rect 68552 6554 68608 6556
rect 68632 6554 68688 6556
rect 68712 6554 68768 6556
rect 68792 6554 68848 6556
rect 68552 6502 68598 6554
rect 68598 6502 68608 6554
rect 68632 6502 68662 6554
rect 68662 6502 68674 6554
rect 68674 6502 68688 6554
rect 68712 6502 68726 6554
rect 68726 6502 68738 6554
rect 68738 6502 68768 6554
rect 68792 6502 68802 6554
rect 68802 6502 68848 6554
rect 68552 6500 68608 6502
rect 68632 6500 68688 6502
rect 68712 6500 68768 6502
rect 68792 6500 68848 6502
rect 79230 10104 79286 10160
rect 77206 9832 77262 9888
rect 78678 9832 78734 9888
rect 74722 9580 74778 9616
rect 74722 9560 74724 9580
rect 74724 9560 74776 9580
rect 74776 9560 74778 9580
rect 74722 9016 74778 9072
rect 75826 7656 75882 7712
rect 76470 9560 76526 9616
rect 77298 9580 77354 9616
rect 77298 9560 77300 9580
rect 77300 9560 77352 9580
rect 77352 9560 77354 9580
rect 76562 7404 76618 7440
rect 76562 7384 76564 7404
rect 76564 7384 76616 7404
rect 76616 7384 76618 7404
rect 79966 9580 80022 9616
rect 79966 9560 79968 9580
rect 79968 9560 80020 9580
rect 80020 9560 80022 9580
rect 78770 7248 78826 7304
rect 81254 9832 81310 9888
rect 83094 10104 83150 10160
rect 83922 10104 83978 10160
rect 84658 10104 84714 10160
rect 85394 10104 85450 10160
rect 80150 7520 80206 7576
rect 86406 9832 86462 9888
rect 82726 6568 82782 6624
rect 90362 10240 90418 10296
rect 88246 9172 88302 9208
rect 88246 9152 88248 9172
rect 88248 9152 88300 9172
rect 88300 9152 88302 9172
rect 87510 8628 87566 8664
rect 87510 8608 87512 8628
rect 87512 8608 87564 8628
rect 87564 8608 87566 8628
rect 85486 7792 85542 7848
rect 84106 6432 84162 6488
rect 78954 6296 79010 6352
rect 68552 5466 68608 5468
rect 68632 5466 68688 5468
rect 68712 5466 68768 5468
rect 68792 5466 68848 5468
rect 68552 5414 68598 5466
rect 68598 5414 68608 5466
rect 68632 5414 68662 5466
rect 68662 5414 68674 5466
rect 68674 5414 68688 5466
rect 68712 5414 68726 5466
rect 68726 5414 68738 5466
rect 68738 5414 68768 5466
rect 68792 5414 68802 5466
rect 68802 5414 68848 5466
rect 68552 5412 68608 5414
rect 68632 5412 68688 5414
rect 68712 5412 68768 5414
rect 68792 5412 68848 5414
rect 80058 4392 80114 4448
rect 68552 4378 68608 4380
rect 68632 4378 68688 4380
rect 68712 4378 68768 4380
rect 68792 4378 68848 4380
rect 68552 4326 68598 4378
rect 68598 4326 68608 4378
rect 68632 4326 68662 4378
rect 68662 4326 68674 4378
rect 68674 4326 68688 4378
rect 68712 4326 68726 4378
rect 68726 4326 68738 4378
rect 68738 4326 68768 4378
rect 68792 4326 68802 4378
rect 68802 4326 68848 4378
rect 68552 4324 68608 4326
rect 68632 4324 68688 4326
rect 68712 4324 68768 4326
rect 68792 4324 68848 4326
rect 78586 3576 78642 3632
rect 68552 3290 68608 3292
rect 68632 3290 68688 3292
rect 68712 3290 68768 3292
rect 68792 3290 68848 3292
rect 68552 3238 68598 3290
rect 68598 3238 68608 3290
rect 68632 3238 68662 3290
rect 68662 3238 68674 3290
rect 68674 3238 68688 3290
rect 68712 3238 68726 3290
rect 68726 3238 68738 3290
rect 68738 3238 68768 3290
rect 68792 3238 68802 3290
rect 68802 3238 68848 3290
rect 68552 3236 68608 3238
rect 68632 3236 68688 3238
rect 68712 3236 68768 3238
rect 68792 3236 68848 3238
rect 67638 3032 67694 3088
rect 68552 2202 68608 2204
rect 68632 2202 68688 2204
rect 68712 2202 68768 2204
rect 68792 2202 68848 2204
rect 68552 2150 68598 2202
rect 68598 2150 68608 2202
rect 68632 2150 68662 2202
rect 68662 2150 68674 2202
rect 68674 2150 68688 2202
rect 68712 2150 68726 2202
rect 68726 2150 68738 2202
rect 68738 2150 68768 2202
rect 68792 2150 68802 2202
rect 68802 2150 68848 2202
rect 68552 2148 68608 2150
rect 68632 2148 68688 2150
rect 68712 2148 68768 2150
rect 68792 2148 68848 2150
rect 68552 1114 68608 1116
rect 68632 1114 68688 1116
rect 68712 1114 68768 1116
rect 68792 1114 68848 1116
rect 68552 1062 68598 1114
rect 68598 1062 68608 1114
rect 68632 1062 68662 1114
rect 68662 1062 68674 1114
rect 68674 1062 68688 1114
rect 68712 1062 68726 1114
rect 68726 1062 68738 1114
rect 68738 1062 68768 1114
rect 68792 1062 68802 1114
rect 68802 1062 68848 1114
rect 68552 1060 68608 1062
rect 68632 1060 68688 1062
rect 68712 1060 68768 1062
rect 68792 1060 68848 1062
rect 72054 1828 72110 1864
rect 72054 1808 72056 1828
rect 72056 1808 72108 1828
rect 72108 1808 72110 1828
rect 71502 992 71558 1048
rect 72238 992 72294 1048
rect 69110 856 69166 912
rect 69570 856 69626 912
rect 70950 856 71006 912
rect 74630 1828 74686 1864
rect 74630 1808 74632 1828
rect 74632 1808 74684 1828
rect 74684 1808 74686 1828
rect 73710 992 73766 1048
rect 72974 856 73030 912
rect 67270 448 67326 504
rect 76470 1264 76526 1320
rect 75734 992 75790 1048
rect 77206 992 77262 1048
rect 74262 856 74318 912
rect 74722 856 74778 912
rect 77298 856 77354 912
rect 78678 1264 78734 1320
rect 79414 992 79470 1048
rect 79966 856 80022 912
rect 84106 3304 84162 3360
rect 81622 1264 81678 1320
rect 80886 992 80942 1048
rect 82358 992 82414 1048
rect 82634 856 82690 912
rect 83830 1264 83886 1320
rect 84842 1964 84898 2000
rect 89350 9444 89406 9480
rect 89350 9424 89352 9444
rect 89352 9424 89404 9444
rect 89404 9424 89406 9444
rect 88982 2488 89038 2544
rect 84842 1944 84844 1964
rect 84844 1944 84896 1964
rect 84896 1944 84898 1964
rect 84566 992 84622 1048
rect 86038 992 86094 1048
rect 88338 1400 88394 1456
rect 89074 1420 89130 1456
rect 89074 1400 89076 1420
rect 89076 1400 89128 1420
rect 89128 1400 89130 1420
rect 89718 8064 89774 8120
rect 89626 2080 89682 2136
rect 90822 8628 90878 8664
rect 90822 8608 90824 8628
rect 90824 8608 90876 8628
rect 90876 8608 90878 8628
rect 91650 9968 91706 10024
rect 89534 1264 89590 1320
rect 90178 1264 90234 1320
rect 92018 9444 92074 9480
rect 92018 9424 92020 9444
rect 92020 9424 92072 9444
rect 92072 9424 92074 9444
rect 91742 9172 91798 9208
rect 91742 9152 91744 9172
rect 91744 9152 91796 9172
rect 91796 9152 91798 9172
rect 92754 9716 92810 9752
rect 92754 9696 92756 9716
rect 92756 9696 92808 9716
rect 92808 9696 92810 9716
rect 91190 2352 91246 2408
rect 92478 6976 92534 7032
rect 91190 1536 91246 1592
rect 91374 1536 91430 1592
rect 90822 1264 90878 1320
rect 92018 1264 92074 1320
rect 86774 856 86830 912
rect 88522 1128 88578 1184
rect 92202 584 92258 640
rect 87510 448 87566 504
rect 53102 312 53158 368
rect 63866 312 63922 368
rect 64602 312 64658 368
rect 65982 312 66038 368
rect 85026 312 85082 368
rect 85486 312 85542 368
rect 92662 4256 92718 4312
rect 92570 3732 92626 3768
rect 92570 3712 92572 3732
rect 92572 3712 92624 3732
rect 92624 3712 92626 3732
rect 92754 4120 92810 4176
rect 92938 3984 92994 4040
rect 92386 1672 92442 1728
rect 92754 1264 92810 1320
rect 92386 856 92442 912
rect 93490 9716 93546 9752
rect 93490 9696 93492 9716
rect 93492 9696 93544 9716
rect 93544 9696 93546 9716
rect 94318 8064 94374 8120
rect 94318 7656 94374 7712
rect 94594 8628 94650 8664
rect 94594 8608 94596 8628
rect 94596 8608 94648 8628
rect 94648 8608 94650 8628
rect 94226 6840 94282 6896
rect 93950 3032 94006 3088
rect 93674 2216 93730 2272
rect 93674 1808 93730 1864
rect 94502 7520 94558 7576
rect 94502 7112 94558 7168
rect 95054 8628 95110 8664
rect 95054 8608 95056 8628
rect 95056 8608 95108 8628
rect 95108 8608 95110 8628
rect 95238 8472 95294 8528
rect 94502 6296 94558 6352
rect 94502 5752 94558 5808
rect 94410 5516 94412 5536
rect 94412 5516 94464 5536
rect 94464 5516 94466 5536
rect 94410 5480 94466 5516
rect 94226 2080 94282 2136
rect 93030 992 93086 1048
rect 92478 584 92534 640
rect 94410 2624 94466 2680
rect 94870 3168 94926 3224
rect 94594 992 94650 1048
rect 95054 6024 95110 6080
rect 95238 3712 95294 3768
rect 95238 3168 95294 3224
rect 95054 1844 95056 1864
rect 95056 1844 95108 1864
rect 95108 1844 95110 1864
rect 95514 4120 95570 4176
rect 95422 2760 95478 2816
rect 95330 2080 95386 2136
rect 95054 1808 95110 1844
rect 95238 1808 95294 1864
rect 95330 1536 95386 1592
rect 96066 9716 96122 9752
rect 96066 9696 96068 9716
rect 96068 9696 96120 9716
rect 96120 9696 96122 9716
rect 96342 9716 96398 9752
rect 96342 9696 96344 9716
rect 96344 9696 96396 9716
rect 96396 9696 96398 9716
rect 95882 8492 95938 8528
rect 95882 8472 95884 8492
rect 95884 8472 95936 8492
rect 95936 8472 95938 8492
rect 95974 8200 96030 8256
rect 96066 5480 96122 5536
rect 96158 3032 96214 3088
rect 96618 10412 96620 10432
rect 96620 10412 96672 10432
rect 96672 10412 96674 10432
rect 96618 10376 96674 10412
rect 96526 8880 96582 8936
rect 96986 9016 97042 9072
rect 98550 8916 98552 8936
rect 98552 8916 98604 8936
rect 98604 8916 98606 8936
rect 97170 8508 97172 8528
rect 97172 8508 97224 8528
rect 97224 8508 97226 8528
rect 97170 8472 97226 8508
rect 97538 8628 97594 8664
rect 97538 8608 97540 8628
rect 97540 8608 97592 8628
rect 97592 8608 97594 8628
rect 97998 8628 98054 8664
rect 97998 8608 98000 8628
rect 98000 8608 98052 8628
rect 98052 8608 98054 8628
rect 98550 8880 98606 8916
rect 96618 7792 96674 7848
rect 96618 4936 96674 4992
rect 96526 4392 96582 4448
rect 96618 3848 96674 3904
rect 95974 2216 96030 2272
rect 96434 2352 96490 2408
rect 96434 2100 96490 2136
rect 96434 2080 96436 2100
rect 96436 2080 96488 2100
rect 96488 2080 96490 2100
rect 96250 1536 96306 1592
rect 97446 6840 97502 6896
rect 97538 5344 97594 5400
rect 97630 3984 97686 4040
rect 97538 3712 97594 3768
rect 97906 6876 97908 6896
rect 97908 6876 97960 6896
rect 97960 6876 97962 6896
rect 97906 6840 97962 6876
rect 98458 5344 98514 5400
rect 99378 9716 99434 9752
rect 99378 9696 99380 9716
rect 99380 9696 99432 9716
rect 99432 9696 99434 9716
rect 99286 9036 99342 9072
rect 99286 9016 99288 9036
rect 99288 9016 99340 9036
rect 99340 9016 99342 9036
rect 99470 8880 99526 8936
rect 99378 8628 99434 8664
rect 99378 8608 99380 8628
rect 99380 8608 99432 8628
rect 99432 8608 99434 8628
rect 98918 8472 98974 8528
rect 96986 2796 96988 2816
rect 96988 2796 97040 2816
rect 97040 2796 97042 2816
rect 96986 2760 97042 2796
rect 96894 2352 96950 2408
rect 96802 1672 96858 1728
rect 96986 1672 97042 1728
rect 94778 584 94834 640
rect 97722 2624 97778 2680
rect 97814 2080 97870 2136
rect 97998 1672 98054 1728
rect 97906 1536 97962 1592
rect 94318 176 94374 232
rect 99102 8336 99158 8392
rect 99102 6432 99158 6488
rect 99470 4820 99526 4856
rect 99470 4800 99472 4820
rect 99472 4800 99524 4820
rect 99524 4800 99526 4820
rect 99838 4392 99894 4448
rect 100482 9716 100538 9752
rect 100482 9696 100484 9716
rect 100484 9696 100536 9716
rect 100536 9696 100538 9716
rect 100298 8508 100300 8528
rect 100300 8508 100352 8528
rect 100352 8508 100354 8528
rect 100298 8472 100354 8508
rect 103242 10240 103298 10296
rect 103886 10240 103942 10296
rect 104714 10240 104770 10296
rect 100666 8336 100722 8392
rect 100666 6976 100722 7032
rect 100482 6432 100538 6488
rect 100206 6160 100262 6216
rect 100022 4800 100078 4856
rect 100022 4528 100078 4584
rect 100298 5636 100354 5672
rect 100298 5616 100300 5636
rect 100300 5616 100352 5636
rect 100352 5616 100354 5636
rect 101218 9172 101274 9208
rect 101218 9152 101220 9172
rect 101220 9152 101272 9172
rect 101272 9152 101274 9172
rect 102351 9274 102407 9276
rect 102431 9274 102487 9276
rect 102511 9274 102567 9276
rect 102591 9274 102647 9276
rect 102351 9222 102397 9274
rect 102397 9222 102407 9274
rect 102431 9222 102461 9274
rect 102461 9222 102473 9274
rect 102473 9222 102487 9274
rect 102511 9222 102525 9274
rect 102525 9222 102537 9274
rect 102537 9222 102567 9274
rect 102591 9222 102601 9274
rect 102601 9222 102647 9274
rect 102351 9220 102407 9222
rect 102431 9220 102487 9222
rect 102511 9220 102567 9222
rect 102591 9220 102647 9222
rect 102046 8200 102102 8256
rect 102351 8186 102407 8188
rect 102431 8186 102487 8188
rect 102511 8186 102567 8188
rect 102591 8186 102647 8188
rect 102351 8134 102397 8186
rect 102397 8134 102407 8186
rect 102431 8134 102461 8186
rect 102461 8134 102473 8186
rect 102473 8134 102487 8186
rect 102511 8134 102525 8186
rect 102525 8134 102537 8186
rect 102537 8134 102567 8186
rect 102591 8134 102601 8186
rect 102601 8134 102647 8186
rect 102351 8132 102407 8134
rect 102431 8132 102487 8134
rect 102511 8132 102567 8134
rect 102591 8132 102647 8134
rect 102874 7656 102930 7712
rect 100666 4664 100722 4720
rect 100298 3984 100354 4040
rect 100850 5888 100906 5944
rect 100298 3440 100354 3496
rect 100482 3440 100538 3496
rect 100482 3168 100538 3224
rect 100758 3168 100814 3224
rect 99194 1264 99250 1320
rect 99286 584 99342 640
rect 101034 3168 101090 3224
rect 101310 6160 101366 6216
rect 101310 5616 101366 5672
rect 102138 7112 102194 7168
rect 102351 7098 102407 7100
rect 102431 7098 102487 7100
rect 102511 7098 102567 7100
rect 102591 7098 102647 7100
rect 102351 7046 102397 7098
rect 102397 7046 102407 7098
rect 102431 7046 102461 7098
rect 102461 7046 102473 7098
rect 102473 7046 102487 7098
rect 102511 7046 102525 7098
rect 102525 7046 102537 7098
rect 102537 7046 102567 7098
rect 102591 7046 102601 7098
rect 102601 7046 102647 7098
rect 102351 7044 102407 7046
rect 102431 7044 102487 7046
rect 102511 7044 102567 7046
rect 102591 7044 102647 7046
rect 101494 5888 101550 5944
rect 101218 3168 101274 3224
rect 101770 6704 101826 6760
rect 102690 6740 102692 6760
rect 102692 6740 102744 6760
rect 102744 6740 102746 6760
rect 102690 6704 102746 6740
rect 101954 6024 102010 6080
rect 102046 5888 102102 5944
rect 101678 5616 101734 5672
rect 102046 4256 102102 4312
rect 102351 6010 102407 6012
rect 102431 6010 102487 6012
rect 102511 6010 102567 6012
rect 102591 6010 102647 6012
rect 102351 5958 102397 6010
rect 102397 5958 102407 6010
rect 102431 5958 102461 6010
rect 102461 5958 102473 6010
rect 102473 5958 102487 6010
rect 102511 5958 102525 6010
rect 102525 5958 102537 6010
rect 102537 5958 102567 6010
rect 102591 5958 102601 6010
rect 102601 5958 102647 6010
rect 102351 5956 102407 5958
rect 102431 5956 102487 5958
rect 102511 5956 102567 5958
rect 102591 5956 102647 5958
rect 102351 4922 102407 4924
rect 102431 4922 102487 4924
rect 102511 4922 102567 4924
rect 102591 4922 102647 4924
rect 102351 4870 102397 4922
rect 102397 4870 102407 4922
rect 102431 4870 102461 4922
rect 102461 4870 102473 4922
rect 102473 4870 102487 4922
rect 102511 4870 102525 4922
rect 102525 4870 102537 4922
rect 102537 4870 102567 4922
rect 102591 4870 102601 4922
rect 102601 4870 102647 4922
rect 102351 4868 102407 4870
rect 102431 4868 102487 4870
rect 102511 4868 102567 4870
rect 102591 4868 102647 4870
rect 102230 4120 102286 4176
rect 102351 3834 102407 3836
rect 102431 3834 102487 3836
rect 102511 3834 102567 3836
rect 102591 3834 102647 3836
rect 102351 3782 102397 3834
rect 102397 3782 102407 3834
rect 102431 3782 102461 3834
rect 102461 3782 102473 3834
rect 102473 3782 102487 3834
rect 102511 3782 102525 3834
rect 102525 3782 102537 3834
rect 102537 3782 102567 3834
rect 102591 3782 102601 3834
rect 102601 3782 102647 3834
rect 102351 3780 102407 3782
rect 102431 3780 102487 3782
rect 102511 3780 102567 3782
rect 102591 3780 102647 3782
rect 105634 10240 105690 10296
rect 106278 10240 106334 10296
rect 103426 8200 103482 8256
rect 103150 3460 103206 3496
rect 103150 3440 103152 3460
rect 103152 3440 103204 3460
rect 103204 3440 103206 3460
rect 102351 2746 102407 2748
rect 102431 2746 102487 2748
rect 102511 2746 102567 2748
rect 102591 2746 102647 2748
rect 102351 2694 102397 2746
rect 102397 2694 102407 2746
rect 102431 2694 102461 2746
rect 102461 2694 102473 2746
rect 102473 2694 102487 2746
rect 102511 2694 102525 2746
rect 102525 2694 102537 2746
rect 102537 2694 102567 2746
rect 102591 2694 102601 2746
rect 102601 2694 102647 2746
rect 102351 2692 102407 2694
rect 102431 2692 102487 2694
rect 102511 2692 102567 2694
rect 102591 2692 102647 2694
rect 101310 2388 101312 2408
rect 101312 2388 101364 2408
rect 101364 2388 101366 2408
rect 101310 2352 101366 2388
rect 100850 1672 100906 1728
rect 102351 1658 102407 1660
rect 102431 1658 102487 1660
rect 102511 1658 102567 1660
rect 102591 1658 102647 1660
rect 102351 1606 102397 1658
rect 102397 1606 102407 1658
rect 102431 1606 102461 1658
rect 102461 1606 102473 1658
rect 102473 1606 102487 1658
rect 102511 1606 102525 1658
rect 102525 1606 102537 1658
rect 102537 1606 102567 1658
rect 102591 1606 102601 1658
rect 102601 1606 102647 1658
rect 102351 1604 102407 1606
rect 102431 1604 102487 1606
rect 102511 1604 102567 1606
rect 102591 1604 102647 1606
rect 100758 856 100814 912
rect 103610 6568 103666 6624
rect 103426 3984 103482 4040
rect 103702 3596 103758 3632
rect 103702 3576 103704 3596
rect 103704 3576 103756 3596
rect 103756 3576 103758 3596
rect 107198 10240 107254 10296
rect 107750 10240 107806 10296
rect 108394 10240 108450 10296
rect 109038 10240 109094 10296
rect 110050 10240 110106 10296
rect 110786 10240 110842 10296
rect 111522 10240 111578 10296
rect 112350 10240 112406 10296
rect 112902 10240 112958 10296
rect 113546 10240 113602 10296
rect 114190 10240 114246 10296
rect 115202 10240 115258 10296
rect 115754 10240 115810 10296
rect 116674 10240 116730 10296
rect 117226 10240 117282 10296
rect 118054 10240 118110 10296
rect 118698 10240 118754 10296
rect 119342 10240 119398 10296
rect 120354 10240 120410 10296
rect 121090 10240 121146 10296
rect 121734 10240 121790 10296
rect 122378 10240 122434 10296
rect 104346 4936 104402 4992
rect 104530 3984 104586 4040
rect 104438 3712 104494 3768
rect 104622 3848 104678 3904
rect 104070 2080 104126 2136
rect 104254 2760 104310 2816
rect 104898 3848 104954 3904
rect 104990 3712 105046 3768
rect 106278 8200 106334 8256
rect 105450 4528 105506 4584
rect 104898 3168 104954 3224
rect 105634 3984 105690 4040
rect 106002 5888 106058 5944
rect 106002 4972 106004 4992
rect 106004 4972 106056 4992
rect 106056 4972 106058 4992
rect 106002 4936 106058 4972
rect 106186 4800 106242 4856
rect 106094 4528 106150 4584
rect 105818 3712 105874 3768
rect 105082 1844 105084 1864
rect 105084 1844 105136 1864
rect 105136 1844 105138 1864
rect 105082 1808 105138 1844
rect 104070 1264 104126 1320
rect 104162 856 104218 912
rect 105726 2760 105782 2816
rect 106278 4256 106334 4312
rect 107198 4256 107254 4312
rect 107106 3984 107162 4040
rect 106186 3476 106188 3496
rect 106188 3476 106240 3496
rect 106240 3476 106242 3496
rect 106186 3440 106242 3476
rect 106002 2488 106058 2544
rect 107566 3984 107622 4040
rect 107382 3440 107438 3496
rect 108210 6180 108266 6216
rect 108210 6160 108212 6180
rect 108212 6160 108264 6180
rect 108264 6160 108266 6180
rect 108026 3984 108082 4040
rect 108118 3440 108174 3496
rect 109038 5772 109094 5808
rect 109038 5752 109040 5772
rect 109040 5752 109092 5772
rect 109092 5752 109094 5772
rect 109130 5072 109186 5128
rect 108670 4936 108726 4992
rect 109222 3984 109278 4040
rect 108854 3712 108910 3768
rect 108946 3168 109002 3224
rect 104070 584 104126 640
rect 103518 312 103574 368
rect 109590 6316 109646 6352
rect 109590 6296 109592 6316
rect 109592 6296 109644 6316
rect 109644 6296 109646 6316
rect 109590 2796 109592 2816
rect 109592 2796 109644 2816
rect 109644 2796 109646 2816
rect 109590 2760 109646 2796
rect 109222 1420 109278 1456
rect 109222 1400 109224 1420
rect 109224 1400 109276 1420
rect 109276 1400 109278 1420
rect 110050 3984 110106 4040
rect 110786 5228 110842 5264
rect 110786 5208 110788 5228
rect 110788 5208 110840 5228
rect 110840 5208 110842 5228
rect 110694 3984 110750 4040
rect 110142 2488 110198 2544
rect 110326 2488 110382 2544
rect 108486 720 108542 776
rect 111246 3984 111302 4040
rect 111430 5480 111486 5536
rect 111430 5208 111486 5264
rect 111338 1420 111394 1456
rect 111338 1400 111340 1420
rect 111340 1400 111392 1420
rect 111392 1400 111394 1420
rect 111706 2760 111762 2816
rect 112166 6840 112222 6896
rect 112350 3984 112406 4040
rect 112350 1128 112406 1184
rect 112902 6160 112958 6216
rect 113086 5752 113142 5808
rect 113086 5072 113142 5128
rect 112994 3984 113050 4040
rect 113822 8064 113878 8120
rect 113454 6316 113510 6352
rect 113454 6296 113456 6316
rect 113456 6296 113508 6316
rect 113508 6296 113510 6316
rect 113362 3440 113418 3496
rect 113546 5344 113602 5400
rect 114006 7792 114062 7848
rect 114558 6568 114614 6624
rect 114466 5480 114522 5536
rect 114742 6296 114798 6352
rect 114834 6160 114890 6216
rect 114558 5344 114614 5400
rect 115478 7384 115534 7440
rect 115018 6432 115074 6488
rect 115662 7268 115718 7304
rect 115662 7248 115664 7268
rect 115664 7248 115716 7268
rect 115716 7248 115718 7268
rect 115018 5208 115074 5264
rect 114650 5072 114706 5128
rect 114558 4528 114614 4584
rect 114926 4664 114982 4720
rect 115018 3576 115074 3632
rect 114926 2896 114982 2952
rect 114558 2216 114614 2272
rect 114558 1400 114614 1456
rect 114834 1400 114890 1456
rect 115110 992 115166 1048
rect 114926 856 114982 912
rect 115570 1400 115626 1456
rect 116214 6740 116216 6760
rect 116216 6740 116268 6760
rect 116268 6740 116270 6760
rect 116214 6704 116270 6740
rect 115938 6024 115994 6080
rect 116030 5208 116086 5264
rect 116030 4664 116086 4720
rect 116582 6876 116584 6896
rect 116584 6876 116636 6896
rect 116636 6876 116638 6896
rect 116582 6840 116638 6876
rect 116490 6024 116546 6080
rect 116490 5888 116546 5944
rect 116398 5752 116454 5808
rect 116950 7928 117006 7984
rect 117594 5244 117596 5264
rect 117596 5244 117648 5264
rect 117648 5244 117650 5264
rect 117594 5208 117650 5244
rect 117226 3304 117282 3360
rect 117226 2760 117282 2816
rect 117870 6296 117926 6352
rect 117870 5888 117926 5944
rect 118146 6160 118202 6216
rect 117318 1400 117374 1456
rect 117686 1964 117742 2000
rect 117686 1944 117688 1964
rect 117688 1944 117740 1964
rect 117740 1944 117742 1964
rect 118882 6704 118938 6760
rect 120262 7792 120318 7848
rect 119250 7112 119306 7168
rect 119986 6840 120042 6896
rect 119434 2488 119490 2544
rect 120814 2624 120870 2680
rect 121090 2624 121146 2680
rect 121366 4664 121422 4720
rect 123206 10240 123262 10296
rect 124034 10240 124090 10296
rect 122102 7384 122158 7440
rect 121918 6024 121974 6080
rect 121918 5652 121920 5672
rect 121920 5652 121972 5672
rect 121972 5652 121974 5672
rect 121918 5616 121974 5652
rect 125598 10376 125654 10432
rect 125230 10240 125286 10296
rect 124126 2760 124182 2816
rect 124126 2624 124182 2680
rect 123482 2080 123538 2136
rect 124126 2080 124182 2136
rect 126334 10240 126390 10296
rect 126978 10240 127034 10296
rect 121826 1808 121882 1864
rect 122102 1844 122104 1864
rect 122104 1844 122156 1864
rect 122156 1844 122158 1864
rect 122102 1808 122158 1844
rect 127714 10240 127770 10296
rect 128266 10240 128322 10296
rect 129278 10240 129334 10296
rect 129646 10240 129702 10296
rect 130750 10240 130806 10296
rect 127714 6160 127770 6216
rect 126978 1400 127034 1456
rect 128450 1400 128506 1456
rect 124402 584 124458 640
rect 125322 584 125378 640
rect 126242 584 126298 640
rect 131486 10240 131542 10296
rect 132130 10240 132186 10296
rect 129186 584 129242 640
rect 117778 448 117834 504
rect 118054 448 118110 504
rect 118698 448 118754 504
rect 119342 448 119398 504
rect 120354 448 120410 504
rect 121090 448 121146 504
rect 121826 448 121882 504
rect 122654 448 122710 504
rect 123390 448 123446 504
rect 127806 448 127862 504
rect 132958 10240 133014 10296
rect 133418 10240 133474 10296
rect 134154 10240 134210 10296
rect 134706 10240 134762 10296
rect 138754 10240 138810 10296
rect 136149 9818 136205 9820
rect 136229 9818 136285 9820
rect 136309 9818 136365 9820
rect 136389 9818 136445 9820
rect 136149 9766 136195 9818
rect 136195 9766 136205 9818
rect 136229 9766 136259 9818
rect 136259 9766 136271 9818
rect 136271 9766 136285 9818
rect 136309 9766 136323 9818
rect 136323 9766 136335 9818
rect 136335 9766 136365 9818
rect 136389 9766 136399 9818
rect 136399 9766 136445 9818
rect 136149 9764 136205 9766
rect 136229 9764 136285 9766
rect 136309 9764 136365 9766
rect 136389 9764 136445 9766
rect 138018 9580 138074 9616
rect 139398 10104 139454 10160
rect 139766 9832 139822 9888
rect 138018 9560 138020 9580
rect 138020 9560 138072 9580
rect 138072 9560 138074 9580
rect 133786 2760 133842 2816
rect 136149 8730 136205 8732
rect 136229 8730 136285 8732
rect 136309 8730 136365 8732
rect 136389 8730 136445 8732
rect 136149 8678 136195 8730
rect 136195 8678 136205 8730
rect 136229 8678 136259 8730
rect 136259 8678 136271 8730
rect 136271 8678 136285 8730
rect 136309 8678 136323 8730
rect 136323 8678 136335 8730
rect 136335 8678 136365 8730
rect 136389 8678 136399 8730
rect 136399 8678 136445 8730
rect 136149 8676 136205 8678
rect 136229 8676 136285 8678
rect 136309 8676 136365 8678
rect 136389 8676 136445 8678
rect 136149 7642 136205 7644
rect 136229 7642 136285 7644
rect 136309 7642 136365 7644
rect 136389 7642 136445 7644
rect 136149 7590 136195 7642
rect 136195 7590 136205 7642
rect 136229 7590 136259 7642
rect 136259 7590 136271 7642
rect 136271 7590 136285 7642
rect 136309 7590 136323 7642
rect 136323 7590 136335 7642
rect 136335 7590 136365 7642
rect 136389 7590 136399 7642
rect 136399 7590 136445 7642
rect 136149 7588 136205 7590
rect 136229 7588 136285 7590
rect 136309 7588 136365 7590
rect 136389 7588 136445 7590
rect 136149 6554 136205 6556
rect 136229 6554 136285 6556
rect 136309 6554 136365 6556
rect 136389 6554 136445 6556
rect 136149 6502 136195 6554
rect 136195 6502 136205 6554
rect 136229 6502 136259 6554
rect 136259 6502 136271 6554
rect 136271 6502 136285 6554
rect 136309 6502 136323 6554
rect 136323 6502 136335 6554
rect 136335 6502 136365 6554
rect 136389 6502 136399 6554
rect 136399 6502 136445 6554
rect 136149 6500 136205 6502
rect 136229 6500 136285 6502
rect 136309 6500 136365 6502
rect 136389 6500 136445 6502
rect 137282 5752 137338 5808
rect 136086 5652 136088 5672
rect 136088 5652 136140 5672
rect 136140 5652 136142 5672
rect 136086 5616 136142 5652
rect 136149 5466 136205 5468
rect 136229 5466 136285 5468
rect 136309 5466 136365 5468
rect 136389 5466 136445 5468
rect 136149 5414 136195 5466
rect 136195 5414 136205 5466
rect 136229 5414 136259 5466
rect 136259 5414 136271 5466
rect 136271 5414 136285 5466
rect 136309 5414 136323 5466
rect 136323 5414 136335 5466
rect 136335 5414 136365 5466
rect 136389 5414 136399 5466
rect 136399 5414 136445 5466
rect 136149 5412 136205 5414
rect 136229 5412 136285 5414
rect 136309 5412 136365 5414
rect 136389 5412 136445 5414
rect 138846 7520 138902 7576
rect 136149 4378 136205 4380
rect 136229 4378 136285 4380
rect 136309 4378 136365 4380
rect 136389 4378 136445 4380
rect 136149 4326 136195 4378
rect 136195 4326 136205 4378
rect 136229 4326 136259 4378
rect 136259 4326 136271 4378
rect 136271 4326 136285 4378
rect 136309 4326 136323 4378
rect 136323 4326 136335 4378
rect 136335 4326 136365 4378
rect 136389 4326 136399 4378
rect 136399 4326 136445 4378
rect 136149 4324 136205 4326
rect 136229 4324 136285 4326
rect 136309 4324 136365 4326
rect 136389 4324 136445 4326
rect 136149 3290 136205 3292
rect 136229 3290 136285 3292
rect 136309 3290 136365 3292
rect 136389 3290 136445 3292
rect 136149 3238 136195 3290
rect 136195 3238 136205 3290
rect 136229 3238 136259 3290
rect 136259 3238 136271 3290
rect 136271 3238 136285 3290
rect 136309 3238 136323 3290
rect 136323 3238 136335 3290
rect 136335 3238 136365 3290
rect 136389 3238 136399 3290
rect 136399 3238 136445 3290
rect 136149 3236 136205 3238
rect 136229 3236 136285 3238
rect 136309 3236 136365 3238
rect 136389 3236 136445 3238
rect 134154 2488 134210 2544
rect 130842 584 130898 640
rect 131670 584 131726 640
rect 136149 2202 136205 2204
rect 136229 2202 136285 2204
rect 136309 2202 136365 2204
rect 136389 2202 136445 2204
rect 136149 2150 136195 2202
rect 136195 2150 136205 2202
rect 136229 2150 136259 2202
rect 136259 2150 136271 2202
rect 136271 2150 136285 2202
rect 136309 2150 136323 2202
rect 136323 2150 136335 2202
rect 136335 2150 136365 2202
rect 136389 2150 136399 2202
rect 136399 2150 136445 2202
rect 136149 2148 136205 2150
rect 136229 2148 136285 2150
rect 136309 2148 136365 2150
rect 136389 2148 136445 2150
rect 135258 1400 135314 1456
rect 138018 1436 138020 1456
rect 138020 1436 138072 1456
rect 138072 1436 138074 1456
rect 138018 1400 138074 1436
rect 139214 4392 139270 4448
rect 136149 1114 136205 1116
rect 136229 1114 136285 1116
rect 136309 1114 136365 1116
rect 136389 1114 136445 1116
rect 136149 1062 136195 1114
rect 136195 1062 136205 1114
rect 136229 1062 136259 1114
rect 136259 1062 136271 1114
rect 136271 1062 136285 1114
rect 136309 1062 136323 1114
rect 136323 1062 136335 1114
rect 136335 1062 136365 1114
rect 136389 1062 136399 1114
rect 136399 1062 136445 1114
rect 136149 1060 136205 1062
rect 136229 1060 136285 1062
rect 136309 1060 136365 1062
rect 136389 1060 136445 1062
rect 139766 6296 139822 6352
rect 139766 5888 139822 5944
rect 139858 4392 139914 4448
rect 139950 3440 140006 3496
rect 140042 2760 140098 2816
rect 143262 10240 143318 10296
rect 140686 10104 140742 10160
rect 141330 10104 141386 10160
rect 140226 1808 140282 1864
rect 139766 992 139822 1048
rect 138846 720 138902 776
rect 134522 584 134578 640
rect 138754 584 138810 640
rect 130750 312 130806 368
rect 132130 312 132186 368
rect 133234 312 133290 368
rect 141974 10104 142030 10160
rect 140686 5616 140742 5672
rect 140962 4020 140964 4040
rect 140964 4020 141016 4040
rect 141016 4020 141018 4040
rect 140962 3984 141018 4020
rect 140870 2760 140926 2816
rect 143538 10104 143594 10160
rect 144550 10104 144606 10160
rect 144918 9832 144974 9888
rect 142434 6704 142490 6760
rect 141514 4936 141570 4992
rect 141606 4392 141662 4448
rect 141514 4120 141570 4176
rect 141790 3984 141846 4040
rect 142066 3032 142122 3088
rect 141606 1844 141608 1864
rect 141608 1844 141660 1864
rect 141660 1844 141662 1864
rect 141606 1808 141662 1844
rect 140686 1400 140742 1456
rect 143538 3848 143594 3904
rect 104162 176 104218 232
rect 140318 176 140374 232
rect 143906 2896 143962 2952
rect 145102 8472 145158 8528
rect 144918 6432 144974 6488
rect 144826 5652 144828 5672
rect 144828 5652 144880 5672
rect 144880 5652 144882 5672
rect 144826 5616 144882 5652
rect 144826 3304 144882 3360
rect 144734 3168 144790 3224
rect 143630 856 143686 912
rect 141790 720 141846 776
rect 144550 1264 144606 1320
rect 144734 856 144790 912
rect 143998 448 144054 504
rect 141422 312 141478 368
rect 144918 720 144974 776
rect 144918 620 144920 640
rect 144920 620 144972 640
rect 144972 620 144974 640
rect 144918 584 144974 620
rect 145838 10104 145894 10160
rect 146298 10104 146354 10160
rect 145562 4120 145618 4176
rect 145470 2796 145472 2816
rect 145472 2796 145524 2816
rect 145524 2796 145526 2816
rect 145470 2760 145526 2796
rect 146298 6296 146354 6352
rect 146390 3576 146446 3632
rect 146482 3440 146538 3496
rect 146298 2352 146354 2408
rect 148414 10512 148470 10568
rect 147126 10104 147182 10160
rect 146666 3712 146722 3768
rect 147218 3460 147274 3496
rect 147218 3440 147220 3460
rect 147220 3440 147272 3460
rect 147272 3440 147274 3460
rect 147586 2080 147642 2136
rect 146850 1672 146906 1728
rect 148506 6024 148562 6080
rect 149058 10240 149114 10296
rect 149702 10104 149758 10160
rect 150990 10104 151046 10160
rect 151634 10104 151690 10160
rect 150070 9832 150126 9888
rect 148322 992 148378 1048
rect 147678 720 147734 776
rect 148414 720 148470 776
rect 146942 312 146998 368
rect 147862 584 147918 640
rect 149334 1672 149390 1728
rect 92202 40 92258 96
rect 98274 40 98330 96
rect 141238 40 141294 96
rect 149978 7928 150034 7984
rect 150070 5480 150126 5536
rect 149978 5208 150034 5264
rect 150254 5208 150310 5264
rect 149978 4800 150034 4856
rect 150162 4800 150218 4856
rect 149886 4684 149942 4720
rect 149886 4664 149888 4684
rect 149888 4664 149940 4684
rect 149940 4664 149942 4684
rect 150070 4256 150126 4312
rect 149610 3168 149666 3224
rect 149610 1944 149666 2000
rect 149978 1944 150034 2000
rect 149610 1672 149666 1728
rect 154302 10376 154358 10432
rect 152278 10104 152334 10160
rect 152830 10104 152886 10160
rect 154210 10104 154266 10160
rect 150346 3576 150402 3632
rect 150346 2896 150402 2952
rect 150254 1536 150310 1592
rect 149518 1128 149574 1184
rect 150622 1400 150678 1456
rect 150438 720 150494 776
rect 155222 9832 155278 9888
rect 151726 5344 151782 5400
rect 151726 5072 151782 5128
rect 151266 2080 151322 2136
rect 151358 992 151414 1048
rect 152002 6432 152058 6488
rect 151910 5108 151912 5128
rect 151912 5108 151964 5128
rect 151964 5108 151966 5128
rect 151910 5072 151966 5108
rect 152462 6724 152518 6760
rect 152462 6704 152464 6724
rect 152464 6704 152516 6724
rect 152516 6704 152518 6724
rect 152094 5652 152096 5672
rect 152096 5652 152148 5672
rect 152148 5652 152150 5672
rect 152094 5616 152150 5652
rect 152002 4020 152004 4040
rect 152004 4020 152056 4040
rect 152056 4020 152058 4040
rect 152002 3984 152058 4020
rect 153106 5072 153162 5128
rect 152922 4936 152978 4992
rect 152370 3848 152426 3904
rect 152002 3168 152058 3224
rect 151726 2352 151782 2408
rect 153566 5480 153622 5536
rect 152922 3304 152978 3360
rect 156694 9444 156750 9480
rect 156694 9424 156696 9444
rect 156696 9424 156748 9444
rect 156748 9424 156750 9444
rect 153934 6976 153990 7032
rect 153842 6724 153898 6760
rect 153842 6704 153844 6724
rect 153844 6704 153896 6724
rect 153896 6704 153898 6724
rect 153658 2932 153660 2952
rect 153660 2932 153712 2952
rect 153712 2932 153714 2952
rect 153658 2896 153714 2932
rect 154578 7656 154634 7712
rect 154762 8064 154818 8120
rect 154762 5208 154818 5264
rect 154578 4528 154634 4584
rect 154026 4120 154082 4176
rect 153106 1536 153162 1592
rect 152094 1400 152150 1456
rect 152462 1264 152518 1320
rect 152370 992 152426 1048
rect 154118 3168 154174 3224
rect 154302 3304 154358 3360
rect 154394 2760 154450 2816
rect 154394 2216 154450 2272
rect 154118 584 154174 640
rect 154486 1264 154542 1320
rect 155038 2896 155094 2952
rect 156050 9036 156106 9072
rect 156050 9016 156052 9036
rect 156052 9016 156104 9036
rect 156104 9016 156106 9036
rect 156050 8628 156106 8664
rect 156050 8608 156052 8628
rect 156052 8608 156104 8628
rect 156104 8608 156106 8628
rect 156050 7792 156106 7848
rect 156142 3712 156198 3768
rect 155866 2896 155922 2952
rect 156418 2760 156474 2816
rect 156234 2488 156290 2544
rect 156602 2488 156658 2544
rect 157430 9036 157486 9072
rect 157430 9016 157432 9036
rect 157432 9016 157484 9036
rect 157484 9016 157486 9036
rect 157706 8472 157762 8528
rect 157062 2896 157118 2952
rect 156970 2624 157026 2680
rect 155958 1400 156014 1456
rect 157246 8336 157302 8392
rect 158718 8084 158774 8120
rect 158718 8064 158720 8084
rect 158720 8064 158772 8084
rect 158772 8064 158774 8084
rect 157798 7384 157854 7440
rect 157246 3712 157302 3768
rect 156602 1672 156658 1728
rect 156786 1672 156842 1728
rect 157246 1400 157302 1456
rect 155774 1128 155830 1184
rect 158166 6432 158222 6488
rect 158534 4800 158590 4856
rect 159362 8336 159418 8392
rect 159454 8084 159510 8120
rect 159454 8064 159456 8084
rect 159456 8064 159508 8084
rect 159508 8064 159510 8084
rect 158626 1264 158682 1320
rect 160926 8336 160982 8392
rect 161018 8084 161074 8120
rect 161018 8064 161020 8084
rect 161020 8064 161072 8084
rect 161072 8064 161074 8084
rect 160006 3576 160062 3632
rect 159362 1128 159418 1184
rect 158442 992 158498 1048
rect 160374 1264 160430 1320
rect 161202 8064 161258 8120
rect 161386 6976 161442 7032
rect 162398 8336 162454 8392
rect 162398 7792 162454 7848
rect 161294 3848 161350 3904
rect 160834 1128 160890 1184
rect 163318 8064 163374 8120
rect 163318 7792 163374 7848
rect 163778 9016 163834 9072
rect 163870 8336 163926 8392
rect 163962 8084 164018 8120
rect 163962 8064 163964 8084
rect 163964 8064 164016 8084
rect 164016 8064 164018 8084
rect 162950 1672 163006 1728
rect 160374 720 160430 776
rect 160558 720 160614 776
rect 160098 584 160154 640
rect 161662 1128 161718 1184
rect 165250 8336 165306 8392
rect 165342 8084 165398 8120
rect 165342 8064 165344 8084
rect 165344 8064 165396 8084
rect 165396 8064 165398 8084
rect 172242 10512 172298 10568
rect 171690 10240 171746 10296
rect 168378 9716 168434 9752
rect 168378 9696 168380 9716
rect 168380 9696 168432 9716
rect 168432 9696 168434 9716
rect 169482 9696 169538 9752
rect 166538 8336 166594 8392
rect 166906 8336 166962 8392
rect 163870 1128 163926 1184
rect 169948 9274 170004 9276
rect 170028 9274 170084 9276
rect 170108 9274 170164 9276
rect 170188 9274 170244 9276
rect 169948 9222 169994 9274
rect 169994 9222 170004 9274
rect 170028 9222 170058 9274
rect 170058 9222 170070 9274
rect 170070 9222 170084 9274
rect 170108 9222 170122 9274
rect 170122 9222 170134 9274
rect 170134 9222 170164 9274
rect 170188 9222 170198 9274
rect 170198 9222 170244 9274
rect 169948 9220 170004 9222
rect 170028 9220 170084 9222
rect 170108 9220 170164 9222
rect 170188 9220 170244 9222
rect 169758 9152 169814 9208
rect 171046 8200 171102 8256
rect 169948 8186 170004 8188
rect 170028 8186 170084 8188
rect 170108 8186 170164 8188
rect 170188 8186 170244 8188
rect 169948 8134 169994 8186
rect 169994 8134 170004 8186
rect 170028 8134 170058 8186
rect 170058 8134 170070 8186
rect 170070 8134 170084 8186
rect 170108 8134 170122 8186
rect 170122 8134 170134 8186
rect 170134 8134 170164 8186
rect 170188 8134 170198 8186
rect 170198 8134 170244 8186
rect 169948 8132 170004 8134
rect 170028 8132 170084 8134
rect 170108 8132 170164 8134
rect 170188 8132 170244 8134
rect 168286 6704 168342 6760
rect 168286 5752 168342 5808
rect 168838 6160 168894 6216
rect 169574 7112 169630 7168
rect 169206 5752 169262 5808
rect 169948 7098 170004 7100
rect 170028 7098 170084 7100
rect 170108 7098 170164 7100
rect 170188 7098 170244 7100
rect 169948 7046 169994 7098
rect 169994 7046 170004 7098
rect 170028 7046 170058 7098
rect 170058 7046 170070 7098
rect 170070 7046 170084 7098
rect 170108 7046 170122 7098
rect 170122 7046 170134 7098
rect 170134 7046 170164 7098
rect 170188 7046 170198 7098
rect 170198 7046 170244 7098
rect 169948 7044 170004 7046
rect 170028 7044 170084 7046
rect 170108 7044 170164 7046
rect 170188 7044 170244 7046
rect 170770 7792 170826 7848
rect 170586 6568 170642 6624
rect 169758 6316 169814 6352
rect 169758 6296 169760 6316
rect 169760 6296 169812 6316
rect 169812 6296 169814 6316
rect 171138 7384 171194 7440
rect 173990 10376 174046 10432
rect 173898 10240 173954 10296
rect 174450 10240 174506 10296
rect 175186 10240 175242 10296
rect 175922 10240 175978 10296
rect 176750 10240 176806 10296
rect 177486 10240 177542 10296
rect 172518 7656 172574 7712
rect 172610 7112 172666 7168
rect 170770 6024 170826 6080
rect 169948 6010 170004 6012
rect 170028 6010 170084 6012
rect 170108 6010 170164 6012
rect 170188 6010 170244 6012
rect 169948 5958 169994 6010
rect 169994 5958 170004 6010
rect 170028 5958 170058 6010
rect 170058 5958 170070 6010
rect 170070 5958 170084 6010
rect 170108 5958 170122 6010
rect 170122 5958 170134 6010
rect 170134 5958 170164 6010
rect 170188 5958 170198 6010
rect 170198 5958 170244 6010
rect 169948 5956 170004 5958
rect 170028 5956 170084 5958
rect 170108 5956 170164 5958
rect 170188 5956 170244 5958
rect 172518 5616 172574 5672
rect 169948 4922 170004 4924
rect 170028 4922 170084 4924
rect 170108 4922 170164 4924
rect 170188 4922 170244 4924
rect 169948 4870 169994 4922
rect 169994 4870 170004 4922
rect 170028 4870 170058 4922
rect 170058 4870 170070 4922
rect 170070 4870 170084 4922
rect 170108 4870 170122 4922
rect 170122 4870 170134 4922
rect 170134 4870 170164 4922
rect 170188 4870 170198 4922
rect 170198 4870 170244 4922
rect 169948 4868 170004 4870
rect 170028 4868 170084 4870
rect 170108 4868 170164 4870
rect 170188 4868 170244 4870
rect 169666 4392 169722 4448
rect 169574 4120 169630 4176
rect 168378 1400 168434 1456
rect 169948 3834 170004 3836
rect 170028 3834 170084 3836
rect 170108 3834 170164 3836
rect 170188 3834 170244 3836
rect 169948 3782 169994 3834
rect 169994 3782 170004 3834
rect 170028 3782 170058 3834
rect 170058 3782 170070 3834
rect 170070 3782 170084 3834
rect 170108 3782 170122 3834
rect 170122 3782 170134 3834
rect 170134 3782 170164 3834
rect 170188 3782 170198 3834
rect 170198 3782 170244 3834
rect 169948 3780 170004 3782
rect 170028 3780 170084 3782
rect 170108 3780 170164 3782
rect 170188 3780 170244 3782
rect 180522 10512 180578 10568
rect 177946 10240 178002 10296
rect 179142 10240 179198 10296
rect 180430 10240 180486 10296
rect 175278 5344 175334 5400
rect 181810 10376 181866 10432
rect 181902 10240 181958 10296
rect 191286 10376 191342 10432
rect 192850 10376 192906 10432
rect 182546 10240 182602 10296
rect 183282 10240 183338 10296
rect 184294 10240 184350 10296
rect 184754 10240 184810 10296
rect 185490 10240 185546 10296
rect 186226 10240 186282 10296
rect 186962 10240 187018 10296
rect 187698 10240 187754 10296
rect 188618 10240 188674 10296
rect 189446 10240 189502 10296
rect 189906 10240 189962 10296
rect 179418 8200 179474 8256
rect 185858 6432 185914 6488
rect 178406 4664 178462 4720
rect 173806 4256 173862 4312
rect 169948 2746 170004 2748
rect 170028 2746 170084 2748
rect 170108 2746 170164 2748
rect 170188 2746 170244 2748
rect 169948 2694 169994 2746
rect 169994 2694 170004 2746
rect 170028 2694 170058 2746
rect 170058 2694 170070 2746
rect 170070 2694 170084 2746
rect 170108 2694 170122 2746
rect 170122 2694 170134 2746
rect 170134 2694 170164 2746
rect 170188 2694 170198 2746
rect 170198 2694 170244 2746
rect 169948 2692 170004 2694
rect 170028 2692 170084 2694
rect 170108 2692 170164 2694
rect 170188 2692 170244 2694
rect 169948 1658 170004 1660
rect 170028 1658 170084 1660
rect 170108 1658 170164 1660
rect 170188 1658 170244 1660
rect 169948 1606 169994 1658
rect 169994 1606 170004 1658
rect 170028 1606 170058 1658
rect 170058 1606 170070 1658
rect 170070 1606 170084 1658
rect 170108 1606 170122 1658
rect 170122 1606 170134 1658
rect 170134 1606 170164 1658
rect 170188 1606 170198 1658
rect 170198 1606 170244 1658
rect 169948 1604 170004 1606
rect 170028 1604 170084 1606
rect 170108 1604 170164 1606
rect 170188 1604 170244 1606
rect 166998 1264 167054 1320
rect 165250 1128 165306 1184
rect 165986 1128 166042 1184
rect 166814 1128 166870 1184
rect 162122 584 162178 640
rect 163502 584 163558 640
rect 164606 584 164662 640
rect 168378 992 168434 1048
rect 170310 992 170366 1048
rect 169022 584 169078 640
rect 171690 584 171746 640
rect 172242 584 172298 640
rect 176658 3032 176714 3088
rect 174726 1844 174728 1864
rect 174728 1844 174780 1864
rect 174780 1844 174782 1864
rect 172978 584 173034 640
rect 173898 584 173954 640
rect 161294 312 161350 368
rect 167918 312 167974 368
rect 174726 1808 174782 1844
rect 174450 584 174506 640
rect 175278 584 175334 640
rect 176842 2216 176898 2272
rect 179418 2080 179474 2136
rect 176658 584 176714 640
rect 176566 448 176622 504
rect 180522 992 180578 1048
rect 177854 584 177910 640
rect 178498 584 178554 640
rect 179142 584 179198 640
rect 179602 584 179658 640
rect 180338 584 180394 640
rect 180522 584 180578 640
rect 189446 6704 189502 6760
rect 189998 6160 190054 6216
rect 186410 3168 186466 3224
rect 181810 448 181866 504
rect 176842 312 176898 368
rect 181718 312 181774 368
rect 160558 176 160614 232
rect 174266 176 174322 232
rect 160006 40 160062 96
rect 183006 448 183062 504
rect 183282 448 183338 504
rect 184294 448 184350 504
rect 186318 1400 186374 1456
rect 184754 448 184810 504
rect 185490 448 185546 504
rect 186962 448 187018 504
rect 190366 2760 190422 2816
rect 191378 10240 191434 10296
rect 191746 2760 191802 2816
rect 192942 10240 192998 10296
rect 194046 10240 194102 10296
rect 194322 10240 194378 10296
rect 195518 10240 195574 10296
rect 195794 10240 195850 10296
rect 195334 8200 195390 8256
rect 196530 10240 196586 10296
rect 197266 10240 197322 10296
rect 198002 10240 198058 10296
rect 199106 10240 199162 10296
rect 199934 10240 199990 10296
rect 191838 1944 191894 2000
rect 192114 1944 192170 2000
rect 194598 1808 194654 1864
rect 196070 1808 196126 1864
rect 188158 448 188214 504
rect 188618 448 188674 504
rect 189446 448 189502 504
rect 191102 448 191158 504
rect 197358 1400 197414 1456
rect 200762 10240 200818 10296
rect 200946 10240 201002 10296
rect 198646 2760 198702 2816
rect 200026 2760 200082 2816
rect 208306 10512 208362 10568
rect 213458 10512 213514 10568
rect 202418 10376 202474 10432
rect 202510 10240 202566 10296
rect 204074 10240 204130 10296
rect 205822 10240 205878 10296
rect 201406 2760 201462 2816
rect 203746 9818 203802 9820
rect 203826 9818 203882 9820
rect 203906 9818 203962 9820
rect 203986 9818 204042 9820
rect 203746 9766 203792 9818
rect 203792 9766 203802 9818
rect 203826 9766 203856 9818
rect 203856 9766 203868 9818
rect 203868 9766 203882 9818
rect 203906 9766 203920 9818
rect 203920 9766 203932 9818
rect 203932 9766 203962 9818
rect 203986 9766 203996 9818
rect 203996 9766 204042 9818
rect 203746 9764 203802 9766
rect 203826 9764 203882 9766
rect 203906 9764 203962 9766
rect 203986 9764 204042 9766
rect 206558 10104 206614 10160
rect 207662 10104 207718 10160
rect 210882 10376 210938 10432
rect 208950 10104 209006 10160
rect 209318 10104 209374 10160
rect 211158 10104 211214 10160
rect 203746 8730 203802 8732
rect 203826 8730 203882 8732
rect 203906 8730 203962 8732
rect 203986 8730 204042 8732
rect 203746 8678 203792 8730
rect 203792 8678 203802 8730
rect 203826 8678 203856 8730
rect 203856 8678 203868 8730
rect 203868 8678 203882 8730
rect 203906 8678 203920 8730
rect 203920 8678 203932 8730
rect 203932 8678 203962 8730
rect 203986 8678 203996 8730
rect 203996 8678 204042 8730
rect 203746 8676 203802 8678
rect 203826 8676 203882 8678
rect 203906 8676 203962 8678
rect 203986 8676 204042 8678
rect 203746 7642 203802 7644
rect 203826 7642 203882 7644
rect 203906 7642 203962 7644
rect 203986 7642 204042 7644
rect 203746 7590 203792 7642
rect 203792 7590 203802 7642
rect 203826 7590 203856 7642
rect 203856 7590 203868 7642
rect 203868 7590 203882 7642
rect 203906 7590 203920 7642
rect 203920 7590 203932 7642
rect 203932 7590 203962 7642
rect 203986 7590 203996 7642
rect 203996 7590 204042 7642
rect 203746 7588 203802 7590
rect 203826 7588 203882 7590
rect 203906 7588 203962 7590
rect 203986 7588 204042 7590
rect 203746 6554 203802 6556
rect 203826 6554 203882 6556
rect 203906 6554 203962 6556
rect 203986 6554 204042 6556
rect 203746 6502 203792 6554
rect 203792 6502 203802 6554
rect 203826 6502 203856 6554
rect 203856 6502 203868 6554
rect 203868 6502 203882 6554
rect 203906 6502 203920 6554
rect 203920 6502 203932 6554
rect 203932 6502 203962 6554
rect 203986 6502 203996 6554
rect 203996 6502 204042 6554
rect 203746 6500 203802 6502
rect 203826 6500 203882 6502
rect 203906 6500 203962 6502
rect 203986 6500 204042 6502
rect 206190 5480 206246 5536
rect 203746 5466 203802 5468
rect 203826 5466 203882 5468
rect 203906 5466 203962 5468
rect 203986 5466 204042 5468
rect 203746 5414 203792 5466
rect 203792 5414 203802 5466
rect 203826 5414 203856 5466
rect 203856 5414 203868 5466
rect 203868 5414 203882 5466
rect 203906 5414 203920 5466
rect 203920 5414 203932 5466
rect 203932 5414 203962 5466
rect 203986 5414 203996 5466
rect 203996 5414 204042 5466
rect 203746 5412 203802 5414
rect 203826 5412 203882 5414
rect 203906 5412 203962 5414
rect 203986 5412 204042 5414
rect 203746 4378 203802 4380
rect 203826 4378 203882 4380
rect 203906 4378 203962 4380
rect 203986 4378 204042 4380
rect 203746 4326 203792 4378
rect 203792 4326 203802 4378
rect 203826 4326 203856 4378
rect 203856 4326 203868 4378
rect 203868 4326 203882 4378
rect 203906 4326 203920 4378
rect 203920 4326 203932 4378
rect 203932 4326 203962 4378
rect 203986 4326 203996 4378
rect 203996 4326 204042 4378
rect 203746 4324 203802 4326
rect 203826 4324 203882 4326
rect 203906 4324 203962 4326
rect 203986 4324 204042 4326
rect 203746 3290 203802 3292
rect 203826 3290 203882 3292
rect 203906 3290 203962 3292
rect 203986 3290 204042 3292
rect 203746 3238 203792 3290
rect 203792 3238 203802 3290
rect 203826 3238 203856 3290
rect 203856 3238 203868 3290
rect 203868 3238 203882 3290
rect 203906 3238 203920 3290
rect 203920 3238 203932 3290
rect 203932 3238 203962 3290
rect 203986 3238 203996 3290
rect 203996 3238 204042 3290
rect 203746 3236 203802 3238
rect 203826 3236 203882 3238
rect 203906 3236 203962 3238
rect 203986 3236 204042 3238
rect 207110 7656 207166 7712
rect 203746 2202 203802 2204
rect 203826 2202 203882 2204
rect 203906 2202 203962 2204
rect 203986 2202 204042 2204
rect 203746 2150 203792 2202
rect 203792 2150 203802 2202
rect 203826 2150 203856 2202
rect 203856 2150 203868 2202
rect 203868 2150 203882 2202
rect 203906 2150 203920 2202
rect 203920 2150 203932 2202
rect 203932 2150 203962 2202
rect 203986 2150 203996 2202
rect 203996 2150 204042 2202
rect 203746 2148 203802 2150
rect 203826 2148 203882 2150
rect 203906 2148 203962 2150
rect 203986 2148 204042 2150
rect 202878 1400 202934 1456
rect 203746 1114 203802 1116
rect 203826 1114 203882 1116
rect 203906 1114 203962 1116
rect 203986 1114 204042 1116
rect 203746 1062 203792 1114
rect 203792 1062 203802 1114
rect 203826 1062 203856 1114
rect 203856 1062 203868 1114
rect 203868 1062 203882 1114
rect 203906 1062 203920 1114
rect 203920 1062 203932 1114
rect 203932 1062 203962 1114
rect 203986 1062 203996 1114
rect 203996 1062 204042 1114
rect 203746 1060 203802 1062
rect 203826 1060 203882 1062
rect 203906 1060 203962 1062
rect 203986 1060 204042 1062
rect 208398 5108 208400 5128
rect 208400 5108 208452 5128
rect 208452 5108 208454 5128
rect 208398 5072 208454 5108
rect 205822 856 205878 912
rect 206558 856 206614 912
rect 207662 856 207718 912
rect 209318 6568 209374 6624
rect 209134 6432 209190 6488
rect 209134 5480 209190 5536
rect 209318 3848 209374 3904
rect 192850 448 192906 504
rect 193586 448 193642 504
rect 195610 448 195666 504
rect 196622 448 196678 504
rect 199934 448 199990 504
rect 201222 448 201278 504
rect 202418 448 202474 504
rect 204074 448 204130 504
rect 208582 1536 208638 1592
rect 208490 448 208546 504
rect 209686 2760 209742 2816
rect 209686 1400 209742 1456
rect 208950 856 209006 912
rect 192574 312 192630 368
rect 208306 312 208362 368
rect 209778 992 209834 1048
rect 209962 3168 210018 3224
rect 212538 10104 212594 10160
rect 211710 9832 211766 9888
rect 216586 10396 216642 10432
rect 216586 10376 216588 10396
rect 216588 10376 216640 10396
rect 216640 10376 216642 10396
rect 213918 10104 213974 10160
rect 214470 10104 214526 10160
rect 216678 10104 216734 10160
rect 215206 9716 215262 9752
rect 215206 9696 215208 9716
rect 215208 9696 215260 9716
rect 215260 9696 215262 9716
rect 215482 9580 215538 9616
rect 215482 9560 215484 9580
rect 215484 9560 215536 9580
rect 215536 9560 215538 9580
rect 212170 4700 212172 4720
rect 212172 4700 212224 4720
rect 212224 4700 212226 4720
rect 212170 4664 212226 4700
rect 211526 3032 211582 3088
rect 210974 176 211030 232
rect 211802 1128 211858 1184
rect 213182 7248 213238 7304
rect 213090 6316 213146 6352
rect 213090 6296 213092 6316
rect 213092 6296 213144 6316
rect 213144 6296 213146 6316
rect 212814 5752 212870 5808
rect 213182 5480 213238 5536
rect 214010 9152 214066 9208
rect 213458 7404 213514 7440
rect 213458 7384 213460 7404
rect 213460 7384 213512 7404
rect 213512 7384 213514 7404
rect 214010 8200 214066 8256
rect 214194 8064 214250 8120
rect 213918 7792 213974 7848
rect 213734 6976 213790 7032
rect 213642 2216 213698 2272
rect 211894 992 211950 1048
rect 212998 332 213054 368
rect 212998 312 213000 332
rect 213000 312 213052 332
rect 213052 312 213054 332
rect 214470 5480 214526 5536
rect 214378 5344 214434 5400
rect 214378 4800 214434 4856
rect 214562 2488 214618 2544
rect 214378 2388 214380 2408
rect 214380 2388 214432 2408
rect 214432 2388 214434 2408
rect 214378 2352 214434 2388
rect 214746 4684 214802 4720
rect 214746 4664 214748 4684
rect 214748 4664 214800 4684
rect 214800 4664 214802 4684
rect 214010 1808 214066 1864
rect 214562 1672 214618 1728
rect 215206 3984 215262 4040
rect 216862 9832 216918 9888
rect 216770 9016 216826 9072
rect 216586 8200 216642 8256
rect 216402 6160 216458 6216
rect 217322 8336 217378 8392
rect 216586 6024 216642 6080
rect 216586 5752 216642 5808
rect 216402 5616 216458 5672
rect 215850 4936 215906 4992
rect 215942 2352 215998 2408
rect 216034 2080 216090 2136
rect 217046 3440 217102 3496
rect 217138 2896 217194 2952
rect 216862 2488 216918 2544
rect 218610 10512 218666 10568
rect 217966 10104 218022 10160
rect 218058 6840 218114 6896
rect 218334 6704 218390 6760
rect 217690 3168 217746 3224
rect 216126 1844 216128 1864
rect 216128 1844 216180 1864
rect 216180 1844 216182 1864
rect 216126 1808 216182 1844
rect 216402 1808 216458 1864
rect 215574 584 215630 640
rect 218242 3984 218298 4040
rect 219254 10104 219310 10160
rect 223486 10532 223542 10568
rect 223486 10512 223488 10532
rect 223488 10512 223540 10532
rect 223540 10512 223542 10532
rect 221830 10376 221886 10432
rect 220358 10240 220414 10296
rect 219070 7656 219126 7712
rect 219070 6976 219126 7032
rect 218978 6568 219034 6624
rect 218978 4664 219034 4720
rect 219070 4256 219126 4312
rect 219254 5888 219310 5944
rect 219254 4120 219310 4176
rect 220542 10104 220598 10160
rect 219438 7792 219494 7848
rect 220082 7520 220138 7576
rect 220082 7112 220138 7168
rect 219438 6024 219494 6080
rect 219438 5208 219494 5264
rect 219438 4392 219494 4448
rect 218886 3712 218942 3768
rect 219162 3304 219218 3360
rect 218334 1420 218390 1456
rect 218334 1400 218336 1420
rect 218336 1400 218388 1420
rect 218388 1400 218390 1420
rect 218058 1300 218060 1320
rect 218060 1300 218112 1320
rect 218112 1300 218114 1320
rect 218058 1264 218114 1300
rect 218058 720 218114 776
rect 216678 448 216734 504
rect 214470 348 214472 368
rect 214472 348 214524 368
rect 214524 348 214526 368
rect 214470 312 214526 348
rect 215574 312 215630 368
rect 218886 1808 218942 1864
rect 219898 6196 219900 6216
rect 219900 6196 219952 6216
rect 219952 6196 219954 6216
rect 219898 6160 219954 6196
rect 219990 5616 220046 5672
rect 223118 10104 223174 10160
rect 222014 9832 222070 9888
rect 220542 8744 220598 8800
rect 220450 6704 220506 6760
rect 220818 8472 220874 8528
rect 220542 4800 220598 4856
rect 219898 2624 219954 2680
rect 219346 1844 219348 1864
rect 219348 1844 219400 1864
rect 219400 1844 219402 1864
rect 219346 1808 219402 1844
rect 219898 1944 219954 2000
rect 220082 1944 220138 2000
rect 220818 4528 220874 4584
rect 220818 3712 220874 3768
rect 221002 2896 221058 2952
rect 221830 6840 221886 6896
rect 221462 3168 221518 3224
rect 220082 1672 220138 1728
rect 219714 1400 219770 1456
rect 221094 2488 221150 2544
rect 219162 584 219218 640
rect 220818 1284 220874 1320
rect 220818 1264 220820 1284
rect 220820 1264 220872 1284
rect 220872 1264 220874 1284
rect 221738 3984 221794 4040
rect 222014 7112 222070 7168
rect 222198 6452 222254 6488
rect 222198 6432 222200 6452
rect 222200 6432 222252 6452
rect 222252 6432 222254 6452
rect 222198 3984 222254 4040
rect 222106 3712 222162 3768
rect 222014 3576 222070 3632
rect 221738 1672 221794 1728
rect 222198 1264 222254 1320
rect 222566 3168 222622 3224
rect 222566 2760 222622 2816
rect 223302 8336 223358 8392
rect 223210 8064 223266 8120
rect 223118 4256 223174 4312
rect 222566 1400 222622 1456
rect 223946 10104 224002 10160
rect 224038 9424 224094 9480
rect 224314 8336 224370 8392
rect 224682 8628 224738 8664
rect 224682 8608 224684 8628
rect 224684 8608 224736 8628
rect 224736 8608 224738 8628
rect 224590 8064 224646 8120
rect 223762 7928 223818 7984
rect 223486 6976 223542 7032
rect 223578 5616 223634 5672
rect 223762 5208 223818 5264
rect 223670 4800 223726 4856
rect 224866 8200 224922 8256
rect 223486 3712 223542 3768
rect 223578 3440 223634 3496
rect 224866 6704 224922 6760
rect 224590 5888 224646 5944
rect 225510 8628 225566 8664
rect 225510 8608 225512 8628
rect 225512 8608 225564 8628
rect 225564 8608 225566 8628
rect 225510 7828 225512 7848
rect 225512 7828 225564 7848
rect 225564 7828 225566 7848
rect 225510 7792 225566 7828
rect 223578 2488 223634 2544
rect 223486 1128 223542 1184
rect 224682 3984 224738 4040
rect 224498 2760 224554 2816
rect 224958 3712 225014 3768
rect 224866 2896 224922 2952
rect 224866 1944 224922 2000
rect 224222 1128 224278 1184
rect 223578 720 223634 776
rect 224774 720 224830 776
rect 220818 312 220874 368
rect 221094 312 221150 368
rect 225418 2624 225474 2680
rect 226246 8628 226302 8664
rect 226246 8608 226248 8628
rect 226248 8608 226300 8628
rect 226300 8608 226302 8628
rect 225970 7520 226026 7576
rect 225786 7112 225842 7168
rect 225970 7112 226026 7168
rect 226154 7928 226210 7984
rect 226246 7792 226302 7848
rect 226154 7520 226210 7576
rect 226246 6452 226302 6488
rect 226246 6432 226248 6452
rect 226248 6432 226300 6452
rect 226300 6432 226302 6452
rect 226246 5752 226302 5808
rect 227258 9016 227314 9072
rect 226982 8628 227038 8664
rect 226982 8608 226984 8628
rect 226984 8608 227036 8628
rect 227036 8608 227038 8628
rect 226706 6840 226762 6896
rect 225694 1128 225750 1184
rect 226430 1980 226432 2000
rect 226432 1980 226484 2000
rect 226484 1980 226486 2000
rect 226430 1944 226486 1980
rect 226522 1672 226578 1728
rect 226338 1400 226394 1456
rect 226522 1400 226578 1456
rect 226246 1264 226302 1320
rect 227074 2352 227130 2408
rect 228270 9444 228326 9480
rect 228270 9424 228272 9444
rect 228272 9424 228324 9444
rect 228324 9424 228326 9444
rect 228086 9152 228142 9208
rect 227350 7112 227406 7168
rect 227442 6976 227498 7032
rect 227626 6704 227682 6760
rect 227626 4528 227682 4584
rect 227902 5888 227958 5944
rect 227810 4564 227812 4584
rect 227812 4564 227864 4584
rect 227864 4564 227866 4584
rect 227810 4528 227866 4564
rect 227718 4256 227774 4312
rect 227626 3712 227682 3768
rect 227718 3576 227774 3632
rect 227626 3304 227682 3360
rect 228362 7928 228418 7984
rect 227902 2352 227958 2408
rect 227994 1128 228050 1184
rect 225970 584 226026 640
rect 227442 584 227498 640
rect 228546 3848 228602 3904
rect 229006 9444 229062 9480
rect 229006 9424 229008 9444
rect 229008 9424 229060 9444
rect 229060 9424 229062 9444
rect 229834 9444 229890 9480
rect 229834 9424 229836 9444
rect 229836 9424 229888 9444
rect 229888 9424 229890 9444
rect 229190 8628 229246 8664
rect 229190 8608 229192 8628
rect 229192 8608 229244 8628
rect 229244 8608 229246 8628
rect 228730 3576 228786 3632
rect 229006 5480 229062 5536
rect 229006 4120 229062 4176
rect 229742 6432 229798 6488
rect 229742 6160 229798 6216
rect 229926 3576 229982 3632
rect 229926 3168 229982 3224
rect 228638 1264 228694 1320
rect 230386 1672 230442 1728
rect 230018 1128 230074 1184
rect 228730 584 228786 640
rect 229466 584 229522 640
rect 230202 448 230258 504
rect 230386 448 230442 504
rect 230294 312 230350 368
rect 230938 8628 230994 8664
rect 230938 8608 230940 8628
rect 230940 8608 230992 8628
rect 230992 8608 230994 8628
rect 231950 9444 232006 9480
rect 231950 9424 231952 9444
rect 231952 9424 232004 9444
rect 232004 9424 232006 9444
rect 233422 9444 233478 9480
rect 233422 9424 233424 9444
rect 233424 9424 233476 9444
rect 233476 9424 233478 9444
rect 232778 9036 232834 9072
rect 232778 9016 232780 9036
rect 232780 9016 232832 9036
rect 232832 9016 232834 9036
rect 231674 8628 231730 8664
rect 231674 8608 231676 8628
rect 231676 8608 231728 8628
rect 231728 8608 231730 8628
rect 230202 176 230258 232
rect 231858 3596 231914 3632
rect 231858 3576 231860 3596
rect 231860 3576 231912 3596
rect 231912 3576 231914 3596
rect 232502 8744 232558 8800
rect 232594 8628 232650 8664
rect 232594 8608 232596 8628
rect 232596 8608 232648 8628
rect 232648 8608 232650 8628
rect 232318 8336 232374 8392
rect 231582 1128 231638 1184
rect 246210 10376 246266 10432
rect 234434 8628 234490 8664
rect 234434 8608 234436 8628
rect 234436 8608 234488 8628
rect 234488 8608 234490 8628
rect 234434 8336 234490 8392
rect 234894 8336 234950 8392
rect 232410 1128 232466 1184
rect 233146 1128 233202 1184
rect 235998 9444 236054 9480
rect 235998 9424 236000 9444
rect 236000 9424 236052 9444
rect 236052 9424 236054 9444
rect 235998 8744 236054 8800
rect 236274 8628 236330 8664
rect 236274 8608 236276 8628
rect 236276 8608 236328 8628
rect 236328 8608 236330 8628
rect 236826 9172 236882 9208
rect 236826 9152 236828 9172
rect 236828 9152 236880 9172
rect 236880 9152 236882 9172
rect 236734 9016 236790 9072
rect 237194 7520 237250 7576
rect 237545 9274 237601 9276
rect 237625 9274 237681 9276
rect 237705 9274 237761 9276
rect 237785 9274 237841 9276
rect 237545 9222 237591 9274
rect 237591 9222 237601 9274
rect 237625 9222 237655 9274
rect 237655 9222 237667 9274
rect 237667 9222 237681 9274
rect 237705 9222 237719 9274
rect 237719 9222 237731 9274
rect 237731 9222 237761 9274
rect 237785 9222 237795 9274
rect 237795 9222 237841 9274
rect 237545 9220 237601 9222
rect 237625 9220 237681 9222
rect 237705 9220 237761 9222
rect 237785 9220 237841 9222
rect 239954 10240 240010 10296
rect 240966 10240 241022 10296
rect 241242 10240 241298 10296
rect 242346 10240 242402 10296
rect 242898 10240 242954 10296
rect 243450 10240 243506 10296
rect 237545 8186 237601 8188
rect 237625 8186 237681 8188
rect 237705 8186 237761 8188
rect 237785 8186 237841 8188
rect 237545 8134 237591 8186
rect 237591 8134 237601 8186
rect 237625 8134 237655 8186
rect 237655 8134 237667 8186
rect 237667 8134 237681 8186
rect 237705 8134 237719 8186
rect 237719 8134 237731 8186
rect 237731 8134 237761 8186
rect 237785 8134 237795 8186
rect 237795 8134 237841 8186
rect 237545 8132 237601 8134
rect 237625 8132 237681 8134
rect 237705 8132 237761 8134
rect 237785 8132 237841 8134
rect 237378 8064 237434 8120
rect 237378 7520 237434 7576
rect 237545 7098 237601 7100
rect 237625 7098 237681 7100
rect 237705 7098 237761 7100
rect 237785 7098 237841 7100
rect 237545 7046 237591 7098
rect 237591 7046 237601 7098
rect 237625 7046 237655 7098
rect 237655 7046 237667 7098
rect 237667 7046 237681 7098
rect 237705 7046 237719 7098
rect 237719 7046 237731 7098
rect 237731 7046 237761 7098
rect 237785 7046 237795 7098
rect 237795 7046 237841 7098
rect 237545 7044 237601 7046
rect 237625 7044 237681 7046
rect 237705 7044 237761 7046
rect 237785 7044 237841 7046
rect 241518 6976 241574 7032
rect 237545 6010 237601 6012
rect 237625 6010 237681 6012
rect 237705 6010 237761 6012
rect 237785 6010 237841 6012
rect 237545 5958 237591 6010
rect 237591 5958 237601 6010
rect 237625 5958 237655 6010
rect 237655 5958 237667 6010
rect 237667 5958 237681 6010
rect 237705 5958 237719 6010
rect 237719 5958 237731 6010
rect 237731 5958 237761 6010
rect 237785 5958 237795 6010
rect 237795 5958 237841 6010
rect 237545 5956 237601 5958
rect 237625 5956 237681 5958
rect 237705 5956 237761 5958
rect 237785 5956 237841 5958
rect 239402 6432 239458 6488
rect 242530 7520 242586 7576
rect 241610 6568 241666 6624
rect 241794 6568 241850 6624
rect 239402 6160 239458 6216
rect 237286 5208 237342 5264
rect 237545 4922 237601 4924
rect 237625 4922 237681 4924
rect 237705 4922 237761 4924
rect 237785 4922 237841 4924
rect 237545 4870 237591 4922
rect 237591 4870 237601 4922
rect 237625 4870 237655 4922
rect 237655 4870 237667 4922
rect 237667 4870 237681 4922
rect 237705 4870 237719 4922
rect 237719 4870 237731 4922
rect 237731 4870 237761 4922
rect 237785 4870 237795 4922
rect 237795 4870 237841 4922
rect 237545 4868 237601 4870
rect 237625 4868 237681 4870
rect 237705 4868 237761 4870
rect 237785 4868 237841 4870
rect 237286 4256 237342 4312
rect 237545 3834 237601 3836
rect 237625 3834 237681 3836
rect 237705 3834 237761 3836
rect 237785 3834 237841 3836
rect 237545 3782 237591 3834
rect 237591 3782 237601 3834
rect 237625 3782 237655 3834
rect 237655 3782 237667 3834
rect 237667 3782 237681 3834
rect 237705 3782 237719 3834
rect 237719 3782 237731 3834
rect 237731 3782 237761 3834
rect 237785 3782 237795 3834
rect 237795 3782 237841 3834
rect 237545 3780 237601 3782
rect 237625 3780 237681 3782
rect 237705 3780 237761 3782
rect 237785 3780 237841 3782
rect 239402 3712 239458 3768
rect 235170 1128 235226 1184
rect 231858 584 231914 640
rect 233882 584 233938 640
rect 234618 584 234674 640
rect 235814 584 235870 640
rect 239402 3168 239458 3224
rect 237010 3032 237066 3088
rect 237545 2746 237601 2748
rect 237625 2746 237681 2748
rect 237705 2746 237761 2748
rect 237785 2746 237841 2748
rect 237545 2694 237591 2746
rect 237591 2694 237601 2746
rect 237625 2694 237655 2746
rect 237655 2694 237667 2746
rect 237667 2694 237681 2746
rect 237705 2694 237719 2746
rect 237719 2694 237731 2746
rect 237731 2694 237761 2746
rect 237785 2694 237795 2746
rect 237795 2694 237841 2746
rect 237545 2692 237601 2694
rect 237625 2692 237681 2694
rect 237705 2692 237761 2694
rect 237785 2692 237841 2694
rect 242898 5344 242954 5400
rect 242898 3168 242954 3224
rect 237545 1658 237601 1660
rect 237625 1658 237681 1660
rect 237705 1658 237761 1660
rect 237785 1658 237841 1660
rect 237545 1606 237591 1658
rect 237591 1606 237601 1658
rect 237625 1606 237655 1658
rect 237655 1606 237667 1658
rect 237667 1606 237681 1658
rect 237705 1606 237719 1658
rect 237719 1606 237731 1658
rect 237731 1606 237761 1658
rect 237785 1606 237795 1658
rect 237795 1606 237841 1658
rect 237545 1604 237601 1606
rect 237625 1604 237681 1606
rect 237705 1604 237761 1606
rect 237785 1604 237841 1606
rect 237378 1536 237434 1592
rect 236826 1128 236882 1184
rect 239954 584 240010 640
rect 240966 584 241022 640
rect 242806 1400 242862 1456
rect 242898 856 242954 912
rect 241242 584 241298 640
rect 241978 584 242034 640
rect 243082 4120 243138 4176
rect 244186 10240 244242 10296
rect 245014 10240 245070 10296
rect 244094 7112 244150 7168
rect 243542 1264 243598 1320
rect 243634 992 243690 1048
rect 243542 856 243598 912
rect 243450 584 243506 640
rect 236274 176 236330 232
rect 245198 8064 245254 8120
rect 246394 10240 246450 10296
rect 247130 10240 247186 10296
rect 247958 10240 248014 10296
rect 248694 10240 248750 10296
rect 249338 10240 249394 10296
rect 250166 10240 250222 10296
rect 251178 10240 251234 10296
rect 246210 5208 246266 5264
rect 246946 8064 247002 8120
rect 246670 7656 246726 7712
rect 250166 7928 250222 7984
rect 248970 6976 249026 7032
rect 248326 6452 248382 6488
rect 248326 6432 248328 6452
rect 248328 6432 248380 6452
rect 248380 6432 248382 6452
rect 246302 5072 246358 5128
rect 245934 4664 245990 4720
rect 245014 2216 245070 2272
rect 245474 3304 245530 3360
rect 247406 5616 247462 5672
rect 246854 2932 246856 2952
rect 246856 2932 246908 2952
rect 246908 2932 246910 2952
rect 246854 2896 246910 2932
rect 244186 584 244242 640
rect 245750 1400 245806 1456
rect 246670 1672 246726 1728
rect 244922 584 244978 640
rect 246946 1536 247002 1592
rect 246946 992 247002 1048
rect 247406 2216 247462 2272
rect 248326 5208 248382 5264
rect 248142 3460 248198 3496
rect 248142 3440 248144 3460
rect 248144 3440 248196 3460
rect 248196 3440 248198 3460
rect 248878 4256 248934 4312
rect 249062 4256 249118 4312
rect 248786 4120 248842 4176
rect 248694 3848 248750 3904
rect 249798 6704 249854 6760
rect 249062 3032 249118 3088
rect 249614 2760 249670 2816
rect 248418 2352 248474 2408
rect 247038 584 247094 640
rect 253846 10376 253902 10432
rect 251546 10240 251602 10296
rect 252282 10240 252338 10296
rect 253754 10240 253810 10296
rect 255042 10240 255098 10296
rect 255318 10240 255374 10296
rect 256422 10240 256478 10296
rect 256698 10240 256754 10296
rect 257710 10240 257766 10296
rect 258262 10240 258318 10296
rect 254122 7928 254178 7984
rect 252098 7420 252100 7440
rect 252100 7420 252152 7440
rect 252152 7420 252154 7440
rect 252098 7384 252154 7420
rect 251178 7284 251180 7304
rect 251180 7284 251232 7304
rect 251232 7284 251234 7304
rect 251178 7248 251234 7284
rect 251638 6296 251694 6352
rect 250350 5480 250406 5536
rect 250166 4256 250222 4312
rect 251086 4800 251142 4856
rect 250534 2932 250536 2952
rect 250536 2932 250588 2952
rect 250588 2932 250590 2952
rect 250534 2896 250590 2932
rect 249706 2488 249762 2544
rect 250994 3032 251050 3088
rect 251086 2624 251142 2680
rect 250810 1944 250866 2000
rect 249798 1400 249854 1456
rect 251270 1844 251272 1864
rect 251272 1844 251324 1864
rect 251324 1844 251326 1864
rect 251270 1808 251326 1844
rect 251362 1536 251418 1592
rect 248510 720 248566 776
rect 248418 584 248474 640
rect 250074 584 250130 640
rect 253478 6160 253534 6216
rect 252650 4256 252706 4312
rect 252558 1536 252614 1592
rect 252650 1400 252706 1456
rect 254306 5480 254362 5536
rect 254030 3596 254086 3632
rect 254030 3576 254032 3596
rect 254032 3576 254084 3596
rect 254084 3576 254086 3596
rect 255134 5344 255190 5400
rect 255134 4528 255190 4584
rect 254122 2216 254178 2272
rect 256422 4392 256478 4448
rect 256514 2896 256570 2952
rect 255226 1400 255282 1456
rect 255686 1128 255742 1184
rect 254858 584 254914 640
rect 253846 448 253902 504
rect 257526 1400 257582 1456
rect 259182 10240 259238 10296
rect 258170 6704 258226 6760
rect 258262 6024 258318 6080
rect 258262 5752 258318 5808
rect 258170 1536 258226 1592
rect 258446 3440 258502 3496
rect 258998 3168 259054 3224
rect 261758 10376 261814 10432
rect 259918 10240 259974 10296
rect 259550 6976 259606 7032
rect 260470 10240 260526 10296
rect 259274 3712 259330 3768
rect 259734 3304 259790 3360
rect 259826 2796 259828 2816
rect 259828 2796 259880 2816
rect 259880 2796 259882 2816
rect 259826 2760 259882 2796
rect 260010 4392 260066 4448
rect 260838 8064 260894 8120
rect 261850 10240 261906 10296
rect 262494 10240 262550 10296
rect 263322 10240 263378 10296
rect 260930 7112 260986 7168
rect 260930 6568 260986 6624
rect 260838 6024 260894 6080
rect 261022 5228 261078 5264
rect 261022 5208 261024 5228
rect 261024 5208 261076 5228
rect 261076 5208 261078 5228
rect 260838 4120 260894 4176
rect 258722 1944 258778 2000
rect 257802 1128 257858 1184
rect 258722 1400 258778 1456
rect 260470 2760 260526 2816
rect 260286 2100 260342 2136
rect 260286 2080 260288 2100
rect 260288 2080 260340 2100
rect 260340 2080 260342 2100
rect 260102 720 260158 776
rect 261666 7404 261722 7440
rect 261666 7384 261668 7404
rect 261668 7384 261720 7404
rect 261720 7384 261722 7404
rect 261758 6432 261814 6488
rect 262034 6432 262090 6488
rect 262218 7928 262274 7984
rect 262586 8200 262642 8256
rect 262310 7248 262366 7304
rect 262678 6704 262734 6760
rect 262126 2760 262182 2816
rect 262586 2760 262642 2816
rect 264334 10240 264390 10296
rect 263874 8356 263930 8392
rect 263874 8336 263876 8356
rect 263876 8336 263928 8356
rect 263928 8336 263930 8356
rect 263966 8200 264022 8256
rect 263230 7112 263286 7168
rect 263414 5616 263470 5672
rect 263230 4800 263286 4856
rect 266266 10376 266322 10432
rect 266174 10240 266230 10296
rect 260470 856 260526 912
rect 256790 584 256846 640
rect 258078 584 258134 640
rect 264886 8084 264942 8120
rect 264886 8064 264888 8084
rect 264888 8064 264940 8084
rect 264940 8064 264942 8084
rect 264886 7812 264942 7848
rect 264886 7792 264888 7812
rect 264888 7792 264940 7812
rect 264940 7792 264942 7812
rect 264794 5888 264850 5944
rect 265346 7656 265402 7712
rect 266358 6840 266414 6896
rect 265990 6704 266046 6760
rect 266358 5752 266414 5808
rect 268198 9988 268254 10024
rect 268198 9968 268200 9988
rect 268200 9968 268252 9988
rect 268252 9968 268254 9988
rect 267554 9460 267556 9480
rect 267556 9460 267608 9480
rect 267608 9460 267610 9480
rect 266266 3984 266322 4040
rect 266910 5244 266912 5264
rect 266912 5244 266964 5264
rect 266964 5244 266966 5264
rect 266910 5208 266966 5244
rect 267278 8372 267280 8392
rect 267280 8372 267332 8392
rect 267332 8372 267334 8392
rect 267278 8336 267334 8372
rect 267554 9424 267610 9460
rect 268106 9696 268162 9752
rect 267738 9424 267794 9480
rect 268014 9288 268070 9344
rect 268014 8336 268070 8392
rect 267738 7948 267794 7984
rect 267738 7928 267740 7948
rect 267740 7928 267792 7948
rect 267792 7928 267794 7948
rect 268014 7964 268016 7984
rect 268016 7964 268068 7984
rect 268068 7964 268070 7984
rect 268014 7928 268070 7964
rect 267922 7656 267978 7712
rect 267738 6996 267794 7032
rect 267738 6976 267740 6996
rect 267740 6976 267792 6996
rect 267792 6976 267794 6996
rect 267646 6704 267702 6760
rect 267646 5480 267702 5536
rect 267922 6976 267978 7032
rect 267922 6860 267978 6896
rect 267922 6840 267924 6860
rect 267924 6840 267976 6860
rect 267976 6840 267978 6860
rect 268290 8472 268346 8528
rect 268842 9696 268898 9752
rect 268290 8064 268346 8120
rect 268106 6432 268162 6488
rect 267278 4392 267334 4448
rect 267738 4936 267794 4992
rect 267738 4528 267794 4584
rect 267738 3732 267794 3768
rect 267738 3712 267740 3732
rect 267740 3712 267792 3732
rect 267792 3712 267794 3732
rect 267554 3440 267610 3496
rect 268014 3712 268070 3768
rect 268474 6024 268530 6080
rect 268290 5772 268346 5808
rect 268290 5752 268292 5772
rect 268292 5752 268344 5772
rect 268344 5752 268346 5772
rect 268474 5616 268530 5672
rect 268474 5072 268530 5128
rect 268290 4664 268346 4720
rect 268014 3440 268070 3496
rect 267922 3032 267978 3088
rect 267922 2796 267924 2816
rect 267924 2796 267976 2816
rect 267976 2796 267978 2816
rect 267922 2760 267978 2796
rect 267922 2624 267978 2680
rect 268474 4392 268530 4448
rect 268382 2488 268438 2544
rect 268750 9152 268806 9208
rect 268658 9016 268714 9072
rect 268658 7656 268714 7712
rect 272154 9968 272210 10024
rect 271343 9818 271399 9820
rect 271423 9818 271479 9820
rect 271503 9818 271559 9820
rect 271583 9818 271639 9820
rect 271343 9766 271389 9818
rect 271389 9766 271399 9818
rect 271423 9766 271453 9818
rect 271453 9766 271465 9818
rect 271465 9766 271479 9818
rect 271503 9766 271517 9818
rect 271517 9766 271529 9818
rect 271529 9766 271559 9818
rect 271583 9766 271593 9818
rect 271593 9766 271639 9818
rect 271343 9764 271399 9766
rect 271423 9764 271479 9766
rect 271503 9764 271559 9766
rect 271583 9764 271639 9766
rect 269026 8880 269082 8936
rect 268750 6296 268806 6352
rect 268658 5888 268714 5944
rect 268658 5480 268714 5536
rect 268566 3304 268622 3360
rect 267738 2080 267794 2136
rect 269026 6568 269082 6624
rect 268934 6160 268990 6216
rect 268842 6024 268898 6080
rect 269026 5908 269082 5944
rect 269026 5888 269028 5908
rect 269028 5888 269080 5908
rect 269080 5888 269082 5908
rect 269026 5208 269082 5264
rect 268934 4800 268990 4856
rect 268842 3576 268898 3632
rect 269486 5616 269542 5672
rect 270498 9580 270554 9616
rect 270498 9560 270500 9580
rect 270500 9560 270552 9580
rect 270552 9560 270554 9580
rect 271970 9424 272026 9480
rect 272154 9424 272210 9480
rect 270314 6160 270370 6216
rect 270498 5616 270554 5672
rect 271970 8880 272026 8936
rect 270682 6296 270738 6352
rect 271343 8730 271399 8732
rect 271423 8730 271479 8732
rect 271503 8730 271559 8732
rect 271583 8730 271639 8732
rect 271343 8678 271389 8730
rect 271389 8678 271399 8730
rect 271423 8678 271453 8730
rect 271453 8678 271465 8730
rect 271465 8678 271479 8730
rect 271503 8678 271517 8730
rect 271517 8678 271529 8730
rect 271529 8678 271559 8730
rect 271583 8678 271593 8730
rect 271593 8678 271639 8730
rect 271343 8676 271399 8678
rect 271423 8676 271479 8678
rect 271503 8676 271559 8678
rect 271583 8676 271639 8678
rect 271786 8200 271842 8256
rect 272154 8084 272210 8120
rect 272154 8064 272156 8084
rect 272156 8064 272208 8084
rect 272208 8064 272210 8084
rect 270958 6704 271014 6760
rect 270774 3984 270830 4040
rect 271786 7928 271842 7984
rect 271142 7656 271198 7712
rect 271786 7656 271842 7712
rect 271343 7642 271399 7644
rect 271423 7642 271479 7644
rect 271503 7642 271559 7644
rect 271583 7642 271639 7644
rect 271343 7590 271389 7642
rect 271389 7590 271399 7642
rect 271423 7590 271453 7642
rect 271453 7590 271465 7642
rect 271465 7590 271479 7642
rect 271503 7590 271517 7642
rect 271517 7590 271529 7642
rect 271529 7590 271559 7642
rect 271583 7590 271593 7642
rect 271593 7590 271639 7642
rect 271343 7588 271399 7590
rect 271423 7588 271479 7590
rect 271503 7588 271559 7590
rect 271583 7588 271639 7590
rect 271142 7540 271198 7576
rect 271142 7520 271144 7540
rect 271144 7520 271196 7540
rect 271196 7520 271198 7540
rect 272154 7928 272210 7984
rect 271970 7384 272026 7440
rect 272062 6568 272118 6624
rect 271343 6554 271399 6556
rect 271423 6554 271479 6556
rect 271503 6554 271559 6556
rect 271583 6554 271639 6556
rect 271343 6502 271389 6554
rect 271389 6502 271399 6554
rect 271423 6502 271453 6554
rect 271453 6502 271465 6554
rect 271465 6502 271479 6554
rect 271503 6502 271517 6554
rect 271517 6502 271529 6554
rect 271529 6502 271559 6554
rect 271583 6502 271593 6554
rect 271593 6502 271639 6554
rect 271343 6500 271399 6502
rect 271423 6500 271479 6502
rect 271503 6500 271559 6502
rect 271583 6500 271639 6502
rect 271142 6432 271198 6488
rect 271878 6432 271934 6488
rect 271326 6296 271382 6352
rect 271326 6024 271382 6080
rect 271694 6024 271750 6080
rect 271142 5888 271198 5944
rect 271142 5516 271144 5536
rect 271144 5516 271196 5536
rect 271196 5516 271198 5536
rect 271142 5480 271198 5516
rect 270682 2796 270684 2816
rect 270684 2796 270736 2816
rect 270736 2796 270738 2816
rect 270682 2760 270738 2796
rect 268842 1808 268898 1864
rect 268014 1264 268070 1320
rect 267922 856 267978 912
rect 267738 720 267794 776
rect 269854 1556 269910 1592
rect 269854 1536 269856 1556
rect 269856 1536 269908 1556
rect 269908 1536 269910 1556
rect 261114 584 261170 640
rect 262862 584 262918 640
rect 263322 584 263378 640
rect 264334 584 264390 640
rect 264978 584 265034 640
rect 265806 584 265862 640
rect 266358 584 266414 640
rect 266910 584 266966 640
rect 267646 584 267702 640
rect 268382 584 268438 640
rect 269762 584 269818 640
rect 255962 312 256018 368
rect 271142 4392 271198 4448
rect 271343 5466 271399 5468
rect 271423 5466 271479 5468
rect 271503 5466 271559 5468
rect 271583 5466 271639 5468
rect 271343 5414 271389 5466
rect 271389 5414 271399 5466
rect 271423 5414 271453 5466
rect 271453 5414 271465 5466
rect 271465 5414 271479 5466
rect 271503 5414 271517 5466
rect 271517 5414 271529 5466
rect 271529 5414 271559 5466
rect 271583 5414 271593 5466
rect 271593 5414 271639 5466
rect 271343 5412 271399 5414
rect 271423 5412 271479 5414
rect 271503 5412 271559 5414
rect 271583 5412 271639 5414
rect 271786 5516 271788 5536
rect 271788 5516 271840 5536
rect 271840 5516 271842 5536
rect 271786 5480 271842 5516
rect 271786 5344 271842 5400
rect 271786 4936 271842 4992
rect 271343 4378 271399 4380
rect 271423 4378 271479 4380
rect 271503 4378 271559 4380
rect 271583 4378 271639 4380
rect 271343 4326 271389 4378
rect 271389 4326 271399 4378
rect 271423 4326 271453 4378
rect 271453 4326 271465 4378
rect 271465 4326 271479 4378
rect 271503 4326 271517 4378
rect 271517 4326 271529 4378
rect 271529 4326 271559 4378
rect 271583 4326 271593 4378
rect 271593 4326 271639 4378
rect 271343 4324 271399 4326
rect 271423 4324 271479 4326
rect 271503 4324 271559 4326
rect 271583 4324 271639 4326
rect 271786 4256 271842 4312
rect 271694 4120 271750 4176
rect 271142 3340 271144 3360
rect 271144 3340 271196 3360
rect 271196 3340 271198 3360
rect 271142 3304 271198 3340
rect 271343 3290 271399 3292
rect 271423 3290 271479 3292
rect 271503 3290 271559 3292
rect 271583 3290 271639 3292
rect 271343 3238 271389 3290
rect 271389 3238 271399 3290
rect 271423 3238 271453 3290
rect 271453 3238 271465 3290
rect 271465 3238 271479 3290
rect 271503 3238 271517 3290
rect 271517 3238 271529 3290
rect 271529 3238 271559 3290
rect 271583 3238 271593 3290
rect 271593 3238 271639 3290
rect 271343 3236 271399 3238
rect 271423 3236 271479 3238
rect 271503 3236 271559 3238
rect 271583 3236 271639 3238
rect 271970 4936 272026 4992
rect 272154 3848 272210 3904
rect 272154 3576 272210 3632
rect 271142 3168 271198 3224
rect 271786 3168 271842 3224
rect 271234 2760 271290 2816
rect 271142 2216 271198 2272
rect 271343 2202 271399 2204
rect 271423 2202 271479 2204
rect 271503 2202 271559 2204
rect 271583 2202 271639 2204
rect 271343 2150 271389 2202
rect 271389 2150 271399 2202
rect 271423 2150 271453 2202
rect 271453 2150 271465 2202
rect 271465 2150 271479 2202
rect 271503 2150 271517 2202
rect 271517 2150 271529 2202
rect 271529 2150 271559 2202
rect 271583 2150 271593 2202
rect 271593 2150 271639 2202
rect 271343 2148 271399 2150
rect 271423 2148 271479 2150
rect 271503 2148 271559 2150
rect 271583 2148 271639 2150
rect 271970 2080 272026 2136
rect 272062 1944 272118 2000
rect 271970 1536 272026 1592
rect 271970 1264 272026 1320
rect 271343 1114 271399 1116
rect 271423 1114 271479 1116
rect 271503 1114 271559 1116
rect 271583 1114 271639 1116
rect 271343 1062 271389 1114
rect 271389 1062 271399 1114
rect 271423 1062 271453 1114
rect 271453 1062 271465 1114
rect 271465 1062 271479 1114
rect 271503 1062 271517 1114
rect 271517 1062 271529 1114
rect 271529 1062 271559 1114
rect 271583 1062 271593 1114
rect 271593 1062 271639 1114
rect 271343 1060 271399 1062
rect 271423 1060 271479 1062
rect 271503 1060 271559 1062
rect 271583 1060 271639 1062
rect 271970 856 272026 912
rect 272154 1536 272210 1592
rect 270774 584 270830 640
rect 270314 312 270370 368
rect 213366 40 213422 96
rect 231398 40 231454 96
<< metal3 >>
rect 52586 10508 52592 10572
rect 52656 10570 52662 10572
rect 53097 10570 53163 10573
rect 81617 10572 81683 10573
rect 81566 10570 81572 10572
rect 52656 10568 53163 10570
rect 52656 10512 53102 10568
rect 53158 10512 53163 10568
rect 52656 10510 53163 10512
rect 81526 10510 81572 10570
rect 81636 10568 81683 10572
rect 81678 10512 81683 10568
rect 52656 10508 52662 10510
rect 53097 10507 53163 10510
rect 81566 10508 81572 10510
rect 81636 10508 81683 10512
rect 82302 10508 82308 10572
rect 82372 10570 82378 10572
rect 82629 10570 82695 10573
rect 86769 10572 86835 10573
rect 86718 10570 86724 10572
rect 82372 10568 82695 10570
rect 82372 10512 82634 10568
rect 82690 10512 82695 10568
rect 82372 10510 82695 10512
rect 86678 10510 86724 10570
rect 86788 10568 86835 10572
rect 86830 10512 86835 10568
rect 82372 10508 82378 10510
rect 81617 10507 81683 10508
rect 82629 10507 82695 10510
rect 86718 10508 86724 10510
rect 86788 10508 86835 10512
rect 147622 10508 147628 10572
rect 147692 10570 147698 10572
rect 148409 10570 148475 10573
rect 172237 10572 172303 10573
rect 172186 10570 172192 10572
rect 147692 10568 148475 10570
rect 147692 10512 148414 10568
rect 148470 10512 148475 10568
rect 147692 10510 148475 10512
rect 172146 10510 172192 10570
rect 172256 10568 172303 10572
rect 172298 10512 172303 10568
rect 147692 10508 147698 10510
rect 86769 10507 86835 10508
rect 148409 10507 148475 10510
rect 172186 10508 172192 10510
rect 172256 10508 172303 10512
rect 179546 10508 179552 10572
rect 179616 10570 179622 10572
rect 180517 10570 180583 10573
rect 179616 10568 180583 10570
rect 179616 10512 180522 10568
rect 180578 10512 180583 10568
rect 179616 10510 180583 10512
rect 179616 10508 179622 10510
rect 172237 10507 172303 10508
rect 180517 10507 180583 10510
rect 207790 10508 207796 10572
rect 207860 10570 207866 10572
rect 208301 10570 208367 10573
rect 207860 10568 208367 10570
rect 207860 10512 208306 10568
rect 208362 10512 208367 10568
rect 207860 10510 208367 10512
rect 207860 10508 207866 10510
rect 208301 10507 208367 10510
rect 212942 10508 212948 10572
rect 213012 10570 213018 10572
rect 213453 10570 213519 10573
rect 213012 10568 213519 10570
rect 213012 10512 213458 10568
rect 213514 10512 213519 10568
rect 213012 10510 213519 10512
rect 213012 10508 213018 10510
rect 213453 10507 213519 10510
rect 218094 10508 218100 10572
rect 218164 10570 218170 10572
rect 218605 10570 218671 10573
rect 223481 10570 223547 10573
rect 218164 10568 218671 10570
rect 218164 10512 218610 10568
rect 218666 10512 218671 10568
rect 218164 10510 218671 10512
rect 218164 10508 218170 10510
rect 218605 10507 218671 10510
rect 220862 10568 223547 10570
rect 220862 10512 223486 10568
rect 223542 10512 223547 10568
rect 220862 10510 223547 10512
rect 72049 10436 72115 10437
rect 71998 10434 72004 10436
rect 71958 10374 72004 10434
rect 72068 10432 72115 10436
rect 72110 10376 72115 10432
rect 71998 10372 72004 10374
rect 72068 10372 72115 10376
rect 72049 10371 72115 10372
rect 96613 10436 96679 10437
rect 96613 10432 96660 10436
rect 96724 10434 96730 10436
rect 96613 10376 96618 10432
rect 96613 10372 96660 10376
rect 96724 10374 96770 10434
rect 96724 10372 96730 10374
rect 125266 10372 125272 10436
rect 125336 10434 125342 10436
rect 125593 10434 125659 10437
rect 154297 10436 154363 10437
rect 154246 10434 154252 10436
rect 125336 10432 125659 10434
rect 125336 10376 125598 10432
rect 125654 10376 125659 10432
rect 125336 10374 125659 10376
rect 154206 10374 154252 10434
rect 154316 10432 154363 10436
rect 154358 10376 154363 10432
rect 125336 10372 125342 10374
rect 96613 10371 96679 10372
rect 125593 10371 125659 10374
rect 154246 10372 154252 10374
rect 154316 10372 154363 10376
rect 172922 10372 172928 10436
rect 172992 10434 172998 10436
rect 173985 10434 174051 10437
rect 172992 10432 174051 10434
rect 172992 10376 173990 10432
rect 174046 10376 174051 10432
rect 172992 10374 174051 10376
rect 172992 10372 172998 10374
rect 154297 10371 154363 10372
rect 173985 10371 174051 10374
rect 181018 10372 181024 10436
rect 181088 10434 181094 10436
rect 181805 10434 181871 10437
rect 181088 10432 181871 10434
rect 181088 10376 181810 10432
rect 181866 10376 181871 10432
rect 181088 10374 181871 10376
rect 181088 10372 181094 10374
rect 181805 10371 181871 10374
rect 190586 10372 190592 10436
rect 190656 10434 190662 10436
rect 191281 10434 191347 10437
rect 192845 10436 192911 10437
rect 202413 10436 202479 10437
rect 190656 10432 191347 10434
rect 190656 10376 191286 10432
rect 191342 10376 191347 10432
rect 190656 10374 191347 10376
rect 190656 10372 190662 10374
rect 191281 10371 191347 10374
rect 192794 10372 192800 10436
rect 192864 10434 192911 10436
rect 192864 10432 192956 10434
rect 192906 10376 192956 10432
rect 192864 10374 192956 10376
rect 192864 10372 192911 10374
rect 202362 10372 202368 10436
rect 202432 10434 202479 10436
rect 202432 10432 202524 10434
rect 202474 10376 202524 10432
rect 202432 10374 202524 10376
rect 202432 10372 202479 10374
rect 209998 10372 210004 10436
rect 210068 10434 210074 10436
rect 210877 10434 210943 10437
rect 210068 10432 210943 10434
rect 210068 10376 210882 10432
rect 210938 10376 210943 10432
rect 210068 10374 210943 10376
rect 210068 10372 210074 10374
rect 192845 10371 192911 10372
rect 202413 10371 202479 10372
rect 210877 10371 210943 10374
rect 216581 10434 216647 10437
rect 220862 10434 220922 10510
rect 223481 10507 223547 10510
rect 216581 10432 220922 10434
rect 216581 10376 216586 10432
rect 216642 10376 220922 10432
rect 216581 10374 220922 10376
rect 216581 10371 216647 10374
rect 221038 10372 221044 10436
rect 221108 10434 221114 10436
rect 221825 10434 221891 10437
rect 221108 10432 221891 10434
rect 221108 10376 221830 10432
rect 221886 10376 221891 10432
rect 221108 10374 221891 10376
rect 221108 10372 221114 10374
rect 221825 10371 221891 10374
rect 245602 10372 245608 10436
rect 245672 10434 245678 10436
rect 246205 10434 246271 10437
rect 245672 10432 246271 10434
rect 245672 10376 246210 10432
rect 246266 10376 246271 10432
rect 245672 10374 246271 10376
rect 245672 10372 245678 10374
rect 246205 10371 246271 10374
rect 252962 10372 252968 10436
rect 253032 10434 253038 10436
rect 253841 10434 253907 10437
rect 253032 10432 253907 10434
rect 253032 10376 253846 10432
rect 253902 10376 253907 10432
rect 253032 10374 253907 10376
rect 253032 10372 253038 10374
rect 253841 10371 253907 10374
rect 261058 10372 261064 10436
rect 261128 10434 261134 10436
rect 261753 10434 261819 10437
rect 261128 10432 261819 10434
rect 261128 10376 261758 10432
rect 261814 10376 261819 10432
rect 261128 10374 261819 10376
rect 261128 10372 261134 10374
rect 261753 10371 261819 10374
rect 265474 10372 265480 10436
rect 265544 10434 265550 10436
rect 266261 10434 266327 10437
rect 265544 10432 266327 10434
rect 265544 10376 266266 10432
rect 266322 10376 266327 10432
rect 265544 10374 266327 10376
rect 265544 10372 265550 10374
rect 266261 10371 266327 10374
rect 31702 10236 31708 10300
rect 31772 10298 31778 10300
rect 32489 10298 32555 10301
rect 31772 10296 32555 10298
rect 31772 10240 32494 10296
rect 32550 10240 32555 10296
rect 31772 10238 32555 10240
rect 31772 10236 31778 10238
rect 32489 10235 32555 10238
rect 34922 10236 34928 10300
rect 34992 10298 34998 10300
rect 35157 10298 35223 10301
rect 34992 10296 35223 10298
rect 34992 10240 35162 10296
rect 35218 10240 35223 10296
rect 34992 10238 35223 10240
rect 34992 10236 34998 10238
rect 35157 10235 35223 10238
rect 35617 10300 35683 10301
rect 35617 10296 35664 10300
rect 35728 10298 35734 10300
rect 36261 10298 36327 10301
rect 36394 10298 36400 10300
rect 35617 10240 35622 10296
rect 35617 10236 35664 10240
rect 35728 10238 35774 10298
rect 36261 10296 36400 10298
rect 36261 10240 36266 10296
rect 36322 10240 36400 10296
rect 36261 10238 36400 10240
rect 35728 10236 35734 10238
rect 35617 10235 35683 10236
rect 36261 10235 36327 10238
rect 36394 10236 36400 10238
rect 36464 10236 36470 10300
rect 36905 10298 36971 10301
rect 37130 10298 37136 10300
rect 36905 10296 37136 10298
rect 36905 10240 36910 10296
rect 36966 10240 37136 10296
rect 36905 10238 37136 10240
rect 36905 10235 36971 10238
rect 37130 10236 37136 10238
rect 37200 10236 37206 10300
rect 37866 10236 37872 10300
rect 37936 10298 37942 10300
rect 38101 10298 38167 10301
rect 37936 10296 38167 10298
rect 37936 10240 38106 10296
rect 38162 10240 38167 10296
rect 37936 10238 38167 10240
rect 37936 10236 37942 10238
rect 38101 10235 38167 10238
rect 38602 10236 38608 10300
rect 38672 10298 38678 10300
rect 38837 10298 38903 10301
rect 38672 10296 38903 10298
rect 38672 10240 38842 10296
rect 38898 10240 38903 10296
rect 38672 10238 38903 10240
rect 38672 10236 38678 10238
rect 38837 10235 38903 10238
rect 39338 10236 39344 10300
rect 39408 10298 39414 10300
rect 39481 10298 39547 10301
rect 39408 10296 39547 10298
rect 39408 10240 39486 10296
rect 39542 10240 39547 10296
rect 39408 10238 39547 10240
rect 39408 10236 39414 10238
rect 39481 10235 39547 10238
rect 40074 10236 40080 10300
rect 40144 10298 40150 10300
rect 40309 10298 40375 10301
rect 40144 10296 40375 10298
rect 40144 10240 40314 10296
rect 40370 10240 40375 10296
rect 40144 10238 40375 10240
rect 40144 10236 40150 10238
rect 40309 10235 40375 10238
rect 40769 10300 40835 10301
rect 40769 10296 40816 10300
rect 40880 10298 40886 10300
rect 41413 10298 41479 10301
rect 41546 10298 41552 10300
rect 40769 10240 40774 10296
rect 40769 10236 40816 10240
rect 40880 10238 40926 10298
rect 41413 10296 41552 10298
rect 41413 10240 41418 10296
rect 41474 10240 41552 10296
rect 41413 10238 41552 10240
rect 40880 10236 40886 10238
rect 40769 10235 40835 10236
rect 41413 10235 41479 10238
rect 41546 10236 41552 10238
rect 41616 10236 41622 10300
rect 42057 10298 42123 10301
rect 42282 10298 42288 10300
rect 42057 10296 42288 10298
rect 42057 10240 42062 10296
rect 42118 10240 42288 10296
rect 42057 10238 42288 10240
rect 42057 10235 42123 10238
rect 42282 10236 42288 10238
rect 42352 10236 42358 10300
rect 43018 10236 43024 10300
rect 43088 10298 43094 10300
rect 43253 10298 43319 10301
rect 43088 10296 43319 10298
rect 43088 10240 43258 10296
rect 43314 10240 43319 10296
rect 43088 10238 43319 10240
rect 43088 10236 43094 10238
rect 43253 10235 43319 10238
rect 43754 10236 43760 10300
rect 43824 10298 43830 10300
rect 43989 10298 44055 10301
rect 43824 10296 44055 10298
rect 43824 10240 43994 10296
rect 44050 10240 44055 10296
rect 43824 10238 44055 10240
rect 43824 10236 43830 10238
rect 43989 10235 44055 10238
rect 44490 10236 44496 10300
rect 44560 10298 44566 10300
rect 44633 10298 44699 10301
rect 44560 10296 44699 10298
rect 44560 10240 44638 10296
rect 44694 10240 44699 10296
rect 44560 10238 44699 10240
rect 44560 10236 44566 10238
rect 44633 10235 44699 10238
rect 45226 10236 45232 10300
rect 45296 10298 45302 10300
rect 45461 10298 45527 10301
rect 45296 10296 45527 10298
rect 45296 10240 45466 10296
rect 45522 10240 45527 10296
rect 45296 10238 45527 10240
rect 45296 10236 45302 10238
rect 45461 10235 45527 10238
rect 45921 10300 45987 10301
rect 45921 10296 45968 10300
rect 46032 10298 46038 10300
rect 46565 10298 46631 10301
rect 46698 10298 46704 10300
rect 45921 10240 45926 10296
rect 45921 10236 45968 10240
rect 46032 10238 46078 10298
rect 46565 10296 46704 10298
rect 46565 10240 46570 10296
rect 46626 10240 46704 10296
rect 46565 10238 46704 10240
rect 46032 10236 46038 10238
rect 45921 10235 45987 10236
rect 46565 10235 46631 10238
rect 46698 10236 46704 10238
rect 46768 10236 46774 10300
rect 47209 10298 47275 10301
rect 48221 10300 48287 10301
rect 47434 10298 47440 10300
rect 47209 10296 47440 10298
rect 47209 10240 47214 10296
rect 47270 10240 47440 10296
rect 47209 10238 47440 10240
rect 47209 10235 47275 10238
rect 47434 10236 47440 10238
rect 47504 10236 47510 10300
rect 48170 10298 48176 10300
rect 48130 10238 48176 10298
rect 48240 10296 48287 10300
rect 48282 10240 48287 10296
rect 48170 10236 48176 10238
rect 48240 10236 48287 10240
rect 48906 10236 48912 10300
rect 48976 10298 48982 10300
rect 49141 10298 49207 10301
rect 48976 10296 49207 10298
rect 48976 10240 49146 10296
rect 49202 10240 49207 10296
rect 48976 10238 49207 10240
rect 48976 10236 48982 10238
rect 48221 10235 48287 10236
rect 49141 10235 49207 10238
rect 49642 10236 49648 10300
rect 49712 10298 49718 10300
rect 49785 10298 49851 10301
rect 49712 10296 49851 10298
rect 49712 10240 49790 10296
rect 49846 10240 49851 10296
rect 49712 10238 49851 10240
rect 49712 10236 49718 10238
rect 49785 10235 49851 10238
rect 50378 10236 50384 10300
rect 50448 10298 50454 10300
rect 50613 10298 50679 10301
rect 50448 10296 50679 10298
rect 50448 10240 50618 10296
rect 50674 10240 50679 10296
rect 50448 10238 50679 10240
rect 50448 10236 50454 10238
rect 50613 10235 50679 10238
rect 51114 10236 51120 10300
rect 51184 10298 51190 10300
rect 51349 10298 51415 10301
rect 51184 10296 51415 10298
rect 51184 10240 51354 10296
rect 51410 10240 51415 10296
rect 51184 10238 51415 10240
rect 51184 10236 51190 10238
rect 51349 10235 51415 10238
rect 51850 10236 51856 10300
rect 51920 10298 51926 10300
rect 52085 10298 52151 10301
rect 53281 10300 53347 10301
rect 53281 10298 53328 10300
rect 51920 10296 52151 10298
rect 51920 10240 52090 10296
rect 52146 10240 52151 10296
rect 51920 10238 52151 10240
rect 53236 10296 53328 10298
rect 53236 10240 53286 10296
rect 53236 10238 53328 10240
rect 51920 10236 51926 10238
rect 52085 10235 52151 10238
rect 53281 10236 53328 10238
rect 53392 10236 53398 10300
rect 53833 10298 53899 10301
rect 54845 10300 54911 10301
rect 54058 10298 54064 10300
rect 53833 10296 54064 10298
rect 53833 10240 53838 10296
rect 53894 10240 54064 10296
rect 53833 10238 54064 10240
rect 53281 10235 53347 10236
rect 53833 10235 53899 10238
rect 54058 10236 54064 10238
rect 54128 10236 54134 10300
rect 54794 10236 54800 10300
rect 54864 10298 54911 10300
rect 54864 10296 54956 10298
rect 54906 10240 54956 10296
rect 54864 10238 54956 10240
rect 54864 10236 54911 10238
rect 55530 10236 55536 10300
rect 55600 10298 55606 10300
rect 55673 10298 55739 10301
rect 55600 10296 55739 10298
rect 55600 10240 55678 10296
rect 55734 10240 55739 10296
rect 55600 10238 55739 10240
rect 55600 10236 55606 10238
rect 54845 10235 54911 10236
rect 55673 10235 55739 10238
rect 56266 10236 56272 10300
rect 56336 10298 56342 10300
rect 56501 10298 56567 10301
rect 56336 10296 56567 10298
rect 56336 10240 56506 10296
rect 56562 10240 56567 10296
rect 56336 10238 56567 10240
rect 56336 10236 56342 10238
rect 56501 10235 56567 10238
rect 57002 10236 57008 10300
rect 57072 10298 57078 10300
rect 57329 10298 57395 10301
rect 57789 10300 57855 10301
rect 57072 10296 57395 10298
rect 57072 10240 57334 10296
rect 57390 10240 57395 10296
rect 57072 10238 57395 10240
rect 57072 10236 57078 10238
rect 57329 10235 57395 10238
rect 57738 10236 57744 10300
rect 57808 10298 57855 10300
rect 57808 10296 57900 10298
rect 57850 10240 57900 10296
rect 57808 10238 57900 10240
rect 57808 10236 57855 10238
rect 58474 10236 58480 10300
rect 58544 10298 58550 10300
rect 58801 10298 58867 10301
rect 59261 10300 59327 10301
rect 58544 10296 58867 10298
rect 58544 10240 58806 10296
rect 58862 10240 58867 10296
rect 58544 10238 58867 10240
rect 58544 10236 58550 10238
rect 57789 10235 57855 10236
rect 58801 10235 58867 10238
rect 59210 10236 59216 10300
rect 59280 10298 59327 10300
rect 59280 10296 59372 10298
rect 59322 10240 59372 10296
rect 59280 10238 59372 10240
rect 59280 10236 59327 10238
rect 59946 10236 59952 10300
rect 60016 10298 60022 10300
rect 60273 10298 60339 10301
rect 60016 10296 60339 10298
rect 60016 10240 60278 10296
rect 60334 10240 60339 10296
rect 60016 10238 60339 10240
rect 60016 10236 60022 10238
rect 59261 10235 59327 10236
rect 60273 10235 60339 10238
rect 60682 10236 60688 10300
rect 60752 10298 60758 10300
rect 61009 10298 61075 10301
rect 60752 10296 61075 10298
rect 60752 10240 61014 10296
rect 61070 10240 61075 10296
rect 60752 10238 61075 10240
rect 60752 10236 60758 10238
rect 61009 10235 61075 10238
rect 61418 10236 61424 10300
rect 61488 10298 61494 10300
rect 61745 10298 61811 10301
rect 61488 10296 61811 10298
rect 61488 10240 61750 10296
rect 61806 10240 61811 10296
rect 61488 10238 61811 10240
rect 61488 10236 61494 10238
rect 61745 10235 61811 10238
rect 62154 10236 62160 10300
rect 62224 10298 62230 10300
rect 62481 10298 62547 10301
rect 62224 10296 62547 10298
rect 62224 10240 62486 10296
rect 62542 10240 62547 10296
rect 62224 10238 62547 10240
rect 62224 10236 62230 10238
rect 62481 10235 62547 10238
rect 62890 10236 62896 10300
rect 62960 10298 62966 10300
rect 63401 10298 63467 10301
rect 62960 10296 63467 10298
rect 62960 10240 63406 10296
rect 63462 10240 63467 10296
rect 62960 10238 63467 10240
rect 62960 10236 62966 10238
rect 63401 10235 63467 10238
rect 63626 10236 63632 10300
rect 63696 10298 63702 10300
rect 63953 10298 64019 10301
rect 63696 10296 64019 10298
rect 63696 10240 63958 10296
rect 64014 10240 64019 10296
rect 63696 10238 64019 10240
rect 63696 10236 63702 10238
rect 63953 10235 64019 10238
rect 64362 10236 64368 10300
rect 64432 10298 64438 10300
rect 64689 10298 64755 10301
rect 64432 10296 64755 10298
rect 64432 10240 64694 10296
rect 64750 10240 64755 10296
rect 64432 10238 64755 10240
rect 64432 10236 64438 10238
rect 64689 10235 64755 10238
rect 65098 10236 65104 10300
rect 65168 10298 65174 10300
rect 65517 10298 65583 10301
rect 65885 10300 65951 10301
rect 65168 10296 65583 10298
rect 65168 10240 65522 10296
rect 65578 10240 65583 10296
rect 65168 10238 65583 10240
rect 65168 10236 65174 10238
rect 65517 10235 65583 10238
rect 65834 10236 65840 10300
rect 65904 10298 65951 10300
rect 65904 10296 65996 10298
rect 65946 10240 65996 10296
rect 65904 10238 65996 10240
rect 65904 10236 65951 10238
rect 66570 10236 66576 10300
rect 66640 10298 66646 10300
rect 67173 10298 67239 10301
rect 66640 10296 67239 10298
rect 66640 10240 67178 10296
rect 67234 10240 67239 10296
rect 66640 10238 67239 10240
rect 66640 10236 66646 10238
rect 65885 10235 65951 10236
rect 67173 10235 67239 10238
rect 89662 10236 89668 10300
rect 89732 10298 89738 10300
rect 90357 10298 90423 10301
rect 103237 10300 103303 10301
rect 89732 10296 90423 10298
rect 89732 10240 90362 10296
rect 90418 10240 90423 10296
rect 89732 10238 90423 10240
rect 89732 10236 89738 10238
rect 90357 10235 90423 10238
rect 103186 10236 103192 10300
rect 103256 10298 103303 10300
rect 103881 10300 103947 10301
rect 104709 10300 104775 10301
rect 103256 10296 103348 10298
rect 103298 10240 103348 10296
rect 103256 10238 103348 10240
rect 103881 10296 103928 10300
rect 103992 10298 103998 10300
rect 104658 10298 104664 10300
rect 103881 10240 103886 10296
rect 103256 10236 103303 10238
rect 103237 10235 103303 10236
rect 103881 10236 103928 10240
rect 103992 10238 104038 10298
rect 104618 10238 104664 10298
rect 104728 10296 104775 10300
rect 104770 10240 104775 10296
rect 103992 10236 103998 10238
rect 104658 10236 104664 10238
rect 104728 10236 104775 10240
rect 105394 10236 105400 10300
rect 105464 10298 105470 10300
rect 105629 10298 105695 10301
rect 105464 10296 105695 10298
rect 105464 10240 105634 10296
rect 105690 10240 105695 10296
rect 105464 10238 105695 10240
rect 105464 10236 105470 10238
rect 103881 10235 103947 10236
rect 104709 10235 104775 10236
rect 105629 10235 105695 10238
rect 106130 10236 106136 10300
rect 106200 10298 106206 10300
rect 106273 10298 106339 10301
rect 106200 10296 106339 10298
rect 106200 10240 106278 10296
rect 106334 10240 106339 10296
rect 106200 10238 106339 10240
rect 106200 10236 106206 10238
rect 106273 10235 106339 10238
rect 106866 10236 106872 10300
rect 106936 10298 106942 10300
rect 107193 10298 107259 10301
rect 106936 10296 107259 10298
rect 106936 10240 107198 10296
rect 107254 10240 107259 10296
rect 106936 10238 107259 10240
rect 106936 10236 106942 10238
rect 107193 10235 107259 10238
rect 107602 10236 107608 10300
rect 107672 10298 107678 10300
rect 107745 10298 107811 10301
rect 108389 10300 108455 10301
rect 108338 10298 108344 10300
rect 107672 10296 107811 10298
rect 107672 10240 107750 10296
rect 107806 10240 107811 10296
rect 107672 10238 107811 10240
rect 108298 10238 108344 10298
rect 108408 10296 108455 10300
rect 108450 10240 108455 10296
rect 107672 10236 107678 10238
rect 107745 10235 107811 10238
rect 108338 10236 108344 10238
rect 108408 10236 108455 10240
rect 108389 10235 108455 10236
rect 109033 10300 109099 10301
rect 109033 10296 109080 10300
rect 109144 10298 109150 10300
rect 109033 10240 109038 10296
rect 109033 10236 109080 10240
rect 109144 10238 109190 10298
rect 109144 10236 109150 10238
rect 109810 10236 109816 10300
rect 109880 10298 109886 10300
rect 110045 10298 110111 10301
rect 109880 10296 110111 10298
rect 109880 10240 110050 10296
rect 110106 10240 110111 10296
rect 109880 10238 110111 10240
rect 109880 10236 109886 10238
rect 109033 10235 109099 10236
rect 110045 10235 110111 10238
rect 110546 10236 110552 10300
rect 110616 10298 110622 10300
rect 110781 10298 110847 10301
rect 110616 10296 110847 10298
rect 110616 10240 110786 10296
rect 110842 10240 110847 10296
rect 110616 10238 110847 10240
rect 110616 10236 110622 10238
rect 110781 10235 110847 10238
rect 111282 10236 111288 10300
rect 111352 10298 111358 10300
rect 111517 10298 111583 10301
rect 111352 10296 111583 10298
rect 111352 10240 111522 10296
rect 111578 10240 111583 10296
rect 111352 10238 111583 10240
rect 111352 10236 111358 10238
rect 111517 10235 111583 10238
rect 112018 10236 112024 10300
rect 112088 10298 112094 10300
rect 112345 10298 112411 10301
rect 112088 10296 112411 10298
rect 112088 10240 112350 10296
rect 112406 10240 112411 10296
rect 112088 10238 112411 10240
rect 112088 10236 112094 10238
rect 112345 10235 112411 10238
rect 112754 10236 112760 10300
rect 112824 10298 112830 10300
rect 112897 10298 112963 10301
rect 113541 10300 113607 10301
rect 113490 10298 113496 10300
rect 112824 10296 112963 10298
rect 112824 10240 112902 10296
rect 112958 10240 112963 10296
rect 112824 10238 112963 10240
rect 113450 10238 113496 10298
rect 113560 10296 113607 10300
rect 113602 10240 113607 10296
rect 112824 10236 112830 10238
rect 112897 10235 112963 10238
rect 113490 10236 113496 10238
rect 113560 10236 113607 10240
rect 113541 10235 113607 10236
rect 114185 10300 114251 10301
rect 114185 10296 114232 10300
rect 114296 10298 114302 10300
rect 114185 10240 114190 10296
rect 114185 10236 114232 10240
rect 114296 10238 114342 10298
rect 114296 10236 114302 10238
rect 114962 10236 114968 10300
rect 115032 10298 115038 10300
rect 115197 10298 115263 10301
rect 115749 10300 115815 10301
rect 115698 10298 115704 10300
rect 115032 10296 115263 10298
rect 115032 10240 115202 10296
rect 115258 10240 115263 10296
rect 115032 10238 115263 10240
rect 115658 10238 115704 10298
rect 115768 10296 115815 10300
rect 115810 10240 115815 10296
rect 115032 10236 115038 10238
rect 114185 10235 114251 10236
rect 115197 10235 115263 10238
rect 115698 10236 115704 10238
rect 115768 10236 115815 10240
rect 116434 10236 116440 10300
rect 116504 10298 116510 10300
rect 116669 10298 116735 10301
rect 117221 10300 117287 10301
rect 117170 10298 117176 10300
rect 116504 10296 116735 10298
rect 116504 10240 116674 10296
rect 116730 10240 116735 10296
rect 116504 10238 116735 10240
rect 117130 10238 117176 10298
rect 117240 10296 117287 10300
rect 117282 10240 117287 10296
rect 116504 10236 116510 10238
rect 115749 10235 115815 10236
rect 116669 10235 116735 10238
rect 117170 10236 117176 10238
rect 117240 10236 117287 10240
rect 117906 10236 117912 10300
rect 117976 10298 117982 10300
rect 118049 10298 118115 10301
rect 118693 10300 118759 10301
rect 117976 10296 118115 10298
rect 117976 10240 118054 10296
rect 118110 10240 118115 10296
rect 117976 10238 118115 10240
rect 117976 10236 117982 10238
rect 117221 10235 117287 10236
rect 118049 10235 118115 10238
rect 118642 10236 118648 10300
rect 118712 10298 118759 10300
rect 119337 10300 119403 10301
rect 118712 10296 118804 10298
rect 118754 10240 118804 10296
rect 118712 10238 118804 10240
rect 119337 10296 119384 10300
rect 119448 10298 119454 10300
rect 119337 10240 119342 10296
rect 118712 10236 118759 10238
rect 118693 10235 118759 10236
rect 119337 10236 119384 10240
rect 119448 10238 119494 10298
rect 119448 10236 119454 10238
rect 120114 10236 120120 10300
rect 120184 10298 120190 10300
rect 120349 10298 120415 10301
rect 120184 10296 120415 10298
rect 120184 10240 120354 10296
rect 120410 10240 120415 10296
rect 120184 10238 120415 10240
rect 120184 10236 120190 10238
rect 119337 10235 119403 10236
rect 120349 10235 120415 10238
rect 120850 10236 120856 10300
rect 120920 10298 120926 10300
rect 121085 10298 121151 10301
rect 120920 10296 121151 10298
rect 120920 10240 121090 10296
rect 121146 10240 121151 10296
rect 120920 10238 121151 10240
rect 120920 10236 120926 10238
rect 121085 10235 121151 10238
rect 121586 10236 121592 10300
rect 121656 10298 121662 10300
rect 121729 10298 121795 10301
rect 122373 10300 122439 10301
rect 121656 10296 121795 10298
rect 121656 10240 121734 10296
rect 121790 10240 121795 10296
rect 121656 10238 121795 10240
rect 121656 10236 121662 10238
rect 121729 10235 121795 10238
rect 122322 10236 122328 10300
rect 122392 10298 122439 10300
rect 122392 10296 122484 10298
rect 122434 10240 122484 10296
rect 122392 10238 122484 10240
rect 122392 10236 122439 10238
rect 123058 10236 123064 10300
rect 123128 10298 123134 10300
rect 123201 10298 123267 10301
rect 123128 10296 123267 10298
rect 123128 10240 123206 10296
rect 123262 10240 123267 10296
rect 123128 10238 123267 10240
rect 123128 10236 123134 10238
rect 122373 10235 122439 10236
rect 123201 10235 123267 10238
rect 123794 10236 123800 10300
rect 123864 10298 123870 10300
rect 124029 10298 124095 10301
rect 123864 10296 124095 10298
rect 123864 10240 124034 10296
rect 124090 10240 124095 10296
rect 123864 10238 124095 10240
rect 123864 10236 123870 10238
rect 124029 10235 124095 10238
rect 124530 10236 124536 10300
rect 124600 10298 124606 10300
rect 125225 10298 125291 10301
rect 124600 10296 125291 10298
rect 124600 10240 125230 10296
rect 125286 10240 125291 10296
rect 124600 10238 125291 10240
rect 124600 10236 124606 10238
rect 125225 10235 125291 10238
rect 126002 10236 126008 10300
rect 126072 10298 126078 10300
rect 126329 10298 126395 10301
rect 126072 10296 126395 10298
rect 126072 10240 126334 10296
rect 126390 10240 126395 10296
rect 126072 10238 126395 10240
rect 126072 10236 126078 10238
rect 126329 10235 126395 10238
rect 126738 10236 126744 10300
rect 126808 10298 126814 10300
rect 126973 10298 127039 10301
rect 126808 10296 127039 10298
rect 126808 10240 126978 10296
rect 127034 10240 127039 10296
rect 126808 10238 127039 10240
rect 126808 10236 126814 10238
rect 126973 10235 127039 10238
rect 127474 10236 127480 10300
rect 127544 10298 127550 10300
rect 127709 10298 127775 10301
rect 128261 10300 128327 10301
rect 128210 10298 128216 10300
rect 127544 10296 127775 10298
rect 127544 10240 127714 10296
rect 127770 10240 127775 10296
rect 127544 10238 127775 10240
rect 128170 10238 128216 10298
rect 128280 10296 128327 10300
rect 128322 10240 128327 10296
rect 127544 10236 127550 10238
rect 127709 10235 127775 10238
rect 128210 10236 128216 10238
rect 128280 10236 128327 10240
rect 128946 10236 128952 10300
rect 129016 10298 129022 10300
rect 129273 10298 129339 10301
rect 129641 10300 129707 10301
rect 129641 10298 129688 10300
rect 129016 10296 129339 10298
rect 129016 10240 129278 10296
rect 129334 10240 129339 10296
rect 129016 10238 129339 10240
rect 129596 10296 129688 10298
rect 129596 10240 129646 10296
rect 129596 10238 129688 10240
rect 129016 10236 129022 10238
rect 128261 10235 128327 10236
rect 129273 10235 129339 10238
rect 129641 10236 129688 10238
rect 129752 10236 129758 10300
rect 130418 10236 130424 10300
rect 130488 10298 130494 10300
rect 130745 10298 130811 10301
rect 130488 10296 130811 10298
rect 130488 10240 130750 10296
rect 130806 10240 130811 10296
rect 130488 10238 130811 10240
rect 130488 10236 130494 10238
rect 129641 10235 129707 10236
rect 130745 10235 130811 10238
rect 131154 10236 131160 10300
rect 131224 10298 131230 10300
rect 131481 10298 131547 10301
rect 131224 10296 131547 10298
rect 131224 10240 131486 10296
rect 131542 10240 131547 10296
rect 131224 10238 131547 10240
rect 131224 10236 131230 10238
rect 131481 10235 131547 10238
rect 131890 10236 131896 10300
rect 131960 10298 131966 10300
rect 132125 10298 132191 10301
rect 131960 10296 132191 10298
rect 131960 10240 132130 10296
rect 132186 10240 132191 10296
rect 131960 10238 132191 10240
rect 131960 10236 131966 10238
rect 132125 10235 132191 10238
rect 132626 10236 132632 10300
rect 132696 10298 132702 10300
rect 132953 10298 133019 10301
rect 133413 10300 133479 10301
rect 134149 10300 134215 10301
rect 132696 10296 133019 10298
rect 132696 10240 132958 10296
rect 133014 10240 133019 10296
rect 132696 10238 133019 10240
rect 132696 10236 132702 10238
rect 132953 10235 133019 10238
rect 133362 10236 133368 10300
rect 133432 10298 133479 10300
rect 133432 10296 133524 10298
rect 133474 10240 133524 10296
rect 133432 10238 133524 10240
rect 133432 10236 133479 10238
rect 134098 10236 134104 10300
rect 134168 10298 134215 10300
rect 134701 10298 134767 10301
rect 134834 10298 134840 10300
rect 134168 10296 134260 10298
rect 134210 10240 134260 10296
rect 134168 10238 134260 10240
rect 134701 10296 134840 10298
rect 134701 10240 134706 10296
rect 134762 10240 134840 10296
rect 134701 10238 134840 10240
rect 134168 10236 134215 10238
rect 133413 10235 133479 10236
rect 134149 10235 134215 10236
rect 134701 10235 134767 10238
rect 134834 10236 134840 10238
rect 134904 10236 134910 10300
rect 138054 10236 138060 10300
rect 138124 10298 138130 10300
rect 138749 10298 138815 10301
rect 138124 10296 138815 10298
rect 138124 10240 138754 10296
rect 138810 10240 138815 10296
rect 138124 10238 138815 10240
rect 138124 10236 138130 10238
rect 138749 10235 138815 10238
rect 142470 10236 142476 10300
rect 142540 10298 142546 10300
rect 143257 10298 143323 10301
rect 142540 10296 143323 10298
rect 142540 10240 143262 10296
rect 143318 10240 143323 10296
rect 142540 10238 143323 10240
rect 142540 10236 142546 10238
rect 143257 10235 143323 10238
rect 148358 10236 148364 10300
rect 148428 10298 148434 10300
rect 149053 10298 149119 10301
rect 148428 10296 149119 10298
rect 148428 10240 149058 10296
rect 149114 10240 149119 10296
rect 148428 10238 149119 10240
rect 148428 10236 148434 10238
rect 149053 10235 149119 10238
rect 171450 10236 171456 10300
rect 171520 10298 171526 10300
rect 171685 10298 171751 10301
rect 171520 10296 171751 10298
rect 171520 10240 171690 10296
rect 171746 10240 171751 10296
rect 171520 10238 171751 10240
rect 171520 10236 171526 10238
rect 171685 10235 171751 10238
rect 173658 10236 173664 10300
rect 173728 10298 173734 10300
rect 173893 10298 173959 10301
rect 174445 10300 174511 10301
rect 175181 10300 175247 10301
rect 175917 10300 175983 10301
rect 174394 10298 174400 10300
rect 173728 10296 173959 10298
rect 173728 10240 173898 10296
rect 173954 10240 173959 10296
rect 173728 10238 173959 10240
rect 174354 10238 174400 10298
rect 174464 10296 174511 10300
rect 175130 10298 175136 10300
rect 174506 10240 174511 10296
rect 173728 10236 173734 10238
rect 173893 10235 173959 10238
rect 174394 10236 174400 10238
rect 174464 10236 174511 10240
rect 175090 10238 175136 10298
rect 175200 10296 175247 10300
rect 175866 10298 175872 10300
rect 175242 10240 175247 10296
rect 175130 10236 175136 10238
rect 175200 10236 175247 10240
rect 175826 10238 175872 10298
rect 175936 10296 175983 10300
rect 175978 10240 175983 10296
rect 175866 10236 175872 10238
rect 175936 10236 175983 10240
rect 176602 10236 176608 10300
rect 176672 10298 176678 10300
rect 176745 10298 176811 10301
rect 176672 10296 176811 10298
rect 176672 10240 176750 10296
rect 176806 10240 176811 10296
rect 176672 10238 176811 10240
rect 176672 10236 176678 10238
rect 174445 10235 174511 10236
rect 175181 10235 175247 10236
rect 175917 10235 175983 10236
rect 176745 10235 176811 10238
rect 177338 10236 177344 10300
rect 177408 10298 177414 10300
rect 177481 10298 177547 10301
rect 177408 10296 177547 10298
rect 177408 10240 177486 10296
rect 177542 10240 177547 10296
rect 177408 10238 177547 10240
rect 177408 10236 177414 10238
rect 177481 10235 177547 10238
rect 177941 10298 178007 10301
rect 178074 10298 178080 10300
rect 177941 10296 178080 10298
rect 177941 10240 177946 10296
rect 178002 10240 178080 10296
rect 177941 10238 178080 10240
rect 177941 10235 178007 10238
rect 178074 10236 178080 10238
rect 178144 10236 178150 10300
rect 178810 10236 178816 10300
rect 178880 10298 178886 10300
rect 179137 10298 179203 10301
rect 178880 10296 179203 10298
rect 178880 10240 179142 10296
rect 179198 10240 179203 10296
rect 178880 10238 179203 10240
rect 178880 10236 178886 10238
rect 179137 10235 179203 10238
rect 180282 10236 180288 10300
rect 180352 10298 180358 10300
rect 180425 10298 180491 10301
rect 180352 10296 180491 10298
rect 180352 10240 180430 10296
rect 180486 10240 180491 10296
rect 180352 10238 180491 10240
rect 180352 10236 180358 10238
rect 180425 10235 180491 10238
rect 181754 10236 181760 10300
rect 181824 10298 181830 10300
rect 181897 10298 181963 10301
rect 182541 10300 182607 10301
rect 183277 10300 183343 10301
rect 182490 10298 182496 10300
rect 181824 10296 181963 10298
rect 181824 10240 181902 10296
rect 181958 10240 181963 10296
rect 181824 10238 181963 10240
rect 182450 10238 182496 10298
rect 182560 10296 182607 10300
rect 183226 10298 183232 10300
rect 182602 10240 182607 10296
rect 181824 10236 181830 10238
rect 181897 10235 181963 10238
rect 182490 10236 182496 10238
rect 182560 10236 182607 10240
rect 183186 10238 183232 10298
rect 183296 10296 183343 10300
rect 183338 10240 183343 10296
rect 183226 10236 183232 10238
rect 183296 10236 183343 10240
rect 183962 10236 183968 10300
rect 184032 10298 184038 10300
rect 184289 10298 184355 10301
rect 184749 10300 184815 10301
rect 185485 10300 185551 10301
rect 186221 10300 186287 10301
rect 186957 10300 187023 10301
rect 187693 10300 187759 10301
rect 184698 10298 184704 10300
rect 184032 10296 184355 10298
rect 184032 10240 184294 10296
rect 184350 10240 184355 10296
rect 184032 10238 184355 10240
rect 184658 10238 184704 10298
rect 184768 10296 184815 10300
rect 185434 10298 185440 10300
rect 184810 10240 184815 10296
rect 184032 10236 184038 10238
rect 182541 10235 182607 10236
rect 183277 10235 183343 10236
rect 184289 10235 184355 10238
rect 184698 10236 184704 10238
rect 184768 10236 184815 10240
rect 185394 10238 185440 10298
rect 185504 10296 185551 10300
rect 186170 10298 186176 10300
rect 185546 10240 185551 10296
rect 185434 10236 185440 10238
rect 185504 10236 185551 10240
rect 186130 10238 186176 10298
rect 186240 10296 186287 10300
rect 186906 10298 186912 10300
rect 186282 10240 186287 10296
rect 186170 10236 186176 10238
rect 186240 10236 186287 10240
rect 186866 10238 186912 10298
rect 186976 10296 187023 10300
rect 187642 10298 187648 10300
rect 187018 10240 187023 10296
rect 186906 10236 186912 10238
rect 186976 10236 187023 10240
rect 187602 10238 187648 10298
rect 187712 10296 187759 10300
rect 187754 10240 187759 10296
rect 187642 10236 187648 10238
rect 187712 10236 187759 10240
rect 188378 10236 188384 10300
rect 188448 10298 188454 10300
rect 188613 10298 188679 10301
rect 188448 10296 188679 10298
rect 188448 10240 188618 10296
rect 188674 10240 188679 10296
rect 188448 10238 188679 10240
rect 188448 10236 188454 10238
rect 184749 10235 184815 10236
rect 185485 10235 185551 10236
rect 186221 10235 186287 10236
rect 186957 10235 187023 10236
rect 187693 10235 187759 10236
rect 188613 10235 188679 10238
rect 189114 10236 189120 10300
rect 189184 10298 189190 10300
rect 189441 10298 189507 10301
rect 189901 10300 189967 10301
rect 191373 10300 191439 10301
rect 189850 10298 189856 10300
rect 189184 10296 189507 10298
rect 189184 10240 189446 10296
rect 189502 10240 189507 10296
rect 189184 10238 189507 10240
rect 189810 10238 189856 10298
rect 189920 10296 189967 10300
rect 189962 10240 189967 10296
rect 189184 10236 189190 10238
rect 189441 10235 189507 10238
rect 189850 10236 189856 10238
rect 189920 10236 189967 10240
rect 191322 10236 191328 10300
rect 191392 10298 191439 10300
rect 191392 10296 191484 10298
rect 191434 10240 191484 10296
rect 191392 10238 191484 10240
rect 191392 10236 191439 10238
rect 192058 10236 192064 10300
rect 192128 10298 192134 10300
rect 192937 10298 193003 10301
rect 192128 10296 193003 10298
rect 192128 10240 192942 10296
rect 192998 10240 193003 10296
rect 192128 10238 193003 10240
rect 192128 10236 192134 10238
rect 189901 10235 189967 10236
rect 191373 10235 191439 10236
rect 192937 10235 193003 10238
rect 193530 10236 193536 10300
rect 193600 10298 193606 10300
rect 194041 10298 194107 10301
rect 194317 10300 194383 10301
rect 193600 10296 194107 10298
rect 193600 10240 194046 10296
rect 194102 10240 194107 10296
rect 193600 10238 194107 10240
rect 193600 10236 193606 10238
rect 194041 10235 194107 10238
rect 194266 10236 194272 10300
rect 194336 10298 194383 10300
rect 194336 10296 194428 10298
rect 194378 10240 194428 10296
rect 194336 10238 194428 10240
rect 194336 10236 194383 10238
rect 195002 10236 195008 10300
rect 195072 10298 195078 10300
rect 195513 10298 195579 10301
rect 195789 10300 195855 10301
rect 196525 10300 196591 10301
rect 197261 10300 197327 10301
rect 197997 10300 198063 10301
rect 195072 10296 195579 10298
rect 195072 10240 195518 10296
rect 195574 10240 195579 10296
rect 195072 10238 195579 10240
rect 195072 10236 195078 10238
rect 194317 10235 194383 10236
rect 195513 10235 195579 10238
rect 195738 10236 195744 10300
rect 195808 10298 195855 10300
rect 195808 10296 195900 10298
rect 195850 10240 195900 10296
rect 195808 10238 195900 10240
rect 195808 10236 195855 10238
rect 196474 10236 196480 10300
rect 196544 10298 196591 10300
rect 196544 10296 196636 10298
rect 196586 10240 196636 10296
rect 196544 10238 196636 10240
rect 196544 10236 196591 10238
rect 197210 10236 197216 10300
rect 197280 10298 197327 10300
rect 197280 10296 197372 10298
rect 197322 10240 197372 10296
rect 197280 10238 197372 10240
rect 197280 10236 197327 10238
rect 197946 10236 197952 10300
rect 198016 10298 198063 10300
rect 198016 10296 198108 10298
rect 198058 10240 198108 10296
rect 198016 10238 198108 10240
rect 198016 10236 198063 10238
rect 198682 10236 198688 10300
rect 198752 10298 198758 10300
rect 199101 10298 199167 10301
rect 198752 10296 199167 10298
rect 198752 10240 199106 10296
rect 199162 10240 199167 10296
rect 198752 10238 199167 10240
rect 198752 10236 198758 10238
rect 195789 10235 195855 10236
rect 196525 10235 196591 10236
rect 197261 10235 197327 10236
rect 197997 10235 198063 10236
rect 199101 10235 199167 10238
rect 199418 10236 199424 10300
rect 199488 10298 199494 10300
rect 199929 10298 199995 10301
rect 199488 10296 199995 10298
rect 199488 10240 199934 10296
rect 199990 10240 199995 10296
rect 199488 10238 199995 10240
rect 199488 10236 199494 10238
rect 199929 10235 199995 10238
rect 200154 10236 200160 10300
rect 200224 10298 200230 10300
rect 200757 10298 200823 10301
rect 200941 10300 201007 10301
rect 200224 10296 200823 10298
rect 200224 10240 200762 10296
rect 200818 10240 200823 10296
rect 200224 10238 200823 10240
rect 200224 10236 200230 10238
rect 200757 10235 200823 10238
rect 200890 10236 200896 10300
rect 200960 10298 201007 10300
rect 200960 10296 201052 10298
rect 201002 10240 201052 10296
rect 200960 10238 201052 10240
rect 200960 10236 201007 10238
rect 201626 10236 201632 10300
rect 201696 10298 201702 10300
rect 202505 10298 202571 10301
rect 201696 10296 202571 10298
rect 201696 10240 202510 10296
rect 202566 10240 202571 10296
rect 201696 10238 202571 10240
rect 201696 10236 201702 10238
rect 200941 10235 201007 10236
rect 202505 10235 202571 10238
rect 203098 10236 203104 10300
rect 203168 10298 203174 10300
rect 204069 10298 204135 10301
rect 203168 10296 204135 10298
rect 203168 10240 204074 10296
rect 204130 10240 204135 10296
rect 203168 10238 204135 10240
rect 203168 10236 203174 10238
rect 204069 10235 204135 10238
rect 205582 10236 205588 10300
rect 205652 10298 205658 10300
rect 205817 10298 205883 10301
rect 220353 10300 220419 10301
rect 220302 10298 220308 10300
rect 205652 10296 205883 10298
rect 205652 10240 205822 10296
rect 205878 10240 205883 10296
rect 205652 10238 205883 10240
rect 220262 10238 220308 10298
rect 220372 10296 220419 10300
rect 220414 10240 220419 10296
rect 205652 10236 205658 10238
rect 205817 10235 205883 10238
rect 220302 10236 220308 10238
rect 220372 10236 220419 10240
rect 239714 10236 239720 10300
rect 239784 10298 239790 10300
rect 239949 10298 240015 10301
rect 239784 10296 240015 10298
rect 239784 10240 239954 10296
rect 240010 10240 240015 10296
rect 239784 10238 240015 10240
rect 239784 10236 239790 10238
rect 220353 10235 220419 10236
rect 239949 10235 240015 10238
rect 240450 10236 240456 10300
rect 240520 10298 240526 10300
rect 240961 10298 241027 10301
rect 241237 10300 241303 10301
rect 241186 10298 241192 10300
rect 240520 10296 241027 10298
rect 240520 10240 240966 10296
rect 241022 10240 241027 10296
rect 240520 10238 241027 10240
rect 241146 10238 241192 10298
rect 241256 10296 241303 10300
rect 241298 10240 241303 10296
rect 240520 10236 240526 10238
rect 240961 10235 241027 10238
rect 241186 10236 241192 10238
rect 241256 10236 241303 10240
rect 241922 10236 241928 10300
rect 241992 10298 241998 10300
rect 242341 10298 242407 10301
rect 241992 10296 242407 10298
rect 241992 10240 242346 10296
rect 242402 10240 242407 10296
rect 241992 10238 242407 10240
rect 241992 10236 241998 10238
rect 241237 10235 241303 10236
rect 242341 10235 242407 10238
rect 242658 10236 242664 10300
rect 242728 10298 242734 10300
rect 242893 10298 242959 10301
rect 243445 10300 243511 10301
rect 244181 10300 244247 10301
rect 243394 10298 243400 10300
rect 242728 10296 242959 10298
rect 242728 10240 242898 10296
rect 242954 10240 242959 10296
rect 242728 10238 242959 10240
rect 243354 10238 243400 10298
rect 243464 10296 243511 10300
rect 244130 10298 244136 10300
rect 243506 10240 243511 10296
rect 242728 10236 242734 10238
rect 242893 10235 242959 10238
rect 243394 10236 243400 10238
rect 243464 10236 243511 10240
rect 244090 10238 244136 10298
rect 244200 10296 244247 10300
rect 244242 10240 244247 10296
rect 244130 10236 244136 10238
rect 244200 10236 244247 10240
rect 244866 10236 244872 10300
rect 244936 10298 244942 10300
rect 245009 10298 245075 10301
rect 246389 10300 246455 10301
rect 247125 10300 247191 10301
rect 246338 10298 246344 10300
rect 244936 10296 245075 10298
rect 244936 10240 245014 10296
rect 245070 10240 245075 10296
rect 244936 10238 245075 10240
rect 246298 10238 246344 10298
rect 246408 10296 246455 10300
rect 247074 10298 247080 10300
rect 246450 10240 246455 10296
rect 244936 10236 244942 10238
rect 243445 10235 243511 10236
rect 244181 10235 244247 10236
rect 245009 10235 245075 10238
rect 246338 10236 246344 10238
rect 246408 10236 246455 10240
rect 247034 10238 247080 10298
rect 247144 10296 247191 10300
rect 247186 10240 247191 10296
rect 247074 10236 247080 10238
rect 247144 10236 247191 10240
rect 247810 10236 247816 10300
rect 247880 10298 247886 10300
rect 247953 10298 248019 10301
rect 247880 10296 248019 10298
rect 247880 10240 247958 10296
rect 248014 10240 248019 10296
rect 247880 10238 248019 10240
rect 247880 10236 247886 10238
rect 246389 10235 246455 10236
rect 247125 10235 247191 10236
rect 247953 10235 248019 10238
rect 248546 10236 248552 10300
rect 248616 10298 248622 10300
rect 248689 10298 248755 10301
rect 249333 10300 249399 10301
rect 249282 10298 249288 10300
rect 248616 10296 248755 10298
rect 248616 10240 248694 10296
rect 248750 10240 248755 10296
rect 248616 10238 248755 10240
rect 249242 10238 249288 10298
rect 249352 10296 249399 10300
rect 249394 10240 249399 10296
rect 248616 10236 248622 10238
rect 248689 10235 248755 10238
rect 249282 10236 249288 10238
rect 249352 10236 249399 10240
rect 250018 10236 250024 10300
rect 250088 10298 250094 10300
rect 250161 10298 250227 10301
rect 250088 10296 250227 10298
rect 250088 10240 250166 10296
rect 250222 10240 250227 10296
rect 250088 10238 250227 10240
rect 250088 10236 250094 10238
rect 249333 10235 249399 10236
rect 250161 10235 250227 10238
rect 250754 10236 250760 10300
rect 250824 10298 250830 10300
rect 251173 10298 251239 10301
rect 251541 10300 251607 10301
rect 252277 10300 252343 10301
rect 253749 10300 253815 10301
rect 251490 10298 251496 10300
rect 250824 10296 251239 10298
rect 250824 10240 251178 10296
rect 251234 10240 251239 10296
rect 250824 10238 251239 10240
rect 251450 10238 251496 10298
rect 251560 10296 251607 10300
rect 252226 10298 252232 10300
rect 251602 10240 251607 10296
rect 250824 10236 250830 10238
rect 251173 10235 251239 10238
rect 251490 10236 251496 10238
rect 251560 10236 251607 10240
rect 252186 10238 252232 10298
rect 252296 10296 252343 10300
rect 253698 10298 253704 10300
rect 252338 10240 252343 10296
rect 252226 10236 252232 10238
rect 252296 10236 252343 10240
rect 253658 10238 253704 10298
rect 253768 10296 253815 10300
rect 253810 10240 253815 10296
rect 253698 10236 253704 10238
rect 253768 10236 253815 10240
rect 254434 10236 254440 10300
rect 254504 10298 254510 10300
rect 255037 10298 255103 10301
rect 254504 10296 255103 10298
rect 254504 10240 255042 10296
rect 255098 10240 255103 10296
rect 254504 10238 255103 10240
rect 254504 10236 254510 10238
rect 251541 10235 251607 10236
rect 252277 10235 252343 10236
rect 253749 10235 253815 10236
rect 255037 10235 255103 10238
rect 255170 10236 255176 10300
rect 255240 10298 255246 10300
rect 255313 10298 255379 10301
rect 255240 10296 255379 10298
rect 255240 10240 255318 10296
rect 255374 10240 255379 10296
rect 255240 10238 255379 10240
rect 255240 10236 255246 10238
rect 255313 10235 255379 10238
rect 255906 10236 255912 10300
rect 255976 10298 255982 10300
rect 256417 10298 256483 10301
rect 256693 10300 256759 10301
rect 256642 10298 256648 10300
rect 255976 10296 256483 10298
rect 255976 10240 256422 10296
rect 256478 10240 256483 10296
rect 255976 10238 256483 10240
rect 256602 10238 256648 10298
rect 256712 10296 256759 10300
rect 256754 10240 256759 10296
rect 255976 10236 255982 10238
rect 256417 10235 256483 10238
rect 256642 10236 256648 10238
rect 256712 10236 256759 10240
rect 257378 10236 257384 10300
rect 257448 10298 257454 10300
rect 257705 10298 257771 10301
rect 257448 10296 257771 10298
rect 257448 10240 257710 10296
rect 257766 10240 257771 10296
rect 257448 10238 257771 10240
rect 257448 10236 257454 10238
rect 256693 10235 256759 10236
rect 257705 10235 257771 10238
rect 258114 10236 258120 10300
rect 258184 10298 258190 10300
rect 258257 10298 258323 10301
rect 258184 10296 258323 10298
rect 258184 10240 258262 10296
rect 258318 10240 258323 10296
rect 258184 10238 258323 10240
rect 258184 10236 258190 10238
rect 258257 10235 258323 10238
rect 258850 10236 258856 10300
rect 258920 10298 258926 10300
rect 259177 10298 259243 10301
rect 258920 10296 259243 10298
rect 258920 10240 259182 10296
rect 259238 10240 259243 10296
rect 258920 10238 259243 10240
rect 258920 10236 258926 10238
rect 259177 10235 259243 10238
rect 259586 10236 259592 10300
rect 259656 10298 259662 10300
rect 259913 10298 259979 10301
rect 259656 10296 259979 10298
rect 259656 10240 259918 10296
rect 259974 10240 259979 10296
rect 259656 10238 259979 10240
rect 259656 10236 259662 10238
rect 259913 10235 259979 10238
rect 260322 10236 260328 10300
rect 260392 10298 260398 10300
rect 260465 10298 260531 10301
rect 261845 10300 261911 10301
rect 260392 10296 260531 10298
rect 260392 10240 260470 10296
rect 260526 10240 260531 10296
rect 260392 10238 260531 10240
rect 260392 10236 260398 10238
rect 260465 10235 260531 10238
rect 261794 10236 261800 10300
rect 261864 10298 261911 10300
rect 262489 10300 262555 10301
rect 263317 10300 263383 10301
rect 262489 10298 262536 10300
rect 261864 10296 261956 10298
rect 261906 10240 261956 10296
rect 261864 10238 261956 10240
rect 262444 10296 262536 10298
rect 262444 10240 262494 10296
rect 262444 10238 262536 10240
rect 261864 10236 261911 10238
rect 261845 10235 261911 10236
rect 262489 10236 262536 10238
rect 262600 10236 262606 10300
rect 263266 10236 263272 10300
rect 263336 10298 263383 10300
rect 263336 10296 263428 10298
rect 263378 10240 263428 10296
rect 263336 10238 263428 10240
rect 263336 10236 263383 10238
rect 264002 10236 264008 10300
rect 264072 10298 264078 10300
rect 264329 10298 264395 10301
rect 266169 10300 266235 10301
rect 266169 10298 266216 10300
rect 264072 10296 264395 10298
rect 264072 10240 264334 10296
rect 264390 10240 264395 10296
rect 264072 10238 264395 10240
rect 266124 10296 266216 10298
rect 266124 10240 266174 10296
rect 266124 10238 266216 10240
rect 264072 10236 264078 10238
rect 262489 10235 262555 10236
rect 263317 10235 263383 10236
rect 264329 10235 264395 10238
rect 266169 10236 266216 10238
rect 266280 10236 266286 10300
rect 266169 10235 266235 10236
rect 1526 10100 1532 10164
rect 1596 10162 1602 10164
rect 1669 10162 1735 10165
rect 1596 10160 1735 10162
rect 1596 10104 1674 10160
rect 1730 10104 1735 10160
rect 1596 10102 1735 10104
rect 1596 10100 1602 10102
rect 1669 10099 1735 10102
rect 2262 10100 2268 10164
rect 2332 10162 2338 10164
rect 2405 10162 2471 10165
rect 2332 10160 2471 10162
rect 2332 10104 2410 10160
rect 2466 10104 2471 10160
rect 2332 10102 2471 10104
rect 2332 10100 2338 10102
rect 2405 10099 2471 10102
rect 3233 10162 3299 10165
rect 3734 10162 3740 10164
rect 3233 10160 3740 10162
rect 3233 10104 3238 10160
rect 3294 10104 3740 10160
rect 3233 10102 3740 10104
rect 3233 10099 3299 10102
rect 3734 10100 3740 10102
rect 3804 10100 3810 10164
rect 4337 10162 4403 10165
rect 4470 10162 4476 10164
rect 4337 10160 4476 10162
rect 4337 10104 4342 10160
rect 4398 10104 4476 10160
rect 4337 10102 4476 10104
rect 4337 10099 4403 10102
rect 4470 10100 4476 10102
rect 4540 10100 4546 10164
rect 5073 10162 5139 10165
rect 5206 10162 5212 10164
rect 5073 10160 5212 10162
rect 5073 10104 5078 10160
rect 5134 10104 5212 10160
rect 5073 10102 5212 10104
rect 5073 10099 5139 10102
rect 5206 10100 5212 10102
rect 5276 10100 5282 10164
rect 5809 10162 5875 10165
rect 5942 10162 5948 10164
rect 5809 10160 5948 10162
rect 5809 10104 5814 10160
rect 5870 10104 5948 10160
rect 5809 10102 5948 10104
rect 5809 10099 5875 10102
rect 5942 10100 5948 10102
rect 6012 10100 6018 10164
rect 6678 10100 6684 10164
rect 6748 10162 6754 10164
rect 6821 10162 6887 10165
rect 6748 10160 6887 10162
rect 6748 10104 6826 10160
rect 6882 10104 6887 10160
rect 6748 10102 6887 10104
rect 6748 10100 6754 10102
rect 6821 10099 6887 10102
rect 7414 10100 7420 10164
rect 7484 10162 7490 10164
rect 7557 10162 7623 10165
rect 7484 10160 7623 10162
rect 7484 10104 7562 10160
rect 7618 10104 7623 10160
rect 7484 10102 7623 10104
rect 7484 10100 7490 10102
rect 7557 10099 7623 10102
rect 8385 10162 8451 10165
rect 9581 10164 9647 10165
rect 8886 10162 8892 10164
rect 8385 10160 8892 10162
rect 8385 10104 8390 10160
rect 8446 10104 8892 10160
rect 8385 10102 8892 10104
rect 8385 10099 8451 10102
rect 8886 10100 8892 10102
rect 8956 10100 8962 10164
rect 9581 10160 9628 10164
rect 9692 10162 9698 10164
rect 10225 10162 10291 10165
rect 10358 10162 10364 10164
rect 9581 10104 9586 10160
rect 9581 10100 9628 10104
rect 9692 10102 9738 10162
rect 10225 10160 10364 10162
rect 10225 10104 10230 10160
rect 10286 10104 10364 10160
rect 10225 10102 10364 10104
rect 9692 10100 9698 10102
rect 9581 10099 9647 10100
rect 10225 10099 10291 10102
rect 10358 10100 10364 10102
rect 10428 10100 10434 10164
rect 10961 10162 11027 10165
rect 11094 10162 11100 10164
rect 10961 10160 11100 10162
rect 10961 10104 10966 10160
rect 11022 10104 11100 10160
rect 10961 10102 11100 10104
rect 10961 10099 11027 10102
rect 11094 10100 11100 10102
rect 11164 10100 11170 10164
rect 11830 10100 11836 10164
rect 11900 10162 11906 10164
rect 11973 10162 12039 10165
rect 11900 10160 12039 10162
rect 11900 10104 11978 10160
rect 12034 10104 12039 10160
rect 11900 10102 12039 10104
rect 11900 10100 11906 10102
rect 11973 10099 12039 10102
rect 12566 10100 12572 10164
rect 12636 10162 12642 10164
rect 12709 10162 12775 10165
rect 12636 10160 12775 10162
rect 12636 10104 12714 10160
rect 12770 10104 12775 10160
rect 12636 10102 12775 10104
rect 12636 10100 12642 10102
rect 12709 10099 12775 10102
rect 13721 10162 13787 10165
rect 14038 10162 14044 10164
rect 13721 10160 14044 10162
rect 13721 10104 13726 10160
rect 13782 10104 14044 10160
rect 13721 10102 14044 10104
rect 13721 10099 13787 10102
rect 14038 10100 14044 10102
rect 14108 10100 14114 10164
rect 14641 10162 14707 10165
rect 14774 10162 14780 10164
rect 14641 10160 14780 10162
rect 14641 10104 14646 10160
rect 14702 10104 14780 10160
rect 14641 10102 14780 10104
rect 14641 10099 14707 10102
rect 14774 10100 14780 10102
rect 14844 10100 14850 10164
rect 15377 10162 15443 10165
rect 15510 10162 15516 10164
rect 15377 10160 15516 10162
rect 15377 10104 15382 10160
rect 15438 10104 15516 10160
rect 15377 10102 15516 10104
rect 15377 10099 15443 10102
rect 15510 10100 15516 10102
rect 15580 10100 15586 10164
rect 16113 10162 16179 10165
rect 16246 10162 16252 10164
rect 16113 10160 16252 10162
rect 16113 10104 16118 10160
rect 16174 10104 16252 10160
rect 16113 10102 16252 10104
rect 16113 10099 16179 10102
rect 16246 10100 16252 10102
rect 16316 10100 16322 10164
rect 16982 10100 16988 10164
rect 17052 10162 17058 10164
rect 17125 10162 17191 10165
rect 17052 10160 17191 10162
rect 17052 10104 17130 10160
rect 17186 10104 17191 10160
rect 17052 10102 17191 10104
rect 17052 10100 17058 10102
rect 17125 10099 17191 10102
rect 17718 10100 17724 10164
rect 17788 10162 17794 10164
rect 17861 10162 17927 10165
rect 17788 10160 17927 10162
rect 17788 10104 17866 10160
rect 17922 10104 17927 10160
rect 17788 10102 17927 10104
rect 17788 10100 17794 10102
rect 17861 10099 17927 10102
rect 18454 10100 18460 10164
rect 18524 10162 18530 10164
rect 18597 10162 18663 10165
rect 18524 10160 18663 10162
rect 18524 10104 18602 10160
rect 18658 10104 18663 10160
rect 18524 10102 18663 10104
rect 18524 10100 18530 10102
rect 18597 10099 18663 10102
rect 71262 10100 71268 10164
rect 71332 10162 71338 10164
rect 71497 10162 71563 10165
rect 71332 10160 71563 10162
rect 71332 10104 71502 10160
rect 71558 10104 71563 10160
rect 71332 10102 71563 10104
rect 71332 10100 71338 10102
rect 71497 10099 71563 10102
rect 79225 10162 79291 10165
rect 83089 10164 83155 10165
rect 79358 10162 79364 10164
rect 79225 10160 79364 10162
rect 79225 10104 79230 10160
rect 79286 10104 79364 10160
rect 79225 10102 79364 10104
rect 79225 10099 79291 10102
rect 79358 10100 79364 10102
rect 79428 10100 79434 10164
rect 83038 10162 83044 10164
rect 82998 10102 83044 10162
rect 83108 10160 83155 10164
rect 83150 10104 83155 10160
rect 83038 10100 83044 10102
rect 83108 10100 83155 10104
rect 83774 10100 83780 10164
rect 83844 10162 83850 10164
rect 83917 10162 83983 10165
rect 83844 10160 83983 10162
rect 83844 10104 83922 10160
rect 83978 10104 83983 10160
rect 83844 10102 83983 10104
rect 83844 10100 83850 10102
rect 83089 10099 83155 10100
rect 83917 10099 83983 10102
rect 84510 10100 84516 10164
rect 84580 10162 84586 10164
rect 84653 10162 84719 10165
rect 84580 10160 84719 10162
rect 84580 10104 84658 10160
rect 84714 10104 84719 10160
rect 84580 10102 84719 10104
rect 84580 10100 84586 10102
rect 84653 10099 84719 10102
rect 85246 10100 85252 10164
rect 85316 10162 85322 10164
rect 85389 10162 85455 10165
rect 85316 10160 85455 10162
rect 85316 10104 85394 10160
rect 85450 10104 85455 10160
rect 85316 10102 85455 10104
rect 85316 10100 85322 10102
rect 85389 10099 85455 10102
rect 138790 10100 138796 10164
rect 138860 10162 138866 10164
rect 139393 10162 139459 10165
rect 138860 10160 139459 10162
rect 138860 10104 139398 10160
rect 139454 10104 139459 10160
rect 138860 10102 139459 10104
rect 138860 10100 138866 10102
rect 139393 10099 139459 10102
rect 140262 10100 140268 10164
rect 140332 10162 140338 10164
rect 140681 10162 140747 10165
rect 140332 10160 140747 10162
rect 140332 10104 140686 10160
rect 140742 10104 140747 10160
rect 140332 10102 140747 10104
rect 140332 10100 140338 10102
rect 140681 10099 140747 10102
rect 140998 10100 141004 10164
rect 141068 10162 141074 10164
rect 141325 10162 141391 10165
rect 141068 10160 141391 10162
rect 141068 10104 141330 10160
rect 141386 10104 141391 10160
rect 141068 10102 141391 10104
rect 141068 10100 141074 10102
rect 141325 10099 141391 10102
rect 141734 10100 141740 10164
rect 141804 10162 141810 10164
rect 141969 10162 142035 10165
rect 141804 10160 142035 10162
rect 141804 10104 141974 10160
rect 142030 10104 142035 10160
rect 141804 10102 142035 10104
rect 141804 10100 141810 10102
rect 141969 10099 142035 10102
rect 143206 10100 143212 10164
rect 143276 10162 143282 10164
rect 143533 10162 143599 10165
rect 143276 10160 143599 10162
rect 143276 10104 143538 10160
rect 143594 10104 143599 10160
rect 143276 10102 143599 10104
rect 143276 10100 143282 10102
rect 143533 10099 143599 10102
rect 143942 10100 143948 10164
rect 144012 10162 144018 10164
rect 144545 10162 144611 10165
rect 144012 10160 144611 10162
rect 144012 10104 144550 10160
rect 144606 10104 144611 10160
rect 144012 10102 144611 10104
rect 144012 10100 144018 10102
rect 144545 10099 144611 10102
rect 145414 10100 145420 10164
rect 145484 10162 145490 10164
rect 145833 10162 145899 10165
rect 145484 10160 145899 10162
rect 145484 10104 145838 10160
rect 145894 10104 145899 10160
rect 145484 10102 145899 10104
rect 145484 10100 145490 10102
rect 145833 10099 145899 10102
rect 146150 10100 146156 10164
rect 146220 10162 146226 10164
rect 146293 10162 146359 10165
rect 146220 10160 146359 10162
rect 146220 10104 146298 10160
rect 146354 10104 146359 10160
rect 146220 10102 146359 10104
rect 146220 10100 146226 10102
rect 146293 10099 146359 10102
rect 146886 10100 146892 10164
rect 146956 10162 146962 10164
rect 147121 10162 147187 10165
rect 146956 10160 147187 10162
rect 146956 10104 147126 10160
rect 147182 10104 147187 10160
rect 146956 10102 147187 10104
rect 146956 10100 146962 10102
rect 147121 10099 147187 10102
rect 149094 10100 149100 10164
rect 149164 10162 149170 10164
rect 149697 10162 149763 10165
rect 149164 10160 149763 10162
rect 149164 10104 149702 10160
rect 149758 10104 149763 10160
rect 149164 10102 149763 10104
rect 149164 10100 149170 10102
rect 149697 10099 149763 10102
rect 150566 10100 150572 10164
rect 150636 10162 150642 10164
rect 150985 10162 151051 10165
rect 150636 10160 151051 10162
rect 150636 10104 150990 10160
rect 151046 10104 151051 10160
rect 150636 10102 151051 10104
rect 150636 10100 150642 10102
rect 150985 10099 151051 10102
rect 151302 10100 151308 10164
rect 151372 10162 151378 10164
rect 151629 10162 151695 10165
rect 151372 10160 151695 10162
rect 151372 10104 151634 10160
rect 151690 10104 151695 10160
rect 151372 10102 151695 10104
rect 151372 10100 151378 10102
rect 151629 10099 151695 10102
rect 152038 10100 152044 10164
rect 152108 10162 152114 10164
rect 152273 10162 152339 10165
rect 152825 10164 152891 10165
rect 152774 10162 152780 10164
rect 152108 10160 152339 10162
rect 152108 10104 152278 10160
rect 152334 10104 152339 10160
rect 152108 10102 152339 10104
rect 152734 10102 152780 10162
rect 152844 10160 152891 10164
rect 152886 10104 152891 10160
rect 152108 10100 152114 10102
rect 152273 10099 152339 10102
rect 152774 10100 152780 10102
rect 152844 10100 152891 10104
rect 153510 10100 153516 10164
rect 153580 10162 153586 10164
rect 154205 10162 154271 10165
rect 153580 10160 154271 10162
rect 153580 10104 154210 10160
rect 154266 10104 154271 10160
rect 153580 10102 154271 10104
rect 153580 10100 153586 10102
rect 152825 10099 152891 10100
rect 154205 10099 154271 10102
rect 206318 10100 206324 10164
rect 206388 10162 206394 10164
rect 206553 10162 206619 10165
rect 206388 10160 206619 10162
rect 206388 10104 206558 10160
rect 206614 10104 206619 10160
rect 206388 10102 206619 10104
rect 206388 10100 206394 10102
rect 206553 10099 206619 10102
rect 207054 10100 207060 10164
rect 207124 10162 207130 10164
rect 207657 10162 207723 10165
rect 207124 10160 207723 10162
rect 207124 10104 207662 10160
rect 207718 10104 207723 10160
rect 207124 10102 207723 10104
rect 207124 10100 207130 10102
rect 207657 10099 207723 10102
rect 208526 10100 208532 10164
rect 208596 10162 208602 10164
rect 208945 10162 209011 10165
rect 209313 10164 209379 10165
rect 209262 10162 209268 10164
rect 208596 10160 209011 10162
rect 208596 10104 208950 10160
rect 209006 10104 209011 10160
rect 208596 10102 209011 10104
rect 209222 10102 209268 10162
rect 209332 10160 209379 10164
rect 209374 10104 209379 10160
rect 208596 10100 208602 10102
rect 208945 10099 209011 10102
rect 209262 10100 209268 10102
rect 209332 10100 209379 10104
rect 210734 10100 210740 10164
rect 210804 10162 210810 10164
rect 211153 10162 211219 10165
rect 210804 10160 211219 10162
rect 210804 10104 211158 10160
rect 211214 10104 211219 10160
rect 210804 10102 211219 10104
rect 210804 10100 210810 10102
rect 209313 10099 209379 10100
rect 211153 10099 211219 10102
rect 212206 10100 212212 10164
rect 212276 10162 212282 10164
rect 212533 10162 212599 10165
rect 212276 10160 212599 10162
rect 212276 10104 212538 10160
rect 212594 10104 212599 10160
rect 212276 10102 212599 10104
rect 212276 10100 212282 10102
rect 212533 10099 212599 10102
rect 213678 10100 213684 10164
rect 213748 10162 213754 10164
rect 213913 10162 213979 10165
rect 214465 10164 214531 10165
rect 214414 10162 214420 10164
rect 213748 10160 213979 10162
rect 213748 10104 213918 10160
rect 213974 10104 213979 10160
rect 213748 10102 213979 10104
rect 214374 10102 214420 10162
rect 214484 10160 214531 10164
rect 214526 10104 214531 10160
rect 213748 10100 213754 10102
rect 213913 10099 213979 10102
rect 214414 10100 214420 10102
rect 214484 10100 214531 10104
rect 215886 10100 215892 10164
rect 215956 10162 215962 10164
rect 216673 10162 216739 10165
rect 215956 10160 216739 10162
rect 215956 10104 216678 10160
rect 216734 10104 216739 10160
rect 215956 10102 216739 10104
rect 215956 10100 215962 10102
rect 214465 10099 214531 10100
rect 216673 10099 216739 10102
rect 217358 10100 217364 10164
rect 217428 10162 217434 10164
rect 217961 10162 218027 10165
rect 217428 10160 218027 10162
rect 217428 10104 217966 10160
rect 218022 10104 218027 10160
rect 217428 10102 218027 10104
rect 217428 10100 217434 10102
rect 217961 10099 218027 10102
rect 218830 10100 218836 10164
rect 218900 10162 218906 10164
rect 219249 10162 219315 10165
rect 218900 10160 219315 10162
rect 218900 10104 219254 10160
rect 219310 10104 219315 10160
rect 218900 10102 219315 10104
rect 218900 10100 218906 10102
rect 219249 10099 219315 10102
rect 219566 10100 219572 10164
rect 219636 10162 219642 10164
rect 220537 10162 220603 10165
rect 219636 10160 220603 10162
rect 219636 10104 220542 10160
rect 220598 10104 220603 10160
rect 219636 10102 220603 10104
rect 219636 10100 219642 10102
rect 220537 10099 220603 10102
rect 222510 10100 222516 10164
rect 222580 10162 222586 10164
rect 223113 10162 223179 10165
rect 222580 10160 223179 10162
rect 222580 10104 223118 10160
rect 223174 10104 223179 10160
rect 222580 10102 223179 10104
rect 222580 10100 222586 10102
rect 223113 10099 223179 10102
rect 223246 10100 223252 10164
rect 223316 10162 223322 10164
rect 223941 10162 224007 10165
rect 223316 10160 224007 10162
rect 223316 10104 223946 10160
rect 224002 10104 224007 10160
rect 223316 10102 224007 10104
rect 223316 10100 223322 10102
rect 223941 10099 224007 10102
rect 91134 9964 91140 10028
rect 91204 10026 91210 10028
rect 91645 10026 91711 10029
rect 91204 10024 91711 10026
rect 91204 9968 91650 10024
rect 91706 9968 91711 10024
rect 91204 9966 91711 9968
rect 91204 9964 91210 9966
rect 91645 9963 91711 9966
rect 268193 10026 268259 10029
rect 272149 10026 272215 10029
rect 268193 10024 272215 10026
rect 268193 9968 268198 10024
rect 268254 9968 272154 10024
rect 272210 9968 272215 10024
rect 268193 9966 272215 9968
rect 268193 9963 268259 9966
rect 272149 9963 272215 9966
rect 2998 9828 3004 9892
rect 3068 9890 3074 9892
rect 3141 9890 3207 9893
rect 8201 9892 8267 9893
rect 8150 9890 8156 9892
rect 3068 9888 3207 9890
rect 3068 9832 3146 9888
rect 3202 9832 3207 9888
rect 3068 9830 3207 9832
rect 8110 9830 8156 9890
rect 8220 9888 8267 9892
rect 8262 9832 8267 9888
rect 3068 9828 3074 9830
rect 3141 9827 3207 9830
rect 8150 9828 8156 9830
rect 8220 9828 8267 9832
rect 13302 9828 13308 9892
rect 13372 9890 13378 9892
rect 13445 9890 13511 9893
rect 13372 9888 13511 9890
rect 13372 9832 13450 9888
rect 13506 9832 13511 9888
rect 13372 9830 13511 9832
rect 13372 9828 13378 9830
rect 8201 9827 8267 9828
rect 13445 9827 13511 9830
rect 19926 9828 19932 9892
rect 19996 9890 20002 9892
rect 23197 9890 23263 9893
rect 19996 9888 23263 9890
rect 19996 9832 23202 9888
rect 23258 9832 23263 9888
rect 19996 9830 23263 9832
rect 19996 9828 20002 9830
rect 23197 9827 23263 9830
rect 69790 9828 69796 9892
rect 69860 9890 69866 9892
rect 70025 9890 70091 9893
rect 77201 9892 77267 9893
rect 78673 9892 78739 9893
rect 77150 9890 77156 9892
rect 69860 9888 70091 9890
rect 69860 9832 70030 9888
rect 70086 9832 70091 9888
rect 69860 9830 70091 9832
rect 77110 9830 77156 9890
rect 77220 9888 77267 9892
rect 78622 9890 78628 9892
rect 77262 9832 77267 9888
rect 69860 9828 69866 9830
rect 70025 9827 70091 9830
rect 77150 9828 77156 9830
rect 77220 9828 77267 9832
rect 78582 9830 78628 9890
rect 78692 9888 78739 9892
rect 78734 9832 78739 9888
rect 78622 9828 78628 9830
rect 78692 9828 78739 9832
rect 80830 9828 80836 9892
rect 80900 9890 80906 9892
rect 81249 9890 81315 9893
rect 80900 9888 81315 9890
rect 80900 9832 81254 9888
rect 81310 9832 81315 9888
rect 80900 9830 81315 9832
rect 80900 9828 80906 9830
rect 77201 9827 77267 9828
rect 78673 9827 78739 9828
rect 81249 9827 81315 9830
rect 85982 9828 85988 9892
rect 86052 9890 86058 9892
rect 86401 9890 86467 9893
rect 86052 9888 86467 9890
rect 86052 9832 86406 9888
rect 86462 9832 86467 9888
rect 86052 9830 86467 9832
rect 86052 9828 86058 9830
rect 86401 9827 86467 9830
rect 139526 9828 139532 9892
rect 139596 9890 139602 9892
rect 139761 9890 139827 9893
rect 139596 9888 139827 9890
rect 139596 9832 139766 9888
rect 139822 9832 139827 9888
rect 139596 9830 139827 9832
rect 139596 9828 139602 9830
rect 139761 9827 139827 9830
rect 144678 9828 144684 9892
rect 144748 9890 144754 9892
rect 144913 9890 144979 9893
rect 144748 9888 144979 9890
rect 144748 9832 144918 9888
rect 144974 9832 144979 9888
rect 144748 9830 144979 9832
rect 144748 9828 144754 9830
rect 144913 9827 144979 9830
rect 149830 9828 149836 9892
rect 149900 9890 149906 9892
rect 150065 9890 150131 9893
rect 149900 9888 150131 9890
rect 149900 9832 150070 9888
rect 150126 9832 150131 9888
rect 149900 9830 150131 9832
rect 149900 9828 149906 9830
rect 150065 9827 150131 9830
rect 154982 9828 154988 9892
rect 155052 9890 155058 9892
rect 155217 9890 155283 9893
rect 155052 9888 155283 9890
rect 155052 9832 155222 9888
rect 155278 9832 155283 9888
rect 155052 9830 155283 9832
rect 155052 9828 155058 9830
rect 155217 9827 155283 9830
rect 211470 9828 211476 9892
rect 211540 9890 211546 9892
rect 211705 9890 211771 9893
rect 211540 9888 211771 9890
rect 211540 9832 211710 9888
rect 211766 9832 211771 9888
rect 211540 9830 211771 9832
rect 211540 9828 211546 9830
rect 211705 9827 211771 9830
rect 216622 9828 216628 9892
rect 216692 9890 216698 9892
rect 216857 9890 216923 9893
rect 216692 9888 216923 9890
rect 216692 9832 216862 9888
rect 216918 9832 216923 9888
rect 216692 9830 216923 9832
rect 216692 9828 216698 9830
rect 216857 9827 216923 9830
rect 221774 9828 221780 9892
rect 221844 9890 221850 9892
rect 222009 9890 222075 9893
rect 221844 9888 222075 9890
rect 221844 9832 222014 9888
rect 222070 9832 222075 9888
rect 221844 9830 222075 9832
rect 221844 9828 221850 9830
rect 222009 9827 222075 9830
rect 68542 9824 68858 9825
rect 68542 9760 68548 9824
rect 68612 9760 68628 9824
rect 68692 9760 68708 9824
rect 68772 9760 68788 9824
rect 68852 9760 68858 9824
rect 68542 9759 68858 9760
rect 136139 9824 136455 9825
rect 136139 9760 136145 9824
rect 136209 9760 136225 9824
rect 136289 9760 136305 9824
rect 136369 9760 136385 9824
rect 136449 9760 136455 9824
rect 136139 9759 136455 9760
rect 203736 9824 204052 9825
rect 203736 9760 203742 9824
rect 203806 9760 203822 9824
rect 203886 9760 203902 9824
rect 203966 9760 203982 9824
rect 204046 9760 204052 9824
rect 203736 9759 204052 9760
rect 271333 9824 271649 9825
rect 271333 9760 271339 9824
rect 271403 9760 271419 9824
rect 271483 9760 271499 9824
rect 271563 9760 271579 9824
rect 271643 9760 271649 9824
rect 271333 9759 271649 9760
rect 25865 9756 25931 9757
rect 25814 9692 25820 9756
rect 25884 9754 25931 9756
rect 25884 9752 25976 9754
rect 25926 9696 25976 9752
rect 25884 9694 25976 9696
rect 25884 9692 25931 9694
rect 26550 9692 26556 9756
rect 26620 9754 26626 9756
rect 27337 9754 27403 9757
rect 26620 9752 27403 9754
rect 26620 9696 27342 9752
rect 27398 9696 27403 9752
rect 26620 9694 27403 9696
rect 26620 9692 26626 9694
rect 25865 9691 25931 9692
rect 27337 9691 27403 9694
rect 29085 9754 29151 9757
rect 30281 9756 30347 9757
rect 29494 9754 29500 9756
rect 29085 9752 29500 9754
rect 29085 9696 29090 9752
rect 29146 9696 29500 9752
rect 29085 9694 29500 9696
rect 29085 9691 29151 9694
rect 29494 9692 29500 9694
rect 29564 9692 29570 9756
rect 30230 9692 30236 9756
rect 30300 9754 30347 9756
rect 30300 9752 30392 9754
rect 30342 9696 30392 9752
rect 30300 9694 30392 9696
rect 30300 9692 30347 9694
rect 92606 9692 92612 9756
rect 92676 9754 92682 9756
rect 92749 9754 92815 9757
rect 92676 9752 92815 9754
rect 92676 9696 92754 9752
rect 92810 9696 92815 9752
rect 92676 9694 92815 9696
rect 92676 9692 92682 9694
rect 30281 9691 30347 9692
rect 92749 9691 92815 9694
rect 93342 9692 93348 9756
rect 93412 9754 93418 9756
rect 93485 9754 93551 9757
rect 93412 9752 93551 9754
rect 93412 9696 93490 9752
rect 93546 9696 93551 9752
rect 93412 9694 93551 9696
rect 93412 9692 93418 9694
rect 93485 9691 93551 9694
rect 95550 9692 95556 9756
rect 95620 9754 95626 9756
rect 96061 9754 96127 9757
rect 96337 9756 96403 9757
rect 95620 9752 96127 9754
rect 95620 9696 96066 9752
rect 96122 9696 96127 9752
rect 95620 9694 96127 9696
rect 95620 9692 95626 9694
rect 96061 9691 96127 9694
rect 96286 9692 96292 9756
rect 96356 9754 96403 9756
rect 96356 9752 96448 9754
rect 96398 9696 96448 9752
rect 96356 9694 96448 9696
rect 96356 9692 96403 9694
rect 98494 9692 98500 9756
rect 98564 9754 98570 9756
rect 99373 9754 99439 9757
rect 98564 9752 99439 9754
rect 98564 9696 99378 9752
rect 99434 9696 99439 9752
rect 98564 9694 99439 9696
rect 98564 9692 98570 9694
rect 96337 9691 96403 9692
rect 99373 9691 99439 9694
rect 99966 9692 99972 9756
rect 100036 9754 100042 9756
rect 100477 9754 100543 9757
rect 100036 9752 100543 9754
rect 100036 9696 100482 9752
rect 100538 9696 100543 9752
rect 100036 9694 100543 9696
rect 100036 9692 100042 9694
rect 100477 9691 100543 9694
rect 167494 9692 167500 9756
rect 167564 9754 167570 9756
rect 168373 9754 168439 9757
rect 167564 9752 168439 9754
rect 167564 9696 168378 9752
rect 168434 9696 168439 9752
rect 167564 9694 168439 9696
rect 167564 9692 167570 9694
rect 168373 9691 168439 9694
rect 168966 9692 168972 9756
rect 169036 9754 169042 9756
rect 169477 9754 169543 9757
rect 169036 9752 169543 9754
rect 169036 9696 169482 9752
rect 169538 9696 169543 9752
rect 169036 9694 169543 9696
rect 169036 9692 169042 9694
rect 169477 9691 169543 9694
rect 215201 9754 215267 9757
rect 268101 9754 268167 9757
rect 268837 9754 268903 9757
rect 215201 9752 268903 9754
rect 215201 9696 215206 9752
rect 215262 9696 268106 9752
rect 268162 9696 268842 9752
rect 268898 9696 268903 9752
rect 215201 9694 268903 9696
rect 215201 9691 215267 9694
rect 268101 9691 268167 9694
rect 268837 9691 268903 9694
rect 69105 9620 69171 9621
rect 69054 9556 69060 9620
rect 69124 9618 69171 9620
rect 70301 9618 70367 9621
rect 70526 9618 70532 9620
rect 69124 9616 69216 9618
rect 69166 9560 69216 9616
rect 69124 9558 69216 9560
rect 70301 9616 70532 9618
rect 70301 9560 70306 9616
rect 70362 9560 70532 9616
rect 70301 9558 70532 9560
rect 69124 9556 69171 9558
rect 69105 9555 69171 9556
rect 70301 9555 70367 9558
rect 70526 9556 70532 9558
rect 70596 9556 70602 9620
rect 72141 9618 72207 9621
rect 74257 9620 74323 9621
rect 72734 9618 72740 9620
rect 72141 9616 72740 9618
rect 72141 9560 72146 9616
rect 72202 9560 72740 9616
rect 72141 9558 72740 9560
rect 72141 9555 72207 9558
rect 72734 9556 72740 9558
rect 72804 9556 72810 9620
rect 74206 9618 74212 9620
rect 74166 9558 74212 9618
rect 74276 9616 74323 9620
rect 74318 9560 74323 9616
rect 74206 9556 74212 9558
rect 74276 9556 74323 9560
rect 74257 9555 74323 9556
rect 74717 9618 74783 9621
rect 76465 9620 76531 9621
rect 75678 9618 75684 9620
rect 74717 9616 75684 9618
rect 74717 9560 74722 9616
rect 74778 9560 75684 9616
rect 74717 9558 75684 9560
rect 74717 9555 74783 9558
rect 75678 9556 75684 9558
rect 75748 9556 75754 9620
rect 76414 9618 76420 9620
rect 76374 9558 76420 9618
rect 76484 9616 76531 9620
rect 76526 9560 76531 9616
rect 76414 9556 76420 9558
rect 76484 9556 76531 9560
rect 76465 9555 76531 9556
rect 77293 9618 77359 9621
rect 77886 9618 77892 9620
rect 77293 9616 77892 9618
rect 77293 9560 77298 9616
rect 77354 9560 77892 9616
rect 77293 9558 77892 9560
rect 77293 9555 77359 9558
rect 77886 9556 77892 9558
rect 77956 9556 77962 9620
rect 79961 9618 80027 9621
rect 80094 9618 80100 9620
rect 79961 9616 80100 9618
rect 79961 9560 79966 9616
rect 80022 9560 80100 9616
rect 79961 9558 80100 9560
rect 79961 9555 80027 9558
rect 80094 9556 80100 9558
rect 80164 9556 80170 9620
rect 137318 9556 137324 9620
rect 137388 9618 137394 9620
rect 138013 9618 138079 9621
rect 137388 9616 138079 9618
rect 137388 9560 138018 9616
rect 138074 9560 138079 9616
rect 137388 9558 138079 9560
rect 137388 9556 137394 9558
rect 138013 9555 138079 9558
rect 215150 9556 215156 9620
rect 215220 9618 215226 9620
rect 215477 9618 215543 9621
rect 215220 9616 215543 9618
rect 215220 9560 215482 9616
rect 215538 9560 215543 9616
rect 215220 9558 215543 9560
rect 215220 9556 215226 9558
rect 215477 9555 215543 9558
rect 270493 9618 270559 9621
rect 270493 9616 272504 9618
rect 270493 9560 270498 9616
rect 270554 9560 272504 9616
rect 270493 9558 272504 9560
rect 270493 9555 270559 9558
rect 89345 9482 89411 9485
rect 92013 9482 92079 9485
rect 89345 9480 92079 9482
rect 89345 9424 89350 9480
rect 89406 9424 92018 9480
rect 92074 9424 92079 9480
rect 89345 9422 92079 9424
rect 89345 9419 89411 9422
rect 92013 9419 92079 9422
rect 156454 9420 156460 9484
rect 156524 9482 156530 9484
rect 156689 9482 156755 9485
rect 224033 9484 224099 9485
rect 156524 9480 156755 9482
rect 156524 9424 156694 9480
rect 156750 9424 156755 9480
rect 156524 9422 156755 9424
rect 156524 9420 156530 9422
rect 156689 9419 156755 9422
rect 223982 9420 223988 9484
rect 224052 9482 224099 9484
rect 224052 9480 224144 9482
rect 224094 9424 224144 9480
rect 224052 9422 224144 9424
rect 224052 9420 224099 9422
rect 227662 9420 227668 9484
rect 227732 9482 227738 9484
rect 228265 9482 228331 9485
rect 227732 9480 228331 9482
rect 227732 9424 228270 9480
rect 228326 9424 228331 9480
rect 227732 9422 228331 9424
rect 227732 9420 227738 9422
rect 224033 9419 224099 9420
rect 228265 9419 228331 9422
rect 228398 9420 228404 9484
rect 228468 9482 228474 9484
rect 229001 9482 229067 9485
rect 229829 9484 229895 9485
rect 229829 9482 229876 9484
rect 228468 9480 229067 9482
rect 228468 9424 229006 9480
rect 229062 9424 229067 9480
rect 228468 9422 229067 9424
rect 229784 9480 229876 9482
rect 229784 9424 229834 9480
rect 229784 9422 229876 9424
rect 228468 9420 228474 9422
rect 229001 9419 229067 9422
rect 229829 9420 229876 9422
rect 229940 9420 229946 9484
rect 231945 9482 232011 9485
rect 232078 9482 232084 9484
rect 231945 9480 232084 9482
rect 231945 9424 231950 9480
rect 232006 9424 232084 9480
rect 231945 9422 232084 9424
rect 229829 9419 229895 9420
rect 231945 9419 232011 9422
rect 232078 9420 232084 9422
rect 232148 9420 232154 9484
rect 233417 9482 233483 9485
rect 233550 9482 233556 9484
rect 233417 9480 233556 9482
rect 233417 9424 233422 9480
rect 233478 9424 233556 9480
rect 233417 9422 233556 9424
rect 233417 9419 233483 9422
rect 233550 9420 233556 9422
rect 233620 9420 233626 9484
rect 235758 9420 235764 9484
rect 235828 9482 235834 9484
rect 235993 9482 236059 9485
rect 267549 9484 267615 9485
rect 267549 9482 267596 9484
rect 235828 9480 236059 9482
rect 235828 9424 235998 9480
rect 236054 9424 236059 9480
rect 235828 9422 236059 9424
rect 267504 9480 267596 9482
rect 267504 9424 267554 9480
rect 267504 9422 267596 9424
rect 235828 9420 235834 9422
rect 235993 9419 236059 9422
rect 267549 9420 267596 9422
rect 267660 9420 267666 9484
rect 267733 9482 267799 9485
rect 271965 9482 272031 9485
rect 267733 9480 272031 9482
rect 267733 9424 267738 9480
rect 267794 9424 271970 9480
rect 272026 9424 272031 9480
rect 267733 9422 272031 9424
rect 267549 9419 267615 9420
rect 267733 9419 267799 9422
rect 271965 9419 272031 9422
rect 272149 9482 272215 9485
rect 272149 9480 272504 9482
rect 272149 9424 272154 9480
rect 272210 9424 272504 9480
rect 272149 9422 272504 9424
rect 272149 9419 272215 9422
rect 268009 9346 268075 9349
rect 268009 9344 272504 9346
rect 268009 9288 268014 9344
rect 268070 9288 272504 9344
rect 268009 9286 272504 9288
rect 268009 9283 268075 9286
rect 34744 9280 35060 9281
rect 34744 9216 34750 9280
rect 34814 9216 34830 9280
rect 34894 9216 34910 9280
rect 34974 9216 34990 9280
rect 35054 9216 35060 9280
rect 34744 9215 35060 9216
rect 102341 9280 102657 9281
rect 102341 9216 102347 9280
rect 102411 9216 102427 9280
rect 102491 9216 102507 9280
rect 102571 9216 102587 9280
rect 102651 9216 102657 9280
rect 102341 9215 102657 9216
rect 169938 9280 170254 9281
rect 169938 9216 169944 9280
rect 170008 9216 170024 9280
rect 170088 9216 170104 9280
rect 170168 9216 170184 9280
rect 170248 9216 170254 9280
rect 169938 9215 170254 9216
rect 237535 9280 237851 9281
rect 237535 9216 237541 9280
rect 237605 9216 237621 9280
rect 237685 9216 237701 9280
rect 237765 9216 237781 9280
rect 237845 9216 237851 9280
rect 237535 9215 237851 9216
rect 790 9148 796 9212
rect 860 9210 866 9212
rect 1393 9210 1459 9213
rect 860 9208 1459 9210
rect 860 9152 1398 9208
rect 1454 9152 1459 9208
rect 860 9150 1459 9152
rect 860 9148 866 9150
rect 1393 9147 1459 9150
rect 23933 9210 23999 9213
rect 24342 9210 24348 9212
rect 23933 9208 24348 9210
rect 23933 9152 23938 9208
rect 23994 9152 24348 9208
rect 23933 9150 24348 9152
rect 23933 9147 23999 9150
rect 24342 9148 24348 9150
rect 24412 9148 24418 9212
rect 32438 9148 32444 9212
rect 32508 9210 32514 9212
rect 33041 9210 33107 9213
rect 88241 9212 88307 9213
rect 32508 9208 33107 9210
rect 32508 9152 33046 9208
rect 33102 9152 33107 9208
rect 32508 9150 33107 9152
rect 32508 9148 32514 9150
rect 33041 9147 33107 9150
rect 88190 9148 88196 9212
rect 88260 9210 88307 9212
rect 91737 9210 91803 9213
rect 91870 9210 91876 9212
rect 88260 9208 88352 9210
rect 88302 9152 88352 9208
rect 88260 9150 88352 9152
rect 91737 9208 91876 9210
rect 91737 9152 91742 9208
rect 91798 9152 91876 9208
rect 91737 9150 91876 9152
rect 88260 9148 88307 9150
rect 88241 9147 88307 9148
rect 91737 9147 91803 9150
rect 91870 9148 91876 9150
rect 91940 9148 91946 9212
rect 100702 9148 100708 9212
rect 100772 9210 100778 9212
rect 101213 9210 101279 9213
rect 100772 9208 101279 9210
rect 100772 9152 101218 9208
rect 101274 9152 101279 9208
rect 100772 9150 101279 9152
rect 100772 9148 100778 9150
rect 101213 9147 101279 9150
rect 168230 9148 168236 9212
rect 168300 9210 168306 9212
rect 169753 9210 169819 9213
rect 168300 9208 169819 9210
rect 168300 9152 169758 9208
rect 169814 9152 169819 9208
rect 168300 9150 169819 9152
rect 168300 9148 168306 9150
rect 169753 9147 169819 9150
rect 214005 9210 214071 9213
rect 228081 9210 228147 9213
rect 214005 9208 228147 9210
rect 214005 9152 214010 9208
rect 214066 9152 228086 9208
rect 228142 9152 228147 9208
rect 214005 9150 228147 9152
rect 214005 9147 214071 9150
rect 228081 9147 228147 9150
rect 236494 9148 236500 9212
rect 236564 9210 236570 9212
rect 236821 9210 236887 9213
rect 236564 9208 236887 9210
rect 236564 9152 236826 9208
rect 236882 9152 236887 9208
rect 236564 9150 236887 9152
rect 236564 9148 236570 9150
rect 236821 9147 236887 9150
rect 268745 9210 268811 9213
rect 268745 9208 272504 9210
rect 268745 9152 268750 9208
rect 268806 9152 272504 9208
rect 268745 9150 272504 9152
rect 268745 9147 268811 9150
rect 73429 9076 73495 9077
rect 73429 9074 73476 9076
rect 73384 9072 73476 9074
rect 73384 9016 73434 9072
rect 73384 9014 73476 9016
rect 73429 9012 73476 9014
rect 73540 9012 73546 9076
rect 74717 9074 74783 9077
rect 74942 9074 74948 9076
rect 74717 9072 74948 9074
rect 74717 9016 74722 9072
rect 74778 9016 74948 9072
rect 74717 9014 74948 9016
rect 73429 9011 73495 9012
rect 74717 9011 74783 9014
rect 74942 9012 74948 9014
rect 75012 9012 75018 9076
rect 96981 9074 97047 9077
rect 99281 9074 99347 9077
rect 96981 9072 99347 9074
rect 96981 9016 96986 9072
rect 97042 9016 99286 9072
rect 99342 9016 99347 9072
rect 96981 9014 99347 9016
rect 96981 9011 97047 9014
rect 99281 9011 99347 9014
rect 156045 9074 156111 9077
rect 157425 9074 157491 9077
rect 156045 9072 157491 9074
rect 156045 9016 156050 9072
rect 156106 9016 157430 9072
rect 157486 9016 157491 9072
rect 156045 9014 157491 9016
rect 156045 9011 156111 9014
rect 157425 9011 157491 9014
rect 163773 9074 163839 9077
rect 213862 9074 213868 9076
rect 163773 9072 213868 9074
rect 163773 9016 163778 9072
rect 163834 9016 213868 9072
rect 163773 9014 213868 9016
rect 163773 9011 163839 9014
rect 213862 9012 213868 9014
rect 213932 9012 213938 9076
rect 216765 9074 216831 9077
rect 227253 9074 227319 9077
rect 216765 9072 227319 9074
rect 216765 9016 216770 9072
rect 216826 9016 227258 9072
rect 227314 9016 227319 9072
rect 216765 9014 227319 9016
rect 216765 9011 216831 9014
rect 227253 9011 227319 9014
rect 232773 9074 232839 9077
rect 236729 9074 236795 9077
rect 232773 9072 236795 9074
rect 232773 9016 232778 9072
rect 232834 9016 236734 9072
rect 236790 9016 236795 9072
rect 232773 9014 236795 9016
rect 232773 9011 232839 9014
rect 236729 9011 236795 9014
rect 268653 9074 268719 9077
rect 268653 9072 272504 9074
rect 268653 9016 268658 9072
rect 268714 9016 272504 9072
rect 268653 9014 272504 9016
rect 268653 9011 268719 9014
rect 22093 8940 22159 8941
rect 22093 8936 22140 8940
rect 22204 8938 22210 8940
rect 22093 8880 22098 8936
rect 22093 8876 22140 8880
rect 22204 8878 22250 8938
rect 22204 8876 22210 8878
rect 96286 8876 96292 8940
rect 96356 8938 96362 8940
rect 96521 8938 96587 8941
rect 96356 8936 96587 8938
rect 96356 8880 96526 8936
rect 96582 8880 96587 8936
rect 96356 8878 96587 8880
rect 96356 8876 96362 8878
rect 22093 8875 22159 8876
rect 96521 8875 96587 8878
rect 98545 8938 98611 8941
rect 99465 8938 99531 8941
rect 227478 8938 227484 8940
rect 98545 8936 99531 8938
rect 98545 8880 98550 8936
rect 98606 8880 99470 8936
rect 99526 8880 99531 8936
rect 98545 8878 99531 8880
rect 98545 8875 98611 8878
rect 99465 8875 99531 8878
rect 220126 8878 227484 8938
rect 68542 8736 68858 8737
rect 68542 8672 68548 8736
rect 68612 8672 68628 8736
rect 68692 8672 68708 8736
rect 68772 8672 68788 8736
rect 68852 8672 68858 8736
rect 68542 8671 68858 8672
rect 136139 8736 136455 8737
rect 136139 8672 136145 8736
rect 136209 8672 136225 8736
rect 136289 8672 136305 8736
rect 136369 8672 136385 8736
rect 136449 8672 136455 8736
rect 136139 8671 136455 8672
rect 203736 8736 204052 8737
rect 203736 8672 203742 8736
rect 203806 8672 203822 8736
rect 203886 8672 203902 8736
rect 203966 8672 203982 8736
rect 204046 8672 204052 8736
rect 203736 8671 204052 8672
rect 21357 8668 21423 8669
rect 21357 8666 21404 8668
rect 21312 8664 21404 8666
rect 21312 8608 21362 8664
rect 21312 8606 21404 8608
rect 21357 8604 21404 8606
rect 21468 8604 21474 8668
rect 27286 8604 27292 8668
rect 27356 8666 27362 8668
rect 27429 8666 27495 8669
rect 27356 8664 27495 8666
rect 27356 8608 27434 8664
rect 27490 8608 27495 8664
rect 27356 8606 27495 8608
rect 27356 8604 27362 8606
rect 21357 8603 21423 8604
rect 27429 8603 27495 8606
rect 28022 8604 28028 8668
rect 28092 8666 28098 8668
rect 28165 8666 28231 8669
rect 28092 8664 28231 8666
rect 28092 8608 28170 8664
rect 28226 8608 28231 8664
rect 28092 8606 28231 8608
rect 28092 8604 28098 8606
rect 28165 8603 28231 8606
rect 28758 8604 28764 8668
rect 28828 8666 28834 8668
rect 28901 8666 28967 8669
rect 31017 8668 31083 8669
rect 87505 8668 87571 8669
rect 28828 8664 28967 8666
rect 28828 8608 28906 8664
rect 28962 8608 28967 8664
rect 28828 8606 28967 8608
rect 28828 8604 28834 8606
rect 28901 8603 28967 8606
rect 30966 8604 30972 8668
rect 31036 8666 31083 8668
rect 31036 8664 31128 8666
rect 31078 8608 31128 8664
rect 31036 8606 31128 8608
rect 31036 8604 31083 8606
rect 87454 8604 87460 8668
rect 87524 8666 87571 8668
rect 87524 8664 87616 8666
rect 87566 8608 87616 8664
rect 87524 8606 87616 8608
rect 87524 8604 87571 8606
rect 90398 8604 90404 8668
rect 90468 8666 90474 8668
rect 90817 8666 90883 8669
rect 90468 8664 90883 8666
rect 90468 8608 90822 8664
rect 90878 8608 90883 8664
rect 90468 8606 90883 8608
rect 90468 8604 90474 8606
rect 31017 8603 31083 8604
rect 87505 8603 87571 8604
rect 90817 8603 90883 8606
rect 94078 8604 94084 8668
rect 94148 8666 94154 8668
rect 94589 8666 94655 8669
rect 94148 8664 94655 8666
rect 94148 8608 94594 8664
rect 94650 8608 94655 8664
rect 94148 8606 94655 8608
rect 94148 8604 94154 8606
rect 94589 8603 94655 8606
rect 94814 8604 94820 8668
rect 94884 8666 94890 8668
rect 95049 8666 95115 8669
rect 94884 8664 95115 8666
rect 94884 8608 95054 8664
rect 95110 8608 95115 8664
rect 94884 8606 95115 8608
rect 94884 8604 94890 8606
rect 95049 8603 95115 8606
rect 97022 8604 97028 8668
rect 97092 8666 97098 8668
rect 97533 8666 97599 8669
rect 97092 8664 97599 8666
rect 97092 8608 97538 8664
rect 97594 8608 97599 8664
rect 97092 8606 97599 8608
rect 97092 8604 97098 8606
rect 97533 8603 97599 8606
rect 97758 8604 97764 8668
rect 97828 8666 97834 8668
rect 97993 8666 98059 8669
rect 97828 8664 98059 8666
rect 97828 8608 97998 8664
rect 98054 8608 98059 8664
rect 97828 8606 98059 8608
rect 97828 8604 97834 8606
rect 97993 8603 98059 8606
rect 99230 8604 99236 8668
rect 99300 8666 99306 8668
rect 99373 8666 99439 8669
rect 99300 8664 99439 8666
rect 99300 8608 99378 8664
rect 99434 8608 99439 8664
rect 99300 8606 99439 8608
rect 99300 8604 99306 8606
rect 99373 8603 99439 8606
rect 155718 8604 155724 8668
rect 155788 8666 155794 8668
rect 156045 8666 156111 8669
rect 220126 8666 220186 8878
rect 227478 8876 227484 8878
rect 227548 8876 227554 8940
rect 269021 8938 269087 8941
rect 271965 8938 272031 8941
rect 269021 8936 271890 8938
rect 269021 8880 269026 8936
rect 269082 8880 271890 8936
rect 269021 8878 271890 8880
rect 269021 8875 269087 8878
rect 220537 8802 220603 8805
rect 226006 8802 226012 8804
rect 220537 8800 226012 8802
rect 220537 8744 220542 8800
rect 220598 8744 226012 8800
rect 220537 8742 226012 8744
rect 220537 8739 220603 8742
rect 226006 8740 226012 8742
rect 226076 8740 226082 8804
rect 232497 8802 232563 8805
rect 235993 8802 236059 8805
rect 232497 8800 236059 8802
rect 232497 8744 232502 8800
rect 232558 8744 235998 8800
rect 236054 8744 236059 8800
rect 232497 8742 236059 8744
rect 271830 8802 271890 8878
rect 271965 8936 272504 8938
rect 271965 8880 271970 8936
rect 272026 8880 272504 8936
rect 271965 8878 272504 8880
rect 271965 8875 272031 8878
rect 271830 8742 272504 8802
rect 232497 8739 232563 8742
rect 235993 8739 236059 8742
rect 271333 8736 271649 8737
rect 271333 8672 271339 8736
rect 271403 8672 271419 8736
rect 271483 8672 271499 8736
rect 271563 8672 271579 8736
rect 271643 8672 271649 8736
rect 271333 8671 271649 8672
rect 224677 8668 224743 8669
rect 225505 8668 225571 8669
rect 226241 8668 226307 8669
rect 226977 8668 227043 8669
rect 229185 8668 229251 8669
rect 224677 8666 224724 8668
rect 155788 8664 156111 8666
rect 155788 8608 156050 8664
rect 156106 8608 156111 8664
rect 155788 8606 156111 8608
rect 155788 8604 155794 8606
rect 156045 8603 156111 8606
rect 214192 8606 220186 8666
rect 224632 8664 224724 8666
rect 224632 8608 224682 8664
rect 224632 8606 224724 8608
rect 95233 8530 95299 8533
rect 95877 8530 95943 8533
rect 95233 8528 95943 8530
rect 95233 8472 95238 8528
rect 95294 8472 95882 8528
rect 95938 8472 95943 8528
rect 95233 8470 95943 8472
rect 95233 8467 95299 8470
rect 95877 8467 95943 8470
rect 97165 8530 97231 8533
rect 98913 8530 98979 8533
rect 100293 8530 100359 8533
rect 97165 8528 100359 8530
rect 97165 8472 97170 8528
rect 97226 8472 98918 8528
rect 98974 8472 100298 8528
rect 100354 8472 100359 8528
rect 97165 8470 100359 8472
rect 97165 8467 97231 8470
rect 98913 8467 98979 8470
rect 100293 8467 100359 8470
rect 145097 8530 145163 8533
rect 157701 8530 157767 8533
rect 145097 8528 157767 8530
rect 145097 8472 145102 8528
rect 145158 8472 157706 8528
rect 157762 8472 157767 8528
rect 145097 8470 157767 8472
rect 145097 8467 145163 8470
rect 157701 8467 157767 8470
rect 20662 8332 20668 8396
rect 20732 8394 20738 8396
rect 21909 8394 21975 8397
rect 22921 8396 22987 8397
rect 23657 8396 23723 8397
rect 20732 8392 21975 8394
rect 20732 8336 21914 8392
rect 21970 8336 21975 8392
rect 20732 8334 21975 8336
rect 20732 8332 20738 8334
rect 21909 8331 21975 8334
rect 22870 8332 22876 8396
rect 22940 8394 22987 8396
rect 22940 8392 23032 8394
rect 22982 8336 23032 8392
rect 22940 8334 23032 8336
rect 22940 8332 22987 8334
rect 23606 8332 23612 8396
rect 23676 8394 23723 8396
rect 23676 8392 23768 8394
rect 23718 8336 23768 8392
rect 23676 8334 23768 8336
rect 23676 8332 23723 8334
rect 25078 8332 25084 8396
rect 25148 8394 25154 8396
rect 25221 8394 25287 8397
rect 25148 8392 25287 8394
rect 25148 8336 25226 8392
rect 25282 8336 25287 8392
rect 25148 8334 25287 8336
rect 25148 8332 25154 8334
rect 22921 8331 22987 8332
rect 23657 8331 23723 8332
rect 25221 8331 25287 8334
rect 99097 8394 99163 8397
rect 100661 8394 100727 8397
rect 157241 8396 157307 8397
rect 157190 8394 157196 8396
rect 99097 8392 100727 8394
rect 99097 8336 99102 8392
rect 99158 8336 100666 8392
rect 100722 8336 100727 8392
rect 99097 8334 100727 8336
rect 157150 8334 157196 8394
rect 157260 8392 157307 8396
rect 157302 8336 157307 8392
rect 99097 8331 99163 8334
rect 100661 8331 100727 8334
rect 157190 8332 157196 8334
rect 157260 8332 157307 8336
rect 158662 8332 158668 8396
rect 158732 8394 158738 8396
rect 159357 8394 159423 8397
rect 158732 8392 159423 8394
rect 158732 8336 159362 8392
rect 159418 8336 159423 8392
rect 158732 8334 159423 8336
rect 158732 8332 158738 8334
rect 157241 8331 157307 8332
rect 159357 8331 159423 8334
rect 160134 8332 160140 8396
rect 160204 8394 160210 8396
rect 160921 8394 160987 8397
rect 160204 8392 160987 8394
rect 160204 8336 160926 8392
rect 160982 8336 160987 8392
rect 160204 8334 160987 8336
rect 160204 8332 160210 8334
rect 160921 8331 160987 8334
rect 161606 8332 161612 8396
rect 161676 8394 161682 8396
rect 162393 8394 162459 8397
rect 161676 8392 162459 8394
rect 161676 8336 162398 8392
rect 162454 8336 162459 8392
rect 161676 8334 162459 8336
rect 161676 8332 161682 8334
rect 162393 8331 162459 8334
rect 163078 8332 163084 8396
rect 163148 8394 163154 8396
rect 163865 8394 163931 8397
rect 163148 8392 163931 8394
rect 163148 8336 163870 8392
rect 163926 8336 163931 8392
rect 163148 8334 163931 8336
rect 163148 8332 163154 8334
rect 163865 8331 163931 8334
rect 164550 8332 164556 8396
rect 164620 8394 164626 8396
rect 165245 8394 165311 8397
rect 164620 8392 165311 8394
rect 164620 8336 165250 8392
rect 165306 8336 165311 8392
rect 164620 8334 165311 8336
rect 164620 8332 164626 8334
rect 165245 8331 165311 8334
rect 166022 8332 166028 8396
rect 166092 8394 166098 8396
rect 166533 8394 166599 8397
rect 166092 8392 166599 8394
rect 166092 8336 166538 8392
rect 166594 8336 166599 8392
rect 166092 8334 166599 8336
rect 166092 8332 166098 8334
rect 166533 8331 166599 8334
rect 166758 8332 166764 8396
rect 166828 8394 166834 8396
rect 166901 8394 166967 8397
rect 166828 8392 166967 8394
rect 166828 8336 166906 8392
rect 166962 8336 166967 8392
rect 166828 8334 166967 8336
rect 166828 8332 166834 8334
rect 166901 8331 166967 8334
rect 95969 8258 96035 8261
rect 102041 8258 102107 8261
rect 95969 8256 102107 8258
rect 95969 8200 95974 8256
rect 96030 8200 102046 8256
rect 102102 8200 102107 8256
rect 95969 8198 102107 8200
rect 95969 8195 96035 8198
rect 102041 8195 102107 8198
rect 103421 8258 103487 8261
rect 106273 8258 106339 8261
rect 103421 8256 106339 8258
rect 103421 8200 103426 8256
rect 103482 8200 106278 8256
rect 106334 8200 106339 8256
rect 103421 8198 106339 8200
rect 103421 8195 103487 8198
rect 106273 8195 106339 8198
rect 171041 8258 171107 8261
rect 179413 8258 179479 8261
rect 171041 8256 179479 8258
rect 171041 8200 171046 8256
rect 171102 8200 179418 8256
rect 179474 8200 179479 8256
rect 171041 8198 179479 8200
rect 171041 8195 171107 8198
rect 179413 8195 179479 8198
rect 195329 8258 195395 8261
rect 214005 8258 214071 8261
rect 195329 8256 214071 8258
rect 195329 8200 195334 8256
rect 195390 8200 214010 8256
rect 214066 8200 214071 8256
rect 195329 8198 214071 8200
rect 195329 8195 195395 8198
rect 214005 8195 214071 8198
rect 34744 8192 35060 8193
rect 34744 8128 34750 8192
rect 34814 8128 34830 8192
rect 34894 8128 34910 8192
rect 34974 8128 34990 8192
rect 35054 8128 35060 8192
rect 34744 8127 35060 8128
rect 102341 8192 102657 8193
rect 102341 8128 102347 8192
rect 102411 8128 102427 8192
rect 102491 8128 102507 8192
rect 102571 8128 102587 8192
rect 102651 8128 102657 8192
rect 102341 8127 102657 8128
rect 169938 8192 170254 8193
rect 169938 8128 169944 8192
rect 170008 8128 170024 8192
rect 170088 8128 170104 8192
rect 170168 8128 170184 8192
rect 170248 8128 170254 8192
rect 169938 8127 170254 8128
rect 214192 8125 214252 8606
rect 224677 8604 224724 8606
rect 224788 8604 224794 8668
rect 225454 8604 225460 8668
rect 225524 8666 225571 8668
rect 225524 8664 225616 8666
rect 225566 8608 225616 8664
rect 225524 8606 225616 8608
rect 225524 8604 225571 8606
rect 226190 8604 226196 8668
rect 226260 8666 226307 8668
rect 226260 8664 226352 8666
rect 226302 8608 226352 8664
rect 226260 8606 226352 8608
rect 226260 8604 226307 8606
rect 226926 8604 226932 8668
rect 226996 8666 227043 8668
rect 226996 8664 227088 8666
rect 227038 8608 227088 8664
rect 226996 8606 227088 8608
rect 226996 8604 227043 8606
rect 229134 8604 229140 8668
rect 229204 8666 229251 8668
rect 229204 8664 229296 8666
rect 229246 8608 229296 8664
rect 229204 8606 229296 8608
rect 229204 8604 229251 8606
rect 230606 8604 230612 8668
rect 230676 8666 230682 8668
rect 230933 8666 230999 8669
rect 230676 8664 230999 8666
rect 230676 8608 230938 8664
rect 230994 8608 230999 8664
rect 230676 8606 230999 8608
rect 230676 8604 230682 8606
rect 224677 8603 224743 8604
rect 225505 8603 225571 8604
rect 226241 8603 226307 8604
rect 226977 8603 227043 8604
rect 229185 8603 229251 8604
rect 230933 8603 230999 8606
rect 231342 8604 231348 8668
rect 231412 8666 231418 8668
rect 231669 8666 231735 8669
rect 231412 8664 231735 8666
rect 231412 8608 231674 8664
rect 231730 8608 231735 8664
rect 231412 8606 231735 8608
rect 231412 8604 231418 8606
rect 231669 8603 231735 8606
rect 232589 8666 232655 8669
rect 232814 8666 232820 8668
rect 232589 8664 232820 8666
rect 232589 8608 232594 8664
rect 232650 8608 232820 8664
rect 232589 8606 232820 8608
rect 232589 8603 232655 8606
rect 232814 8604 232820 8606
rect 232884 8604 232890 8668
rect 234286 8604 234292 8668
rect 234356 8666 234362 8668
rect 234429 8666 234495 8669
rect 234356 8664 234495 8666
rect 234356 8608 234434 8664
rect 234490 8608 234495 8664
rect 234356 8606 234495 8608
rect 234356 8604 234362 8606
rect 234429 8603 234495 8606
rect 236269 8666 236335 8669
rect 237230 8666 237236 8668
rect 236269 8664 237236 8666
rect 236269 8608 236274 8664
rect 236330 8608 237236 8664
rect 236269 8606 237236 8608
rect 236269 8603 236335 8606
rect 237230 8604 237236 8606
rect 237300 8604 237306 8668
rect 272304 8606 272504 8666
rect 220813 8530 220879 8533
rect 227294 8530 227300 8532
rect 220813 8528 227300 8530
rect 220813 8472 220818 8528
rect 220874 8472 227300 8528
rect 220813 8470 227300 8472
rect 220813 8467 220879 8470
rect 227294 8468 227300 8470
rect 227364 8468 227370 8532
rect 268285 8530 268351 8533
rect 268285 8528 272504 8530
rect 268285 8472 268290 8528
rect 268346 8472 272504 8528
rect 268285 8470 272504 8472
rect 268285 8467 268351 8470
rect 217317 8394 217383 8397
rect 223297 8394 223363 8397
rect 217317 8392 223363 8394
rect 217317 8336 217322 8392
rect 217378 8336 223302 8392
rect 223358 8336 223363 8392
rect 217317 8334 223363 8336
rect 217317 8331 217383 8334
rect 223297 8331 223363 8334
rect 224309 8396 224375 8397
rect 224309 8392 224356 8396
rect 224420 8394 224426 8396
rect 232313 8394 232379 8397
rect 234429 8394 234495 8397
rect 224309 8336 224314 8392
rect 224309 8332 224356 8336
rect 224420 8334 224466 8394
rect 232313 8392 234495 8394
rect 232313 8336 232318 8392
rect 232374 8336 234434 8392
rect 234490 8336 234495 8392
rect 232313 8334 234495 8336
rect 224420 8332 224426 8334
rect 224309 8331 224375 8332
rect 232313 8331 232379 8334
rect 234429 8331 234495 8334
rect 234889 8394 234955 8397
rect 235022 8394 235028 8396
rect 234889 8392 235028 8394
rect 234889 8336 234894 8392
rect 234950 8336 235028 8392
rect 234889 8334 235028 8336
rect 234889 8331 234955 8334
rect 235022 8332 235028 8334
rect 235092 8332 235098 8396
rect 263869 8394 263935 8397
rect 267273 8394 267339 8397
rect 263869 8392 267339 8394
rect 263869 8336 263874 8392
rect 263930 8336 267278 8392
rect 267334 8336 267339 8392
rect 263869 8334 267339 8336
rect 263869 8331 263935 8334
rect 267273 8331 267339 8334
rect 268009 8394 268075 8397
rect 268009 8392 272504 8394
rect 268009 8336 268014 8392
rect 268070 8336 272504 8392
rect 268009 8334 272504 8336
rect 268009 8331 268075 8334
rect 216581 8258 216647 8261
rect 224861 8258 224927 8261
rect 262581 8258 262647 8261
rect 216581 8256 224927 8258
rect 216581 8200 216586 8256
rect 216642 8200 224866 8256
rect 224922 8200 224927 8256
rect 216581 8198 224927 8200
rect 216581 8195 216647 8198
rect 224861 8195 224927 8198
rect 239446 8256 262647 8258
rect 239446 8200 262586 8256
rect 262642 8200 262647 8256
rect 239446 8198 262647 8200
rect 237535 8192 237851 8193
rect 237535 8128 237541 8192
rect 237605 8128 237621 8192
rect 237685 8128 237701 8192
rect 237765 8128 237781 8192
rect 237845 8128 237851 8192
rect 237535 8127 237851 8128
rect 88926 8060 88932 8124
rect 88996 8122 89002 8124
rect 89713 8122 89779 8125
rect 88996 8120 89779 8122
rect 88996 8064 89718 8120
rect 89774 8064 89779 8120
rect 88996 8062 89779 8064
rect 88996 8060 89002 8062
rect 89713 8059 89779 8062
rect 94313 8122 94379 8125
rect 96838 8122 96844 8124
rect 94313 8120 96844 8122
rect 94313 8064 94318 8120
rect 94374 8064 96844 8120
rect 94313 8062 96844 8064
rect 94313 8059 94379 8062
rect 96838 8060 96844 8062
rect 96908 8060 96914 8124
rect 113817 8122 113883 8125
rect 154757 8122 154823 8125
rect 113817 8120 154823 8122
rect 113817 8064 113822 8120
rect 113878 8064 154762 8120
rect 154818 8064 154823 8120
rect 113817 8062 154823 8064
rect 113817 8059 113883 8062
rect 154757 8059 154823 8062
rect 157926 8060 157932 8124
rect 157996 8122 158002 8124
rect 158713 8122 158779 8125
rect 159449 8124 159515 8125
rect 157996 8120 158779 8122
rect 157996 8064 158718 8120
rect 158774 8064 158779 8120
rect 157996 8062 158779 8064
rect 157996 8060 158002 8062
rect 158713 8059 158779 8062
rect 159398 8060 159404 8124
rect 159468 8122 159515 8124
rect 159468 8120 159560 8122
rect 159510 8064 159560 8120
rect 159468 8062 159560 8064
rect 159468 8060 159515 8062
rect 160870 8060 160876 8124
rect 160940 8122 160946 8124
rect 161013 8122 161079 8125
rect 160940 8120 161079 8122
rect 160940 8064 161018 8120
rect 161074 8064 161079 8120
rect 160940 8062 161079 8064
rect 160940 8060 160946 8062
rect 159449 8059 159515 8060
rect 161013 8059 161079 8062
rect 161197 8122 161263 8125
rect 163313 8122 163379 8125
rect 161197 8120 163379 8122
rect 161197 8064 161202 8120
rect 161258 8064 163318 8120
rect 163374 8064 163379 8120
rect 161197 8062 163379 8064
rect 161197 8059 161263 8062
rect 163313 8059 163379 8062
rect 163814 8060 163820 8124
rect 163884 8122 163890 8124
rect 163957 8122 164023 8125
rect 165337 8124 165403 8125
rect 163884 8120 164023 8122
rect 163884 8064 163962 8120
rect 164018 8064 164023 8120
rect 163884 8062 164023 8064
rect 163884 8060 163890 8062
rect 163957 8059 164023 8062
rect 165286 8060 165292 8124
rect 165356 8122 165403 8124
rect 214189 8122 214255 8125
rect 165356 8120 165448 8122
rect 165398 8064 165448 8120
rect 165356 8062 165448 8064
rect 195930 8120 214255 8122
rect 195930 8064 214194 8120
rect 214250 8064 214255 8120
rect 195930 8062 214255 8064
rect 165356 8060 165403 8062
rect 165337 8059 165403 8060
rect 52177 7986 52243 7989
rect 116945 7986 117011 7989
rect 52177 7984 117011 7986
rect 52177 7928 52182 7984
rect 52238 7928 116950 7984
rect 117006 7928 117011 7984
rect 52177 7926 117011 7928
rect 52177 7923 52243 7926
rect 116945 7923 117011 7926
rect 149973 7986 150039 7989
rect 195930 7986 195990 8062
rect 214189 8059 214255 8062
rect 223205 8122 223271 8125
rect 224585 8122 224651 8125
rect 237373 8122 237439 8125
rect 223205 8120 224050 8122
rect 223205 8064 223210 8120
rect 223266 8064 224050 8120
rect 223205 8062 224050 8064
rect 223205 8059 223271 8062
rect 223757 7986 223823 7989
rect 149973 7984 195990 7986
rect 149973 7928 149978 7984
rect 150034 7928 195990 7984
rect 149973 7926 195990 7928
rect 215250 7984 223823 7986
rect 215250 7928 223762 7984
rect 223818 7928 223823 7984
rect 215250 7926 223823 7928
rect 223990 7986 224050 8062
rect 224585 8120 237439 8122
rect 224585 8064 224590 8120
rect 224646 8064 237378 8120
rect 237434 8064 237439 8120
rect 224585 8062 237439 8064
rect 224585 8059 224651 8062
rect 237373 8059 237439 8062
rect 226149 7986 226215 7989
rect 223990 7984 226215 7986
rect 223990 7928 226154 7984
rect 226210 7928 226215 7984
rect 223990 7926 226215 7928
rect 149973 7923 150039 7926
rect 85481 7850 85547 7853
rect 96613 7850 96679 7853
rect 114001 7850 114067 7853
rect 85481 7848 94514 7850
rect 85481 7792 85486 7848
rect 85542 7792 94514 7848
rect 85481 7790 94514 7792
rect 85481 7787 85547 7790
rect 75821 7714 75887 7717
rect 94313 7714 94379 7717
rect 75821 7712 94379 7714
rect 75821 7656 75826 7712
rect 75882 7656 94318 7712
rect 94374 7656 94379 7712
rect 75821 7654 94379 7656
rect 94454 7714 94514 7790
rect 96613 7848 114067 7850
rect 96613 7792 96618 7848
rect 96674 7792 114006 7848
rect 114062 7792 114067 7848
rect 96613 7790 114067 7792
rect 96613 7787 96679 7790
rect 114001 7787 114067 7790
rect 120257 7850 120323 7853
rect 156045 7850 156111 7853
rect 162393 7852 162459 7853
rect 120257 7848 156111 7850
rect 120257 7792 120262 7848
rect 120318 7792 156050 7848
rect 156106 7792 156111 7848
rect 120257 7790 156111 7792
rect 120257 7787 120323 7790
rect 156045 7787 156111 7790
rect 162342 7788 162348 7852
rect 162412 7850 162459 7852
rect 163313 7850 163379 7853
rect 170765 7850 170831 7853
rect 162412 7848 162504 7850
rect 162454 7792 162504 7848
rect 162412 7790 162504 7792
rect 163313 7848 170831 7850
rect 163313 7792 163318 7848
rect 163374 7792 170770 7848
rect 170826 7792 170831 7848
rect 163313 7790 170831 7792
rect 162412 7788 162459 7790
rect 162393 7787 162459 7788
rect 163313 7787 163379 7790
rect 170765 7787 170831 7790
rect 213913 7850 213979 7853
rect 215250 7850 215310 7926
rect 223757 7923 223823 7926
rect 226149 7923 226215 7926
rect 228357 7986 228423 7989
rect 239446 7986 239506 8198
rect 262581 8195 262647 8198
rect 263961 8258 264027 8261
rect 271781 8258 271847 8261
rect 263961 8256 271847 8258
rect 263961 8200 263966 8256
rect 264022 8200 271786 8256
rect 271842 8200 271847 8256
rect 263961 8198 271847 8200
rect 263961 8195 264027 8198
rect 271781 8195 271847 8198
rect 272014 8198 272504 8258
rect 245193 8122 245259 8125
rect 228357 7984 239506 7986
rect 228357 7928 228362 7984
rect 228418 7928 239506 7984
rect 228357 7926 239506 7928
rect 244230 8120 245259 8122
rect 244230 8064 245198 8120
rect 245254 8064 245259 8120
rect 244230 8062 245259 8064
rect 228357 7923 228423 7926
rect 213913 7848 215310 7850
rect 213913 7792 213918 7848
rect 213974 7792 215310 7848
rect 213913 7790 215310 7792
rect 219433 7850 219499 7853
rect 225505 7850 225571 7853
rect 219433 7848 225571 7850
rect 219433 7792 219438 7848
rect 219494 7792 225510 7848
rect 225566 7792 225571 7848
rect 219433 7790 225571 7792
rect 213913 7787 213979 7790
rect 219433 7787 219499 7790
rect 225505 7787 225571 7790
rect 226241 7850 226307 7853
rect 244230 7850 244290 8062
rect 245193 8059 245259 8062
rect 246941 8122 247007 8125
rect 260833 8122 260899 8125
rect 264881 8124 264947 8125
rect 246941 8120 260899 8122
rect 246941 8064 246946 8120
rect 247002 8064 260838 8120
rect 260894 8064 260899 8120
rect 246941 8062 260899 8064
rect 246941 8059 247007 8062
rect 260833 8059 260899 8062
rect 264830 8060 264836 8124
rect 264900 8122 264947 8124
rect 268285 8122 268351 8125
rect 272014 8122 272074 8198
rect 264900 8120 264992 8122
rect 264942 8064 264992 8120
rect 264900 8062 264992 8064
rect 268285 8120 272074 8122
rect 268285 8064 268290 8120
rect 268346 8064 272074 8120
rect 268285 8062 272074 8064
rect 272149 8122 272215 8125
rect 272149 8120 272504 8122
rect 272149 8064 272154 8120
rect 272210 8064 272504 8120
rect 272149 8062 272504 8064
rect 264900 8060 264947 8062
rect 264881 8059 264947 8060
rect 268285 8059 268351 8062
rect 272149 8059 272215 8062
rect 250161 7986 250227 7989
rect 254117 7986 254183 7989
rect 250161 7984 254183 7986
rect 250161 7928 250166 7984
rect 250222 7928 254122 7984
rect 254178 7928 254183 7984
rect 250161 7926 254183 7928
rect 250161 7923 250227 7926
rect 254117 7923 254183 7926
rect 262213 7986 262279 7989
rect 267733 7986 267799 7989
rect 262213 7984 267799 7986
rect 262213 7928 262218 7984
rect 262274 7928 267738 7984
rect 267794 7928 267799 7984
rect 262213 7926 267799 7928
rect 262213 7923 262279 7926
rect 267733 7923 267799 7926
rect 268009 7986 268075 7989
rect 271781 7986 271847 7989
rect 268009 7984 271847 7986
rect 268009 7928 268014 7984
rect 268070 7928 271786 7984
rect 271842 7928 271847 7984
rect 268009 7926 271847 7928
rect 268009 7923 268075 7926
rect 271781 7923 271847 7926
rect 272149 7986 272215 7989
rect 272149 7984 272504 7986
rect 272149 7928 272154 7984
rect 272210 7928 272504 7984
rect 272149 7926 272504 7928
rect 272149 7923 272215 7926
rect 226241 7848 244290 7850
rect 226241 7792 226246 7848
rect 226302 7792 244290 7848
rect 226241 7790 244290 7792
rect 264881 7850 264947 7853
rect 264881 7848 272504 7850
rect 264881 7792 264886 7848
rect 264942 7792 272504 7848
rect 264881 7790 272504 7792
rect 226241 7787 226307 7790
rect 264881 7787 264947 7790
rect 102869 7714 102935 7717
rect 94454 7712 102935 7714
rect 94454 7656 102874 7712
rect 102930 7656 102935 7712
rect 94454 7654 102935 7656
rect 75821 7651 75887 7654
rect 94313 7651 94379 7654
rect 102869 7651 102935 7654
rect 154573 7714 154639 7717
rect 172513 7714 172579 7717
rect 154573 7712 172579 7714
rect 154573 7656 154578 7712
rect 154634 7656 172518 7712
rect 172574 7656 172579 7712
rect 154573 7654 172579 7656
rect 154573 7651 154639 7654
rect 172513 7651 172579 7654
rect 207105 7714 207171 7717
rect 219065 7714 219131 7717
rect 246665 7714 246731 7717
rect 207105 7712 215310 7714
rect 207105 7656 207110 7712
rect 207166 7656 215310 7712
rect 207105 7654 215310 7656
rect 207105 7651 207171 7654
rect 68542 7648 68858 7649
rect 68542 7584 68548 7648
rect 68612 7584 68628 7648
rect 68692 7584 68708 7648
rect 68772 7584 68788 7648
rect 68852 7584 68858 7648
rect 68542 7583 68858 7584
rect 136139 7648 136455 7649
rect 136139 7584 136145 7648
rect 136209 7584 136225 7648
rect 136289 7584 136305 7648
rect 136369 7584 136385 7648
rect 136449 7584 136455 7648
rect 136139 7583 136455 7584
rect 203736 7648 204052 7649
rect 203736 7584 203742 7648
rect 203806 7584 203822 7648
rect 203886 7584 203902 7648
rect 203966 7584 203982 7648
rect 204046 7584 204052 7648
rect 203736 7583 204052 7584
rect 80145 7578 80211 7581
rect 94497 7578 94563 7581
rect 80145 7576 94563 7578
rect 80145 7520 80150 7576
rect 80206 7520 94502 7576
rect 94558 7520 94563 7576
rect 80145 7518 94563 7520
rect 80145 7515 80211 7518
rect 94497 7515 94563 7518
rect 138841 7578 138907 7581
rect 215250 7578 215310 7654
rect 219065 7712 246731 7714
rect 219065 7656 219070 7712
rect 219126 7656 246670 7712
rect 246726 7656 246731 7712
rect 219065 7654 246731 7656
rect 219065 7651 219131 7654
rect 246665 7651 246731 7654
rect 265341 7714 265407 7717
rect 267774 7714 267780 7716
rect 265341 7712 267780 7714
rect 265341 7656 265346 7712
rect 265402 7656 267780 7712
rect 265341 7654 267780 7656
rect 265341 7651 265407 7654
rect 267774 7652 267780 7654
rect 267844 7652 267850 7716
rect 267917 7714 267983 7717
rect 268653 7714 268719 7717
rect 271137 7714 271203 7717
rect 267917 7712 268578 7714
rect 267917 7656 267922 7712
rect 267978 7656 268578 7712
rect 267917 7654 268578 7656
rect 267917 7651 267983 7654
rect 219934 7578 219940 7580
rect 138841 7576 167010 7578
rect 138841 7520 138846 7576
rect 138902 7520 167010 7576
rect 138841 7518 167010 7520
rect 215250 7518 219940 7578
rect 138841 7515 138907 7518
rect 76557 7442 76623 7445
rect 115473 7442 115539 7445
rect 76557 7440 115539 7442
rect 76557 7384 76562 7440
rect 76618 7384 115478 7440
rect 115534 7384 115539 7440
rect 76557 7382 115539 7384
rect 76557 7379 76623 7382
rect 115473 7379 115539 7382
rect 122097 7442 122163 7445
rect 157793 7442 157859 7445
rect 122097 7440 157859 7442
rect 122097 7384 122102 7440
rect 122158 7384 157798 7440
rect 157854 7384 157859 7440
rect 122097 7382 157859 7384
rect 166950 7442 167010 7518
rect 219934 7516 219940 7518
rect 220004 7516 220010 7580
rect 220077 7578 220143 7581
rect 225965 7578 226031 7581
rect 220077 7576 226031 7578
rect 220077 7520 220082 7576
rect 220138 7520 225970 7576
rect 226026 7520 226031 7576
rect 220077 7518 226031 7520
rect 220077 7515 220143 7518
rect 225965 7515 226031 7518
rect 226149 7578 226215 7581
rect 237189 7578 237255 7581
rect 226149 7576 237255 7578
rect 226149 7520 226154 7576
rect 226210 7520 237194 7576
rect 237250 7520 237255 7576
rect 226149 7518 237255 7520
rect 226149 7515 226215 7518
rect 237189 7515 237255 7518
rect 237373 7578 237439 7581
rect 242525 7578 242591 7581
rect 237373 7576 242591 7578
rect 237373 7520 237378 7576
rect 237434 7520 242530 7576
rect 242586 7520 242591 7576
rect 237373 7518 242591 7520
rect 268518 7578 268578 7654
rect 268653 7712 271203 7714
rect 268653 7656 268658 7712
rect 268714 7656 271142 7712
rect 271198 7656 271203 7712
rect 268653 7654 271203 7656
rect 268653 7651 268719 7654
rect 271137 7651 271203 7654
rect 271781 7714 271847 7717
rect 271781 7712 272504 7714
rect 271781 7656 271786 7712
rect 271842 7656 272504 7712
rect 271781 7654 272504 7656
rect 271781 7651 271847 7654
rect 271333 7648 271649 7649
rect 271333 7584 271339 7648
rect 271403 7584 271419 7648
rect 271483 7584 271499 7648
rect 271563 7584 271579 7648
rect 271643 7584 271649 7648
rect 271333 7583 271649 7584
rect 271137 7578 271203 7581
rect 268518 7576 271203 7578
rect 268518 7520 271142 7576
rect 271198 7520 271203 7576
rect 268518 7518 271203 7520
rect 237373 7515 237439 7518
rect 242525 7515 242591 7518
rect 271137 7515 271203 7518
rect 271830 7518 272504 7578
rect 171133 7442 171199 7445
rect 166950 7440 171199 7442
rect 166950 7384 171138 7440
rect 171194 7384 171199 7440
rect 166950 7382 171199 7384
rect 122097 7379 122163 7382
rect 157793 7379 157859 7382
rect 171133 7379 171199 7382
rect 213453 7442 213519 7445
rect 252093 7442 252159 7445
rect 213453 7440 252159 7442
rect 213453 7384 213458 7440
rect 213514 7384 252098 7440
rect 252154 7384 252159 7440
rect 213453 7382 252159 7384
rect 213453 7379 213519 7382
rect 252093 7379 252159 7382
rect 261661 7442 261727 7445
rect 271830 7442 271890 7518
rect 261661 7440 271890 7442
rect 261661 7384 261666 7440
rect 261722 7384 271890 7440
rect 261661 7382 271890 7384
rect 271965 7442 272031 7445
rect 271965 7440 272504 7442
rect 271965 7384 271970 7440
rect 272026 7384 272504 7440
rect 271965 7382 272504 7384
rect 261661 7379 261727 7382
rect 271965 7379 272031 7382
rect 78765 7306 78831 7309
rect 115657 7306 115723 7309
rect 78765 7304 115723 7306
rect 78765 7248 78770 7304
rect 78826 7248 115662 7304
rect 115718 7248 115723 7304
rect 78765 7246 115723 7248
rect 78765 7243 78831 7246
rect 115657 7243 115723 7246
rect 213177 7306 213243 7309
rect 251173 7306 251239 7309
rect 213177 7304 251239 7306
rect 213177 7248 213182 7304
rect 213238 7248 251178 7304
rect 251234 7248 251239 7304
rect 213177 7246 251239 7248
rect 213177 7243 213243 7246
rect 251173 7243 251239 7246
rect 262305 7306 262371 7309
rect 262305 7304 272504 7306
rect 262305 7248 262310 7304
rect 262366 7248 272504 7304
rect 262305 7246 272504 7248
rect 262305 7243 262371 7246
rect 94497 7170 94563 7173
rect 102133 7170 102199 7173
rect 94497 7168 102199 7170
rect 94497 7112 94502 7168
rect 94558 7112 102138 7168
rect 102194 7112 102199 7168
rect 94497 7110 102199 7112
rect 94497 7107 94563 7110
rect 102133 7107 102199 7110
rect 119245 7170 119311 7173
rect 169569 7170 169635 7173
rect 119245 7168 169635 7170
rect 119245 7112 119250 7168
rect 119306 7112 169574 7168
rect 169630 7112 169635 7168
rect 119245 7110 169635 7112
rect 119245 7107 119311 7110
rect 169569 7107 169635 7110
rect 172605 7170 172671 7173
rect 220077 7170 220143 7173
rect 172605 7168 220143 7170
rect 172605 7112 172610 7168
rect 172666 7112 220082 7168
rect 220138 7112 220143 7168
rect 172605 7110 220143 7112
rect 172605 7107 172671 7110
rect 220077 7107 220143 7110
rect 222009 7170 222075 7173
rect 225781 7170 225847 7173
rect 222009 7168 225847 7170
rect 222009 7112 222014 7168
rect 222070 7112 225786 7168
rect 225842 7112 225847 7168
rect 222009 7110 225847 7112
rect 222009 7107 222075 7110
rect 225781 7107 225847 7110
rect 225965 7170 226031 7173
rect 227345 7170 227411 7173
rect 225965 7168 227411 7170
rect 225965 7112 225970 7168
rect 226026 7112 227350 7168
rect 227406 7112 227411 7168
rect 225965 7110 227411 7112
rect 225965 7107 226031 7110
rect 227345 7107 227411 7110
rect 244089 7170 244155 7173
rect 260925 7170 260991 7173
rect 244089 7168 260991 7170
rect 244089 7112 244094 7168
rect 244150 7112 260930 7168
rect 260986 7112 260991 7168
rect 244089 7110 260991 7112
rect 244089 7107 244155 7110
rect 260925 7107 260991 7110
rect 263225 7170 263291 7173
rect 263225 7168 272504 7170
rect 263225 7112 263230 7168
rect 263286 7112 272504 7168
rect 263225 7110 272504 7112
rect 263225 7107 263291 7110
rect 34744 7104 35060 7105
rect 34744 7040 34750 7104
rect 34814 7040 34830 7104
rect 34894 7040 34910 7104
rect 34974 7040 34990 7104
rect 35054 7040 35060 7104
rect 34744 7039 35060 7040
rect 102341 7104 102657 7105
rect 102341 7040 102347 7104
rect 102411 7040 102427 7104
rect 102491 7040 102507 7104
rect 102571 7040 102587 7104
rect 102651 7040 102657 7104
rect 102341 7039 102657 7040
rect 169938 7104 170254 7105
rect 169938 7040 169944 7104
rect 170008 7040 170024 7104
rect 170088 7040 170104 7104
rect 170168 7040 170184 7104
rect 170248 7040 170254 7104
rect 169938 7039 170254 7040
rect 237535 7104 237851 7105
rect 237535 7040 237541 7104
rect 237605 7040 237621 7104
rect 237685 7040 237701 7104
rect 237765 7040 237781 7104
rect 237845 7040 237851 7104
rect 237535 7039 237851 7040
rect 92473 7034 92539 7037
rect 100661 7034 100727 7037
rect 92473 7032 100727 7034
rect 92473 6976 92478 7032
rect 92534 6976 100666 7032
rect 100722 6976 100727 7032
rect 92473 6974 100727 6976
rect 92473 6971 92539 6974
rect 100661 6971 100727 6974
rect 153929 7034 153995 7037
rect 161381 7034 161447 7037
rect 153929 7032 161447 7034
rect 153929 6976 153934 7032
rect 153990 6976 161386 7032
rect 161442 6976 161447 7032
rect 153929 6974 161447 6976
rect 153929 6971 153995 6974
rect 161381 6971 161447 6974
rect 213729 7034 213795 7037
rect 219065 7034 219131 7037
rect 213729 7032 219131 7034
rect 213729 6976 213734 7032
rect 213790 6976 219070 7032
rect 219126 6976 219131 7032
rect 213729 6974 219131 6976
rect 213729 6971 213795 6974
rect 219065 6971 219131 6974
rect 223481 7034 223547 7037
rect 227437 7034 227503 7037
rect 223481 7032 227503 7034
rect 223481 6976 223486 7032
rect 223542 6976 227442 7032
rect 227498 6976 227503 7032
rect 223481 6974 227503 6976
rect 223481 6971 223547 6974
rect 227437 6971 227503 6974
rect 241513 7034 241579 7037
rect 248965 7034 249031 7037
rect 241513 7032 249031 7034
rect 241513 6976 241518 7032
rect 241574 6976 248970 7032
rect 249026 6976 249031 7032
rect 241513 6974 249031 6976
rect 241513 6971 241579 6974
rect 248965 6971 249031 6974
rect 259545 7034 259611 7037
rect 267733 7034 267799 7037
rect 259545 7032 267799 7034
rect 259545 6976 259550 7032
rect 259606 6976 267738 7032
rect 267794 6976 267799 7032
rect 259545 6974 267799 6976
rect 259545 6971 259611 6974
rect 267733 6971 267799 6974
rect 267917 7034 267983 7037
rect 267917 7032 272504 7034
rect 267917 6976 267922 7032
rect 267978 6976 272504 7032
rect 267917 6974 272504 6976
rect 267917 6971 267983 6974
rect 19241 6900 19307 6901
rect 19190 6898 19196 6900
rect 19150 6838 19196 6898
rect 19260 6896 19307 6900
rect 19302 6840 19307 6896
rect 19190 6836 19196 6838
rect 19260 6836 19307 6840
rect 19241 6835 19307 6836
rect 94221 6900 94287 6901
rect 94221 6896 94268 6900
rect 94332 6898 94338 6900
rect 97441 6898 97507 6901
rect 97901 6898 97967 6901
rect 94221 6840 94226 6896
rect 94221 6836 94268 6840
rect 94332 6838 94378 6898
rect 97441 6896 97967 6898
rect 97441 6840 97446 6896
rect 97502 6840 97906 6896
rect 97962 6840 97967 6896
rect 97441 6838 97967 6840
rect 94332 6836 94338 6838
rect 94221 6835 94287 6836
rect 97441 6835 97507 6838
rect 97901 6835 97967 6838
rect 107142 6836 107148 6900
rect 107212 6898 107218 6900
rect 112161 6898 112227 6901
rect 107212 6896 112227 6898
rect 107212 6840 112166 6896
rect 112222 6840 112227 6896
rect 107212 6838 112227 6840
rect 107212 6836 107218 6838
rect 112161 6835 112227 6838
rect 116577 6898 116643 6901
rect 119981 6898 120047 6901
rect 116577 6896 120047 6898
rect 116577 6840 116582 6896
rect 116638 6840 119986 6896
rect 120042 6840 120047 6896
rect 116577 6838 120047 6840
rect 116577 6835 116643 6838
rect 119981 6835 120047 6838
rect 218053 6898 218119 6901
rect 221825 6898 221891 6901
rect 218053 6896 221891 6898
rect 218053 6840 218058 6896
rect 218114 6840 221830 6896
rect 221886 6840 221891 6896
rect 218053 6838 221891 6840
rect 218053 6835 218119 6838
rect 221825 6835 221891 6838
rect 226701 6898 226767 6901
rect 266353 6898 266419 6901
rect 266854 6898 266860 6900
rect 226701 6896 234630 6898
rect 226701 6840 226706 6896
rect 226762 6840 234630 6896
rect 226701 6838 234630 6840
rect 226701 6835 226767 6838
rect 101765 6762 101831 6765
rect 102685 6762 102751 6765
rect 101765 6760 102751 6762
rect 101765 6704 101770 6760
rect 101826 6704 102690 6760
rect 102746 6704 102751 6760
rect 101765 6702 102751 6704
rect 101765 6699 101831 6702
rect 102685 6699 102751 6702
rect 116209 6762 116275 6765
rect 118877 6762 118943 6765
rect 142429 6762 142495 6765
rect 116209 6760 118943 6762
rect 116209 6704 116214 6760
rect 116270 6704 118882 6760
rect 118938 6704 118943 6760
rect 116209 6702 118943 6704
rect 116209 6699 116275 6702
rect 118877 6699 118943 6702
rect 128310 6760 142495 6762
rect 128310 6704 142434 6760
rect 142490 6704 142495 6760
rect 128310 6702 142495 6704
rect 82721 6626 82787 6629
rect 103605 6626 103671 6629
rect 82721 6624 103671 6626
rect 82721 6568 82726 6624
rect 82782 6568 103610 6624
rect 103666 6568 103671 6624
rect 82721 6566 103671 6568
rect 82721 6563 82787 6566
rect 103605 6563 103671 6566
rect 114553 6626 114619 6629
rect 128310 6626 128370 6702
rect 142429 6699 142495 6702
rect 152457 6762 152523 6765
rect 153837 6762 153903 6765
rect 152457 6760 153903 6762
rect 152457 6704 152462 6760
rect 152518 6704 153842 6760
rect 153898 6704 153903 6760
rect 152457 6702 153903 6704
rect 152457 6699 152523 6702
rect 153837 6699 153903 6702
rect 168281 6762 168347 6765
rect 189441 6762 189507 6765
rect 168281 6760 189507 6762
rect 168281 6704 168286 6760
rect 168342 6704 189446 6760
rect 189502 6704 189507 6760
rect 168281 6702 189507 6704
rect 168281 6699 168347 6702
rect 189441 6699 189507 6702
rect 218329 6762 218395 6765
rect 220445 6762 220511 6765
rect 218329 6760 220511 6762
rect 218329 6704 218334 6760
rect 218390 6704 220450 6760
rect 220506 6704 220511 6760
rect 218329 6702 220511 6704
rect 218329 6699 218395 6702
rect 220445 6699 220511 6702
rect 220854 6700 220860 6764
rect 220924 6762 220930 6764
rect 224861 6762 224927 6765
rect 220924 6760 224927 6762
rect 220924 6704 224866 6760
rect 224922 6704 224927 6760
rect 220924 6702 224927 6704
rect 220924 6700 220930 6702
rect 224861 6699 224927 6702
rect 227478 6700 227484 6764
rect 227548 6762 227554 6764
rect 227621 6762 227687 6765
rect 227548 6760 227687 6762
rect 227548 6704 227626 6760
rect 227682 6704 227687 6760
rect 227548 6702 227687 6704
rect 234570 6762 234630 6838
rect 266353 6896 266860 6898
rect 266353 6840 266358 6896
rect 266414 6840 266860 6896
rect 266353 6838 266860 6840
rect 266353 6835 266419 6838
rect 266854 6836 266860 6838
rect 266924 6836 266930 6900
rect 267917 6898 267983 6901
rect 267917 6896 272504 6898
rect 267917 6840 267922 6896
rect 267978 6840 272504 6896
rect 267917 6838 272504 6840
rect 267917 6835 267983 6838
rect 249006 6762 249012 6764
rect 234570 6702 249012 6762
rect 227548 6700 227554 6702
rect 227621 6699 227687 6702
rect 249006 6700 249012 6702
rect 249076 6700 249082 6764
rect 249793 6762 249859 6765
rect 258165 6762 258231 6765
rect 262673 6762 262739 6765
rect 249793 6760 258231 6762
rect 249793 6704 249798 6760
rect 249854 6704 258170 6760
rect 258226 6704 258231 6760
rect 249793 6702 258231 6704
rect 249793 6699 249859 6702
rect 258165 6699 258231 6702
rect 258766 6760 262739 6762
rect 258766 6704 262678 6760
rect 262734 6704 262739 6760
rect 258766 6702 262739 6704
rect 114553 6624 128370 6626
rect 114553 6568 114558 6624
rect 114614 6568 128370 6624
rect 114553 6566 128370 6568
rect 114553 6563 114619 6566
rect 151670 6564 151676 6628
rect 151740 6626 151746 6628
rect 170581 6626 170647 6629
rect 151740 6624 170647 6626
rect 151740 6568 170586 6624
rect 170642 6568 170647 6624
rect 151740 6566 170647 6568
rect 151740 6564 151746 6566
rect 170581 6563 170647 6566
rect 209313 6626 209379 6629
rect 218973 6626 219039 6629
rect 241605 6626 241671 6629
rect 209313 6624 219039 6626
rect 209313 6568 209318 6624
rect 209374 6568 218978 6624
rect 219034 6568 219039 6624
rect 209313 6566 219039 6568
rect 209313 6563 209379 6566
rect 218973 6563 219039 6566
rect 220126 6624 241671 6626
rect 220126 6568 241610 6624
rect 241666 6568 241671 6624
rect 220126 6566 241671 6568
rect 68542 6560 68858 6561
rect 68542 6496 68548 6560
rect 68612 6496 68628 6560
rect 68692 6496 68708 6560
rect 68772 6496 68788 6560
rect 68852 6496 68858 6560
rect 68542 6495 68858 6496
rect 136139 6560 136455 6561
rect 136139 6496 136145 6560
rect 136209 6496 136225 6560
rect 136289 6496 136305 6560
rect 136369 6496 136385 6560
rect 136449 6496 136455 6560
rect 136139 6495 136455 6496
rect 203736 6560 204052 6561
rect 203736 6496 203742 6560
rect 203806 6496 203822 6560
rect 203886 6496 203902 6560
rect 203966 6496 203982 6560
rect 204046 6496 204052 6560
rect 203736 6495 204052 6496
rect 84101 6490 84167 6493
rect 99097 6490 99163 6493
rect 84101 6488 99163 6490
rect 84101 6432 84106 6488
rect 84162 6432 99102 6488
rect 99158 6432 99163 6488
rect 84101 6430 99163 6432
rect 84101 6427 84167 6430
rect 99097 6427 99163 6430
rect 100477 6490 100543 6493
rect 115013 6490 115079 6493
rect 100477 6488 115079 6490
rect 100477 6432 100482 6488
rect 100538 6432 115018 6488
rect 115074 6432 115079 6488
rect 100477 6430 115079 6432
rect 100477 6427 100543 6430
rect 115013 6427 115079 6430
rect 144913 6490 144979 6493
rect 151997 6490 152063 6493
rect 144913 6488 152063 6490
rect 144913 6432 144918 6488
rect 144974 6432 152002 6488
rect 152058 6432 152063 6488
rect 144913 6430 152063 6432
rect 144913 6427 144979 6430
rect 151997 6427 152063 6430
rect 158161 6490 158227 6493
rect 185853 6490 185919 6493
rect 158161 6488 185919 6490
rect 158161 6432 158166 6488
rect 158222 6432 185858 6488
rect 185914 6432 185919 6488
rect 158161 6430 185919 6432
rect 158161 6427 158227 6430
rect 185853 6427 185919 6430
rect 209129 6490 209195 6493
rect 220126 6490 220186 6566
rect 241605 6563 241671 6566
rect 241789 6626 241855 6629
rect 258766 6626 258826 6702
rect 262673 6699 262739 6702
rect 265985 6762 266051 6765
rect 267641 6762 267707 6765
rect 265985 6760 267707 6762
rect 265985 6704 265990 6760
rect 266046 6704 267646 6760
rect 267702 6704 267707 6760
rect 265985 6702 267707 6704
rect 265985 6699 266051 6702
rect 267641 6699 267707 6702
rect 270953 6762 271019 6765
rect 270953 6760 272504 6762
rect 270953 6704 270958 6760
rect 271014 6704 272504 6760
rect 270953 6702 272504 6704
rect 270953 6699 271019 6702
rect 241789 6624 258826 6626
rect 241789 6568 241794 6624
rect 241850 6568 258826 6624
rect 241789 6566 258826 6568
rect 260925 6626 260991 6629
rect 269021 6626 269087 6629
rect 260925 6624 269087 6626
rect 260925 6568 260930 6624
rect 260986 6568 269026 6624
rect 269082 6568 269087 6624
rect 260925 6566 269087 6568
rect 241789 6563 241855 6566
rect 260925 6563 260991 6566
rect 269021 6563 269087 6566
rect 272057 6626 272123 6629
rect 272057 6624 272504 6626
rect 272057 6568 272062 6624
rect 272118 6568 272504 6624
rect 272057 6566 272504 6568
rect 272057 6563 272123 6566
rect 271333 6560 271649 6561
rect 271333 6496 271339 6560
rect 271403 6496 271419 6560
rect 271483 6496 271499 6560
rect 271563 6496 271579 6560
rect 271643 6496 271649 6560
rect 271333 6495 271649 6496
rect 209129 6488 220186 6490
rect 209129 6432 209134 6488
rect 209190 6432 220186 6488
rect 209129 6430 220186 6432
rect 222193 6490 222259 6493
rect 226241 6490 226307 6493
rect 222193 6488 226307 6490
rect 222193 6432 222198 6488
rect 222254 6432 226246 6488
rect 226302 6432 226307 6488
rect 222193 6430 226307 6432
rect 209129 6427 209195 6430
rect 222193 6427 222259 6430
rect 226241 6427 226307 6430
rect 229737 6490 229803 6493
rect 239397 6490 239463 6493
rect 229737 6488 239463 6490
rect 229737 6432 229742 6488
rect 229798 6432 239402 6488
rect 239458 6432 239463 6488
rect 229737 6430 239463 6432
rect 229737 6427 229803 6430
rect 239397 6427 239463 6430
rect 248321 6490 248387 6493
rect 261753 6490 261819 6493
rect 262029 6490 262095 6493
rect 248321 6488 262095 6490
rect 248321 6432 248326 6488
rect 248382 6432 261758 6488
rect 261814 6432 262034 6488
rect 262090 6432 262095 6488
rect 248321 6430 262095 6432
rect 248321 6427 248387 6430
rect 261753 6427 261819 6430
rect 262029 6427 262095 6430
rect 268101 6490 268167 6493
rect 271137 6490 271203 6493
rect 268101 6488 271203 6490
rect 268101 6432 268106 6488
rect 268162 6432 271142 6488
rect 271198 6432 271203 6488
rect 268101 6430 271203 6432
rect 268101 6427 268167 6430
rect 271137 6427 271203 6430
rect 271873 6490 271939 6493
rect 271873 6488 272504 6490
rect 271873 6432 271878 6488
rect 271934 6432 272504 6488
rect 271873 6430 272504 6432
rect 271873 6427 271939 6430
rect 78949 6354 79015 6357
rect 93894 6354 93900 6356
rect 78949 6352 93900 6354
rect 78949 6296 78954 6352
rect 79010 6296 93900 6352
rect 78949 6294 93900 6296
rect 78949 6291 79015 6294
rect 93894 6292 93900 6294
rect 93964 6292 93970 6356
rect 94497 6354 94563 6357
rect 109585 6354 109651 6357
rect 94497 6352 109651 6354
rect 94497 6296 94502 6352
rect 94558 6296 109590 6352
rect 109646 6296 109651 6352
rect 94497 6294 109651 6296
rect 94497 6291 94563 6294
rect 109585 6291 109651 6294
rect 113449 6354 113515 6357
rect 114737 6354 114803 6357
rect 113449 6352 114803 6354
rect 113449 6296 113454 6352
rect 113510 6296 114742 6352
rect 114798 6296 114803 6352
rect 113449 6294 114803 6296
rect 113449 6291 113515 6294
rect 114737 6291 114803 6294
rect 117865 6354 117931 6357
rect 139761 6354 139827 6357
rect 117865 6352 139827 6354
rect 117865 6296 117870 6352
rect 117926 6296 139766 6352
rect 139822 6296 139827 6352
rect 117865 6294 139827 6296
rect 117865 6291 117931 6294
rect 139761 6291 139827 6294
rect 146293 6354 146359 6357
rect 169753 6354 169819 6357
rect 146293 6352 169819 6354
rect 146293 6296 146298 6352
rect 146354 6296 169758 6352
rect 169814 6296 169819 6352
rect 146293 6294 169819 6296
rect 146293 6291 146359 6294
rect 169753 6291 169819 6294
rect 213085 6354 213151 6357
rect 251633 6354 251699 6357
rect 213085 6352 251699 6354
rect 213085 6296 213090 6352
rect 213146 6296 251638 6352
rect 251694 6296 251699 6352
rect 213085 6294 251699 6296
rect 213085 6291 213151 6294
rect 251633 6291 251699 6294
rect 268745 6354 268811 6357
rect 270677 6354 270743 6357
rect 271086 6354 271092 6356
rect 268745 6352 270602 6354
rect 268745 6296 268750 6352
rect 268806 6296 270602 6352
rect 268745 6294 270602 6296
rect 268745 6291 268811 6294
rect 53741 6218 53807 6221
rect 100201 6218 100267 6221
rect 53741 6216 100267 6218
rect 53741 6160 53746 6216
rect 53802 6160 100206 6216
rect 100262 6160 100267 6216
rect 53741 6158 100267 6160
rect 53741 6155 53807 6158
rect 100201 6155 100267 6158
rect 101305 6218 101371 6221
rect 108205 6218 108271 6221
rect 101305 6216 108271 6218
rect 101305 6160 101310 6216
rect 101366 6160 108210 6216
rect 108266 6160 108271 6216
rect 101305 6158 108271 6160
rect 101305 6155 101371 6158
rect 108205 6155 108271 6158
rect 112897 6218 112963 6221
rect 114829 6218 114895 6221
rect 112897 6216 114895 6218
rect 112897 6160 112902 6216
rect 112958 6160 114834 6216
rect 114890 6160 114895 6216
rect 112897 6158 114895 6160
rect 112897 6155 112963 6158
rect 114829 6155 114895 6158
rect 118141 6218 118207 6221
rect 127709 6218 127775 6221
rect 168833 6218 168899 6221
rect 118141 6216 168899 6218
rect 118141 6160 118146 6216
rect 118202 6160 127714 6216
rect 127770 6160 168838 6216
rect 168894 6160 168899 6216
rect 118141 6158 168899 6160
rect 118141 6155 118207 6158
rect 127709 6155 127775 6158
rect 168833 6155 168899 6158
rect 189993 6218 190059 6221
rect 216397 6218 216463 6221
rect 189993 6216 216463 6218
rect 189993 6160 189998 6216
rect 190054 6160 216402 6216
rect 216458 6160 216463 6216
rect 189993 6158 216463 6160
rect 189993 6155 190059 6158
rect 216397 6155 216463 6158
rect 219893 6218 219959 6221
rect 229737 6218 229803 6221
rect 239397 6218 239463 6221
rect 253473 6218 253539 6221
rect 219893 6216 229803 6218
rect 219893 6160 219898 6216
rect 219954 6160 229742 6216
rect 229798 6160 229803 6216
rect 219893 6158 229803 6160
rect 219893 6155 219959 6158
rect 229737 6155 229803 6158
rect 234570 6158 238034 6218
rect 95049 6082 95115 6085
rect 101949 6082 102015 6085
rect 95049 6080 102015 6082
rect 95049 6024 95054 6080
rect 95110 6024 101954 6080
rect 102010 6024 102015 6080
rect 95049 6022 102015 6024
rect 95049 6019 95115 6022
rect 101949 6019 102015 6022
rect 115933 6082 115999 6085
rect 116485 6082 116551 6085
rect 115933 6080 116551 6082
rect 115933 6024 115938 6080
rect 115994 6024 116490 6080
rect 116546 6024 116551 6080
rect 115933 6022 116551 6024
rect 115933 6019 115999 6022
rect 116485 6019 116551 6022
rect 121913 6082 121979 6085
rect 148501 6082 148567 6085
rect 121913 6080 148567 6082
rect 121913 6024 121918 6080
rect 121974 6024 148506 6080
rect 148562 6024 148567 6080
rect 121913 6022 148567 6024
rect 121913 6019 121979 6022
rect 148501 6019 148567 6022
rect 170765 6082 170831 6085
rect 216581 6082 216647 6085
rect 170765 6080 216647 6082
rect 170765 6024 170770 6080
rect 170826 6024 216586 6080
rect 216642 6024 216647 6080
rect 170765 6022 216647 6024
rect 170765 6019 170831 6022
rect 216581 6019 216647 6022
rect 219433 6082 219499 6085
rect 234570 6082 234630 6158
rect 219433 6080 234630 6082
rect 219433 6024 219438 6080
rect 219494 6024 234630 6080
rect 219433 6022 234630 6024
rect 237974 6082 238034 6158
rect 239397 6216 253539 6218
rect 239397 6160 239402 6216
rect 239458 6160 253478 6216
rect 253534 6160 253539 6216
rect 239397 6158 253539 6160
rect 239397 6155 239463 6158
rect 253473 6155 253539 6158
rect 268510 6156 268516 6220
rect 268580 6218 268586 6220
rect 268929 6218 268995 6221
rect 268580 6216 268995 6218
rect 268580 6160 268934 6216
rect 268990 6160 268995 6216
rect 268580 6158 268995 6160
rect 268580 6156 268586 6158
rect 268929 6155 268995 6158
rect 269982 6156 269988 6220
rect 270052 6218 270058 6220
rect 270309 6218 270375 6221
rect 270052 6216 270375 6218
rect 270052 6160 270314 6216
rect 270370 6160 270375 6216
rect 270052 6158 270375 6160
rect 270542 6218 270602 6294
rect 270677 6352 271092 6354
rect 270677 6296 270682 6352
rect 270738 6296 271092 6352
rect 270677 6294 271092 6296
rect 270677 6291 270743 6294
rect 271086 6292 271092 6294
rect 271156 6292 271162 6356
rect 271321 6354 271387 6357
rect 271321 6352 272504 6354
rect 271321 6296 271326 6352
rect 271382 6296 272504 6352
rect 271321 6294 272504 6296
rect 271321 6291 271387 6294
rect 270542 6158 272504 6218
rect 270052 6156 270058 6158
rect 270309 6155 270375 6158
rect 258257 6082 258323 6085
rect 237974 6080 258323 6082
rect 237974 6024 258262 6080
rect 258318 6024 258323 6080
rect 237974 6022 258323 6024
rect 219433 6019 219499 6022
rect 258257 6019 258323 6022
rect 260833 6082 260899 6085
rect 268469 6082 268535 6085
rect 260833 6080 268535 6082
rect 260833 6024 260838 6080
rect 260894 6024 268474 6080
rect 268530 6024 268535 6080
rect 260833 6022 268535 6024
rect 260833 6019 260899 6022
rect 268469 6019 268535 6022
rect 268837 6082 268903 6085
rect 271321 6082 271387 6085
rect 268837 6080 271387 6082
rect 268837 6024 268842 6080
rect 268898 6024 271326 6080
rect 271382 6024 271387 6080
rect 268837 6022 271387 6024
rect 268837 6019 268903 6022
rect 271321 6019 271387 6022
rect 271689 6082 271755 6085
rect 271689 6080 272504 6082
rect 271689 6024 271694 6080
rect 271750 6024 272504 6080
rect 271689 6022 272504 6024
rect 271689 6019 271755 6022
rect 34744 6016 35060 6017
rect 34744 5952 34750 6016
rect 34814 5952 34830 6016
rect 34894 5952 34910 6016
rect 34974 5952 34990 6016
rect 35054 5952 35060 6016
rect 34744 5951 35060 5952
rect 102341 6016 102657 6017
rect 102341 5952 102347 6016
rect 102411 5952 102427 6016
rect 102491 5952 102507 6016
rect 102571 5952 102587 6016
rect 102651 5952 102657 6016
rect 102341 5951 102657 5952
rect 169938 6016 170254 6017
rect 169938 5952 169944 6016
rect 170008 5952 170024 6016
rect 170088 5952 170104 6016
rect 170168 5952 170184 6016
rect 170248 5952 170254 6016
rect 169938 5951 170254 5952
rect 237535 6016 237851 6017
rect 237535 5952 237541 6016
rect 237605 5952 237621 6016
rect 237685 5952 237701 6016
rect 237765 5952 237781 6016
rect 237845 5952 237851 6016
rect 237535 5951 237851 5952
rect 42793 5946 42859 5949
rect 100845 5946 100911 5949
rect 42793 5944 100911 5946
rect 42793 5888 42798 5944
rect 42854 5888 100850 5944
rect 100906 5888 100911 5944
rect 42793 5886 100911 5888
rect 42793 5883 42859 5886
rect 100845 5883 100911 5886
rect 101489 5946 101555 5949
rect 102041 5946 102107 5949
rect 101489 5944 102107 5946
rect 101489 5888 101494 5944
rect 101550 5888 102046 5944
rect 102102 5888 102107 5944
rect 101489 5886 102107 5888
rect 101489 5883 101555 5886
rect 102041 5883 102107 5886
rect 105997 5946 106063 5949
rect 116485 5946 116551 5949
rect 117865 5946 117931 5949
rect 105997 5944 117931 5946
rect 105997 5888 106002 5944
rect 106058 5888 116490 5944
rect 116546 5888 117870 5944
rect 117926 5888 117931 5944
rect 105997 5886 117931 5888
rect 105997 5883 106063 5886
rect 116485 5883 116551 5886
rect 117865 5883 117931 5886
rect 139761 5946 139827 5949
rect 219249 5946 219315 5949
rect 224585 5946 224651 5949
rect 227897 5946 227963 5949
rect 139761 5944 169218 5946
rect 139761 5888 139766 5944
rect 139822 5888 169218 5944
rect 139761 5886 169218 5888
rect 139761 5883 139827 5886
rect 169158 5813 169218 5886
rect 219249 5944 227963 5946
rect 219249 5888 219254 5944
rect 219310 5888 224590 5944
rect 224646 5888 227902 5944
rect 227958 5888 227963 5944
rect 219249 5886 227963 5888
rect 219249 5883 219315 5886
rect 224585 5883 224651 5886
rect 227897 5883 227963 5886
rect 264789 5946 264855 5949
rect 268653 5946 268719 5949
rect 264789 5944 268719 5946
rect 264789 5888 264794 5944
rect 264850 5888 268658 5944
rect 268714 5888 268719 5944
rect 264789 5886 268719 5888
rect 264789 5883 264855 5886
rect 268653 5883 268719 5886
rect 269021 5946 269087 5949
rect 271137 5946 271203 5949
rect 269021 5944 270970 5946
rect 269021 5888 269026 5944
rect 269082 5888 270970 5944
rect 269021 5886 270970 5888
rect 269021 5883 269087 5886
rect 94497 5810 94563 5813
rect 109033 5810 109099 5813
rect 94497 5808 109099 5810
rect 94497 5752 94502 5808
rect 94558 5752 109038 5808
rect 109094 5752 109099 5808
rect 94497 5750 109099 5752
rect 94497 5747 94563 5750
rect 109033 5747 109099 5750
rect 113081 5810 113147 5813
rect 116393 5810 116459 5813
rect 113081 5808 116459 5810
rect 113081 5752 113086 5808
rect 113142 5752 116398 5808
rect 116454 5752 116459 5808
rect 113081 5750 116459 5752
rect 113081 5747 113147 5750
rect 116393 5747 116459 5750
rect 137277 5810 137343 5813
rect 168281 5810 168347 5813
rect 137277 5808 168347 5810
rect 137277 5752 137282 5808
rect 137338 5752 168286 5808
rect 168342 5752 168347 5808
rect 137277 5750 168347 5752
rect 169158 5810 169267 5813
rect 212809 5810 212875 5813
rect 169158 5808 212875 5810
rect 169158 5752 169206 5808
rect 169262 5752 212814 5808
rect 212870 5752 212875 5808
rect 169158 5750 212875 5752
rect 137277 5747 137343 5750
rect 168281 5747 168347 5750
rect 169201 5747 169267 5750
rect 212809 5747 212875 5750
rect 213862 5748 213868 5812
rect 213932 5810 213938 5812
rect 216581 5810 216647 5813
rect 226241 5810 226307 5813
rect 258257 5810 258323 5813
rect 266353 5812 266419 5813
rect 213932 5808 216647 5810
rect 213932 5752 216586 5808
rect 216642 5752 216647 5808
rect 213932 5750 216647 5752
rect 213932 5748 213938 5750
rect 216581 5747 216647 5750
rect 216814 5750 224970 5810
rect 53281 5674 53347 5677
rect 100293 5674 100359 5677
rect 101305 5674 101371 5677
rect 53281 5672 95434 5674
rect 53281 5616 53286 5672
rect 53342 5616 95434 5672
rect 53281 5614 95434 5616
rect 53281 5611 53347 5614
rect 94405 5538 94471 5541
rect 95182 5538 95188 5540
rect 94405 5536 95188 5538
rect 94405 5480 94410 5536
rect 94466 5480 95188 5536
rect 94405 5478 95188 5480
rect 94405 5475 94471 5478
rect 95182 5476 95188 5478
rect 95252 5476 95258 5540
rect 68542 5472 68858 5473
rect 68542 5408 68548 5472
rect 68612 5408 68628 5472
rect 68692 5408 68708 5472
rect 68772 5408 68788 5472
rect 68852 5408 68858 5472
rect 68542 5407 68858 5408
rect 19333 5266 19399 5269
rect 36261 5266 36327 5269
rect 19333 5264 36327 5266
rect 19333 5208 19338 5264
rect 19394 5208 36266 5264
rect 36322 5208 36327 5264
rect 19333 5206 36327 5208
rect 95374 5266 95434 5614
rect 100293 5672 101371 5674
rect 100293 5616 100298 5672
rect 100354 5616 101310 5672
rect 101366 5616 101371 5672
rect 100293 5614 101371 5616
rect 100293 5611 100359 5614
rect 101305 5611 101371 5614
rect 101673 5674 101739 5677
rect 121913 5674 121979 5677
rect 101673 5672 121979 5674
rect 101673 5616 101678 5672
rect 101734 5616 121918 5672
rect 121974 5616 121979 5672
rect 101673 5614 121979 5616
rect 101673 5611 101739 5614
rect 121913 5611 121979 5614
rect 136081 5674 136147 5677
rect 140681 5674 140747 5677
rect 136081 5672 140747 5674
rect 136081 5616 136086 5672
rect 136142 5616 140686 5672
rect 140742 5616 140747 5672
rect 136081 5614 140747 5616
rect 136081 5611 136147 5614
rect 140681 5611 140747 5614
rect 144821 5674 144887 5677
rect 151854 5674 151860 5676
rect 144821 5672 151860 5674
rect 144821 5616 144826 5672
rect 144882 5616 151860 5672
rect 144821 5614 151860 5616
rect 144821 5611 144887 5614
rect 151854 5612 151860 5614
rect 151924 5612 151930 5676
rect 152089 5674 152155 5677
rect 172513 5674 172579 5677
rect 152089 5672 172579 5674
rect 152089 5616 152094 5672
rect 152150 5616 172518 5672
rect 172574 5616 172579 5672
rect 152089 5614 172579 5616
rect 152089 5611 152155 5614
rect 172513 5611 172579 5614
rect 216397 5674 216463 5677
rect 216814 5674 216874 5750
rect 216397 5672 216874 5674
rect 216397 5616 216402 5672
rect 216458 5616 216874 5672
rect 216397 5614 216874 5616
rect 219985 5674 220051 5677
rect 223573 5674 223639 5677
rect 219985 5672 223639 5674
rect 219985 5616 219990 5672
rect 220046 5616 223578 5672
rect 223634 5616 223639 5672
rect 219985 5614 223639 5616
rect 224910 5674 224970 5750
rect 226241 5808 258323 5810
rect 226241 5752 226246 5808
rect 226302 5752 258262 5808
rect 258318 5752 258323 5808
rect 226241 5750 258323 5752
rect 226241 5747 226307 5750
rect 258257 5747 258323 5750
rect 266302 5748 266308 5812
rect 266372 5810 266419 5812
rect 268285 5810 268351 5813
rect 270910 5810 270970 5886
rect 271137 5944 272504 5946
rect 271137 5888 271142 5944
rect 271198 5888 272504 5944
rect 271137 5886 272504 5888
rect 271137 5883 271203 5886
rect 266372 5808 266464 5810
rect 266414 5752 266464 5808
rect 266372 5750 266464 5752
rect 268285 5808 270786 5810
rect 268285 5752 268290 5808
rect 268346 5752 270786 5808
rect 268285 5750 270786 5752
rect 270910 5750 272504 5810
rect 266372 5748 266419 5750
rect 266353 5747 266419 5748
rect 268285 5747 268351 5750
rect 247401 5674 247467 5677
rect 224910 5672 247467 5674
rect 224910 5616 247406 5672
rect 247462 5616 247467 5672
rect 224910 5614 247467 5616
rect 216397 5611 216463 5614
rect 219985 5611 220051 5614
rect 223573 5611 223639 5614
rect 247401 5611 247467 5614
rect 263409 5674 263475 5677
rect 268469 5674 268535 5677
rect 263409 5672 268535 5674
rect 263409 5616 263414 5672
rect 263470 5616 268474 5672
rect 268530 5616 268535 5672
rect 263409 5614 268535 5616
rect 263409 5611 263475 5614
rect 268469 5611 268535 5614
rect 269246 5612 269252 5676
rect 269316 5674 269322 5676
rect 269481 5674 269547 5677
rect 270493 5676 270559 5677
rect 270493 5674 270540 5676
rect 269316 5672 269547 5674
rect 269316 5616 269486 5672
rect 269542 5616 269547 5672
rect 269316 5614 269547 5616
rect 270448 5672 270540 5674
rect 270448 5616 270498 5672
rect 270448 5614 270540 5616
rect 269316 5612 269322 5614
rect 269481 5611 269547 5614
rect 270493 5612 270540 5614
rect 270604 5612 270610 5676
rect 270726 5674 270786 5750
rect 270726 5614 272504 5674
rect 270493 5611 270559 5612
rect 96061 5538 96127 5541
rect 111425 5538 111491 5541
rect 114461 5538 114527 5541
rect 96061 5536 96170 5538
rect 96061 5480 96066 5536
rect 96122 5480 96170 5536
rect 96061 5475 96170 5480
rect 111425 5536 114527 5538
rect 111425 5480 111430 5536
rect 111486 5480 114466 5536
rect 114522 5480 114527 5536
rect 111425 5478 114527 5480
rect 111425 5475 111491 5478
rect 114461 5475 114527 5478
rect 150065 5538 150131 5541
rect 153561 5538 153627 5541
rect 150065 5536 153627 5538
rect 150065 5480 150070 5536
rect 150126 5480 153566 5536
rect 153622 5480 153627 5536
rect 150065 5478 153627 5480
rect 150065 5475 150131 5478
rect 153561 5475 153627 5478
rect 206185 5538 206251 5541
rect 209129 5538 209195 5541
rect 206185 5536 209195 5538
rect 206185 5480 206190 5536
rect 206246 5480 209134 5536
rect 209190 5480 209195 5536
rect 206185 5478 209195 5480
rect 206185 5475 206251 5478
rect 209129 5475 209195 5478
rect 213177 5538 213243 5541
rect 214465 5538 214531 5541
rect 220854 5538 220860 5540
rect 213177 5536 220860 5538
rect 213177 5480 213182 5536
rect 213238 5480 214470 5536
rect 214526 5480 220860 5536
rect 213177 5478 220860 5480
rect 213177 5475 213243 5478
rect 214465 5475 214531 5478
rect 220854 5476 220860 5478
rect 220924 5476 220930 5540
rect 229001 5538 229067 5541
rect 250345 5538 250411 5541
rect 229001 5536 250411 5538
rect 229001 5480 229006 5536
rect 229062 5480 250350 5536
rect 250406 5480 250411 5536
rect 229001 5478 250411 5480
rect 229001 5475 229067 5478
rect 250345 5475 250411 5478
rect 254301 5538 254367 5541
rect 267641 5538 267707 5541
rect 254301 5536 267707 5538
rect 254301 5480 254306 5536
rect 254362 5480 267646 5536
rect 267702 5480 267707 5536
rect 254301 5478 267707 5480
rect 254301 5475 254367 5478
rect 267641 5475 267707 5478
rect 268653 5538 268719 5541
rect 271137 5538 271203 5541
rect 268653 5536 271203 5538
rect 268653 5480 268658 5536
rect 268714 5480 271142 5536
rect 271198 5480 271203 5536
rect 268653 5478 271203 5480
rect 268653 5475 268719 5478
rect 271137 5475 271203 5478
rect 271781 5538 271847 5541
rect 271781 5536 272504 5538
rect 271781 5480 271786 5536
rect 271842 5480 272504 5536
rect 271781 5478 272504 5480
rect 271781 5475 271847 5478
rect 96110 5402 96170 5475
rect 136139 5472 136455 5473
rect 136139 5408 136145 5472
rect 136209 5408 136225 5472
rect 136289 5408 136305 5472
rect 136369 5408 136385 5472
rect 136449 5408 136455 5472
rect 136139 5407 136455 5408
rect 203736 5472 204052 5473
rect 203736 5408 203742 5472
rect 203806 5408 203822 5472
rect 203886 5408 203902 5472
rect 203966 5408 203982 5472
rect 204046 5408 204052 5472
rect 203736 5407 204052 5408
rect 271333 5472 271649 5473
rect 271333 5408 271339 5472
rect 271403 5408 271419 5472
rect 271483 5408 271499 5472
rect 271563 5408 271579 5472
rect 271643 5408 271649 5472
rect 271333 5407 271649 5408
rect 97533 5402 97599 5405
rect 96110 5400 97599 5402
rect 96110 5344 97538 5400
rect 97594 5344 97599 5400
rect 96110 5342 97599 5344
rect 97533 5339 97599 5342
rect 98453 5402 98519 5405
rect 113030 5402 113036 5404
rect 98453 5400 113036 5402
rect 98453 5344 98458 5400
rect 98514 5344 113036 5400
rect 98453 5342 113036 5344
rect 98453 5339 98519 5342
rect 113030 5340 113036 5342
rect 113100 5340 113106 5404
rect 113541 5402 113607 5405
rect 114553 5402 114619 5405
rect 113541 5400 114619 5402
rect 113541 5344 113546 5400
rect 113602 5344 114558 5400
rect 114614 5344 114619 5400
rect 113541 5342 114619 5344
rect 113541 5339 113607 5342
rect 114553 5339 114619 5342
rect 151721 5402 151787 5405
rect 175273 5402 175339 5405
rect 151721 5400 175339 5402
rect 151721 5344 151726 5400
rect 151782 5344 175278 5400
rect 175334 5344 175339 5400
rect 151721 5342 175339 5344
rect 151721 5339 151787 5342
rect 175273 5339 175339 5342
rect 214373 5402 214439 5405
rect 242893 5402 242959 5405
rect 214373 5400 242959 5402
rect 214373 5344 214378 5400
rect 214434 5344 242898 5400
rect 242954 5344 242959 5400
rect 214373 5342 242959 5344
rect 214373 5339 214439 5342
rect 242893 5339 242959 5342
rect 249006 5340 249012 5404
rect 249076 5402 249082 5404
rect 255129 5402 255195 5405
rect 249076 5400 255195 5402
rect 249076 5344 255134 5400
rect 255190 5344 255195 5400
rect 249076 5342 255195 5344
rect 249076 5340 249082 5342
rect 255129 5339 255195 5342
rect 271781 5402 271847 5405
rect 271781 5400 272504 5402
rect 271781 5344 271786 5400
rect 271842 5344 272504 5400
rect 271781 5342 272504 5344
rect 271781 5339 271847 5342
rect 110781 5266 110847 5269
rect 95374 5264 110847 5266
rect 95374 5208 110786 5264
rect 110842 5208 110847 5264
rect 95374 5206 110847 5208
rect 19333 5203 19399 5206
rect 36261 5203 36327 5206
rect 110781 5203 110847 5206
rect 111425 5266 111491 5269
rect 115013 5266 115079 5269
rect 111425 5264 115079 5266
rect 111425 5208 111430 5264
rect 111486 5208 115018 5264
rect 115074 5208 115079 5264
rect 111425 5206 115079 5208
rect 111425 5203 111491 5206
rect 115013 5203 115079 5206
rect 116025 5266 116091 5269
rect 117589 5266 117655 5269
rect 116025 5264 117655 5266
rect 116025 5208 116030 5264
rect 116086 5208 117594 5264
rect 117650 5208 117655 5264
rect 116025 5206 117655 5208
rect 116025 5203 116091 5206
rect 117589 5203 117655 5206
rect 149973 5266 150039 5269
rect 150249 5266 150315 5269
rect 149973 5264 150315 5266
rect 149973 5208 149978 5264
rect 150034 5208 150254 5264
rect 150310 5208 150315 5264
rect 149973 5206 150315 5208
rect 149973 5203 150039 5206
rect 150249 5203 150315 5206
rect 154757 5266 154823 5269
rect 219433 5266 219499 5269
rect 154757 5264 219499 5266
rect 154757 5208 154762 5264
rect 154818 5208 219438 5264
rect 219494 5208 219499 5264
rect 154757 5206 219499 5208
rect 154757 5203 154823 5206
rect 219433 5203 219499 5206
rect 219934 5204 219940 5268
rect 220004 5266 220010 5268
rect 223757 5266 223823 5269
rect 237281 5266 237347 5269
rect 220004 5264 223823 5266
rect 220004 5208 223762 5264
rect 223818 5208 223823 5264
rect 220004 5206 223823 5208
rect 220004 5204 220010 5206
rect 223757 5203 223823 5206
rect 224910 5264 237347 5266
rect 224910 5208 237286 5264
rect 237342 5208 237347 5264
rect 224910 5206 237347 5208
rect 42609 5130 42675 5133
rect 46657 5130 46723 5133
rect 42609 5128 46723 5130
rect 42609 5072 42614 5128
rect 42670 5072 46662 5128
rect 46718 5072 46723 5128
rect 42609 5070 46723 5072
rect 42609 5067 42675 5070
rect 46657 5067 46723 5070
rect 47117 5130 47183 5133
rect 109125 5130 109191 5133
rect 47117 5128 109191 5130
rect 47117 5072 47122 5128
rect 47178 5072 109130 5128
rect 109186 5072 109191 5128
rect 47117 5070 109191 5072
rect 47117 5067 47183 5070
rect 109125 5067 109191 5070
rect 113081 5130 113147 5133
rect 114645 5130 114711 5133
rect 151721 5130 151787 5133
rect 113081 5128 114711 5130
rect 113081 5072 113086 5128
rect 113142 5072 114650 5128
rect 114706 5072 114711 5128
rect 113081 5070 114711 5072
rect 113081 5067 113147 5070
rect 114645 5067 114711 5070
rect 118650 5128 151787 5130
rect 118650 5072 151726 5128
rect 151782 5072 151787 5128
rect 118650 5070 151787 5072
rect 36813 4994 36879 4997
rect 96613 4994 96679 4997
rect 36813 4992 96679 4994
rect 36813 4936 36818 4992
rect 36874 4936 96618 4992
rect 96674 4936 96679 4992
rect 36813 4934 96679 4936
rect 36813 4931 36879 4934
rect 96613 4931 96679 4934
rect 104341 4994 104407 4997
rect 105997 4994 106063 4997
rect 104341 4992 106063 4994
rect 104341 4936 104346 4992
rect 104402 4936 106002 4992
rect 106058 4936 106063 4992
rect 104341 4934 106063 4936
rect 104341 4931 104407 4934
rect 105997 4931 106063 4934
rect 108665 4994 108731 4997
rect 118650 4994 118710 5070
rect 151721 5067 151787 5070
rect 151905 5130 151971 5133
rect 153101 5130 153167 5133
rect 151905 5128 153167 5130
rect 151905 5072 151910 5128
rect 151966 5072 153106 5128
rect 153162 5072 153167 5128
rect 151905 5070 153167 5072
rect 151905 5067 151971 5070
rect 153101 5067 153167 5070
rect 208393 5130 208459 5133
rect 224910 5130 224970 5206
rect 237281 5203 237347 5206
rect 246205 5266 246271 5269
rect 248321 5266 248387 5269
rect 246205 5264 248387 5266
rect 246205 5208 246210 5264
rect 246266 5208 248326 5264
rect 248382 5208 248387 5264
rect 246205 5206 248387 5208
rect 246205 5203 246271 5206
rect 248321 5203 248387 5206
rect 261017 5266 261083 5269
rect 266905 5266 266971 5269
rect 261017 5264 266971 5266
rect 261017 5208 261022 5264
rect 261078 5208 266910 5264
rect 266966 5208 266971 5264
rect 261017 5206 266971 5208
rect 261017 5203 261083 5206
rect 266905 5203 266971 5206
rect 269021 5266 269087 5269
rect 269021 5264 272504 5266
rect 269021 5208 269026 5264
rect 269082 5208 272504 5264
rect 269021 5206 272504 5208
rect 269021 5203 269087 5206
rect 246297 5130 246363 5133
rect 208393 5128 224970 5130
rect 208393 5072 208398 5128
rect 208454 5072 224970 5128
rect 208393 5070 224970 5072
rect 234570 5128 246363 5130
rect 234570 5072 246302 5128
rect 246358 5072 246363 5128
rect 234570 5070 246363 5072
rect 208393 5067 208459 5070
rect 108665 4992 118710 4994
rect 108665 4936 108670 4992
rect 108726 4936 118710 4992
rect 108665 4934 118710 4936
rect 141509 4994 141575 4997
rect 152917 4994 152983 4997
rect 141509 4992 152983 4994
rect 141509 4936 141514 4992
rect 141570 4936 152922 4992
rect 152978 4936 152983 4992
rect 141509 4934 152983 4936
rect 108665 4931 108731 4934
rect 141509 4931 141575 4934
rect 152917 4931 152983 4934
rect 215845 4994 215911 4997
rect 234570 4994 234630 5070
rect 246297 5067 246363 5070
rect 268469 5130 268535 5133
rect 268469 5128 272504 5130
rect 268469 5072 268474 5128
rect 268530 5072 272504 5128
rect 268469 5070 272504 5072
rect 268469 5067 268535 5070
rect 215845 4992 234630 4994
rect 215845 4936 215850 4992
rect 215906 4936 234630 4992
rect 215845 4934 234630 4936
rect 267733 4994 267799 4997
rect 271781 4994 271847 4997
rect 267733 4992 271847 4994
rect 267733 4936 267738 4992
rect 267794 4936 271786 4992
rect 271842 4936 271847 4992
rect 267733 4934 271847 4936
rect 215845 4931 215911 4934
rect 267733 4931 267799 4934
rect 271781 4931 271847 4934
rect 271965 4994 272031 4997
rect 271965 4992 272504 4994
rect 271965 4936 271970 4992
rect 272026 4936 272504 4992
rect 271965 4934 272504 4936
rect 271965 4931 272031 4934
rect 34744 4928 35060 4929
rect 34744 4864 34750 4928
rect 34814 4864 34830 4928
rect 34894 4864 34910 4928
rect 34974 4864 34990 4928
rect 35054 4864 35060 4928
rect 34744 4863 35060 4864
rect 102341 4928 102657 4929
rect 102341 4864 102347 4928
rect 102411 4864 102427 4928
rect 102491 4864 102507 4928
rect 102571 4864 102587 4928
rect 102651 4864 102657 4928
rect 102341 4863 102657 4864
rect 169938 4928 170254 4929
rect 169938 4864 169944 4928
rect 170008 4864 170024 4928
rect 170088 4864 170104 4928
rect 170168 4864 170184 4928
rect 170248 4864 170254 4928
rect 169938 4863 170254 4864
rect 237535 4928 237851 4929
rect 237535 4864 237541 4928
rect 237605 4864 237621 4928
rect 237685 4864 237701 4928
rect 237765 4864 237781 4928
rect 237845 4864 237851 4928
rect 237535 4863 237851 4864
rect 99465 4858 99531 4861
rect 100017 4858 100083 4861
rect 99465 4856 100083 4858
rect 99465 4800 99470 4856
rect 99526 4800 100022 4856
rect 100078 4800 100083 4856
rect 99465 4798 100083 4800
rect 99465 4795 99531 4798
rect 100017 4795 100083 4798
rect 106038 4796 106044 4860
rect 106108 4858 106114 4860
rect 106181 4858 106247 4861
rect 106108 4856 106247 4858
rect 106108 4800 106186 4856
rect 106242 4800 106247 4856
rect 106108 4798 106247 4800
rect 106108 4796 106114 4798
rect 106181 4795 106247 4798
rect 110270 4796 110276 4860
rect 110340 4858 110346 4860
rect 149973 4858 150039 4861
rect 110340 4856 150039 4858
rect 110340 4800 149978 4856
rect 150034 4800 150039 4856
rect 110340 4798 150039 4800
rect 110340 4796 110346 4798
rect 149973 4795 150039 4798
rect 150157 4858 150223 4861
rect 158529 4858 158595 4861
rect 150157 4856 158595 4858
rect 150157 4800 150162 4856
rect 150218 4800 158534 4856
rect 158590 4800 158595 4856
rect 150157 4798 158595 4800
rect 150157 4795 150223 4798
rect 158529 4795 158595 4798
rect 214373 4858 214439 4861
rect 220537 4858 220603 4861
rect 214373 4856 220603 4858
rect 214373 4800 214378 4856
rect 214434 4800 220542 4856
rect 220598 4800 220603 4856
rect 214373 4798 220603 4800
rect 214373 4795 214439 4798
rect 220537 4795 220603 4798
rect 223665 4858 223731 4861
rect 225086 4858 225092 4860
rect 223665 4856 225092 4858
rect 223665 4800 223670 4856
rect 223726 4800 225092 4856
rect 223665 4798 225092 4800
rect 223665 4795 223731 4798
rect 225086 4796 225092 4798
rect 225156 4796 225162 4860
rect 251081 4858 251147 4861
rect 263225 4858 263291 4861
rect 251081 4856 263291 4858
rect 251081 4800 251086 4856
rect 251142 4800 263230 4856
rect 263286 4800 263291 4856
rect 251081 4798 263291 4800
rect 251081 4795 251147 4798
rect 263225 4795 263291 4798
rect 268929 4858 268995 4861
rect 268929 4856 272504 4858
rect 268929 4800 268934 4856
rect 268990 4800 272504 4856
rect 268929 4798 272504 4800
rect 268929 4795 268995 4798
rect 100661 4722 100727 4725
rect 114921 4722 114987 4725
rect 100661 4720 114987 4722
rect 100661 4664 100666 4720
rect 100722 4664 114926 4720
rect 114982 4664 114987 4720
rect 100661 4662 114987 4664
rect 100661 4659 100727 4662
rect 114921 4659 114987 4662
rect 116025 4722 116091 4725
rect 121361 4722 121427 4725
rect 116025 4720 121427 4722
rect 116025 4664 116030 4720
rect 116086 4664 121366 4720
rect 121422 4664 121427 4720
rect 116025 4662 121427 4664
rect 116025 4659 116091 4662
rect 121361 4659 121427 4662
rect 149881 4722 149947 4725
rect 178401 4722 178467 4725
rect 149881 4720 178467 4722
rect 149881 4664 149886 4720
rect 149942 4664 178406 4720
rect 178462 4664 178467 4720
rect 149881 4662 178467 4664
rect 149881 4659 149947 4662
rect 178401 4659 178467 4662
rect 212165 4722 212231 4725
rect 214741 4722 214807 4725
rect 212165 4720 214807 4722
rect 212165 4664 212170 4720
rect 212226 4664 214746 4720
rect 214802 4664 214807 4720
rect 212165 4662 214807 4664
rect 212165 4659 212231 4662
rect 214741 4659 214807 4662
rect 218973 4722 219039 4725
rect 245929 4722 245995 4725
rect 218973 4720 245995 4722
rect 218973 4664 218978 4720
rect 219034 4664 245934 4720
rect 245990 4664 245995 4720
rect 218973 4662 245995 4664
rect 218973 4659 219039 4662
rect 245929 4659 245995 4662
rect 268285 4722 268351 4725
rect 268285 4720 272504 4722
rect 268285 4664 268290 4720
rect 268346 4664 272504 4720
rect 268285 4662 272504 4664
rect 268285 4659 268351 4662
rect 43529 4586 43595 4589
rect 100017 4586 100083 4589
rect 43529 4584 100083 4586
rect 43529 4528 43534 4584
rect 43590 4528 100022 4584
rect 100078 4528 100083 4584
rect 43529 4526 100083 4528
rect 43529 4523 43595 4526
rect 100017 4523 100083 4526
rect 105445 4586 105511 4589
rect 106089 4586 106155 4589
rect 105445 4584 106155 4586
rect 105445 4528 105450 4584
rect 105506 4528 106094 4584
rect 106150 4528 106155 4584
rect 105445 4526 106155 4528
rect 105445 4523 105511 4526
rect 106089 4523 106155 4526
rect 114553 4586 114619 4589
rect 154573 4586 154639 4589
rect 220813 4586 220879 4589
rect 114553 4584 220879 4586
rect 114553 4528 114558 4584
rect 114614 4528 154578 4584
rect 154634 4528 220818 4584
rect 220874 4528 220879 4584
rect 114553 4526 220879 4528
rect 114553 4523 114619 4526
rect 154573 4523 154639 4526
rect 220813 4523 220879 4526
rect 226190 4524 226196 4588
rect 226260 4586 226266 4588
rect 227621 4586 227687 4589
rect 226260 4584 227687 4586
rect 226260 4528 227626 4584
rect 227682 4528 227687 4584
rect 226260 4526 227687 4528
rect 226260 4524 226266 4526
rect 227621 4523 227687 4526
rect 227805 4586 227871 4589
rect 255129 4586 255195 4589
rect 227805 4584 255195 4586
rect 227805 4528 227810 4584
rect 227866 4528 255134 4584
rect 255190 4528 255195 4584
rect 227805 4526 255195 4528
rect 227805 4523 227871 4526
rect 255129 4523 255195 4526
rect 267733 4586 267799 4589
rect 267733 4584 271890 4586
rect 267733 4528 267738 4584
rect 267794 4528 271890 4584
rect 267733 4526 271890 4528
rect 272304 4526 272504 4586
rect 267733 4523 267799 4526
rect 80053 4450 80119 4453
rect 96521 4450 96587 4453
rect 80053 4448 96587 4450
rect 80053 4392 80058 4448
rect 80114 4392 96526 4448
rect 96582 4392 96587 4448
rect 80053 4390 96587 4392
rect 80053 4387 80119 4390
rect 96521 4387 96587 4390
rect 99833 4450 99899 4453
rect 139209 4450 139275 4453
rect 139853 4450 139919 4453
rect 99833 4448 109050 4450
rect 99833 4392 99838 4448
rect 99894 4392 109050 4448
rect 99833 4390 109050 4392
rect 99833 4387 99899 4390
rect 68542 4384 68858 4385
rect 68542 4320 68548 4384
rect 68612 4320 68628 4384
rect 68692 4320 68708 4384
rect 68772 4320 68788 4384
rect 68852 4320 68858 4384
rect 68542 4319 68858 4320
rect 92657 4314 92723 4317
rect 102041 4314 102107 4317
rect 92657 4312 102107 4314
rect 92657 4256 92662 4312
rect 92718 4256 102046 4312
rect 102102 4256 102107 4312
rect 92657 4254 102107 4256
rect 92657 4251 92723 4254
rect 102041 4251 102107 4254
rect 106273 4314 106339 4317
rect 107193 4314 107259 4317
rect 106273 4312 107259 4314
rect 106273 4256 106278 4312
rect 106334 4256 107198 4312
rect 107254 4256 107259 4312
rect 106273 4254 107259 4256
rect 106273 4251 106339 4254
rect 107193 4251 107259 4254
rect 42609 4178 42675 4181
rect 47117 4178 47183 4181
rect 42609 4176 47183 4178
rect 42609 4120 42614 4176
rect 42670 4120 47122 4176
rect 47178 4120 47183 4176
rect 42609 4118 47183 4120
rect 42609 4115 42675 4118
rect 47117 4115 47183 4118
rect 92749 4178 92815 4181
rect 95509 4178 95575 4181
rect 92749 4176 95575 4178
rect 92749 4120 92754 4176
rect 92810 4120 95514 4176
rect 95570 4120 95575 4176
rect 92749 4118 95575 4120
rect 92749 4115 92815 4118
rect 95509 4115 95575 4118
rect 96470 4116 96476 4180
rect 96540 4178 96546 4180
rect 102225 4178 102291 4181
rect 96540 4176 102291 4178
rect 96540 4120 102230 4176
rect 102286 4120 102291 4176
rect 96540 4118 102291 4120
rect 108990 4178 109050 4390
rect 139209 4448 139919 4450
rect 139209 4392 139214 4448
rect 139270 4392 139858 4448
rect 139914 4392 139919 4448
rect 139209 4390 139919 4392
rect 139209 4387 139275 4390
rect 139853 4387 139919 4390
rect 141601 4450 141667 4453
rect 169661 4450 169727 4453
rect 141601 4448 169727 4450
rect 141601 4392 141606 4448
rect 141662 4392 169666 4448
rect 169722 4392 169727 4448
rect 141601 4390 169727 4392
rect 141601 4387 141667 4390
rect 169661 4387 169727 4390
rect 219433 4450 219499 4453
rect 256417 4450 256483 4453
rect 219433 4448 256483 4450
rect 219433 4392 219438 4448
rect 219494 4392 256422 4448
rect 256478 4392 256483 4448
rect 219433 4390 256483 4392
rect 219433 4387 219499 4390
rect 256417 4387 256483 4390
rect 260005 4450 260071 4453
rect 267273 4450 267339 4453
rect 260005 4448 267339 4450
rect 260005 4392 260010 4448
rect 260066 4392 267278 4448
rect 267334 4392 267339 4448
rect 260005 4390 267339 4392
rect 260005 4387 260071 4390
rect 267273 4387 267339 4390
rect 268469 4450 268535 4453
rect 271137 4450 271203 4453
rect 268469 4448 271203 4450
rect 268469 4392 268474 4448
rect 268530 4392 271142 4448
rect 271198 4392 271203 4448
rect 268469 4390 271203 4392
rect 271830 4450 271890 4526
rect 271830 4390 272504 4450
rect 268469 4387 268535 4390
rect 271137 4387 271203 4390
rect 136139 4384 136455 4385
rect 136139 4320 136145 4384
rect 136209 4320 136225 4384
rect 136289 4320 136305 4384
rect 136369 4320 136385 4384
rect 136449 4320 136455 4384
rect 136139 4319 136455 4320
rect 203736 4384 204052 4385
rect 203736 4320 203742 4384
rect 203806 4320 203822 4384
rect 203886 4320 203902 4384
rect 203966 4320 203982 4384
rect 204046 4320 204052 4384
rect 203736 4319 204052 4320
rect 271333 4384 271649 4385
rect 271333 4320 271339 4384
rect 271403 4320 271419 4384
rect 271483 4320 271499 4384
rect 271563 4320 271579 4384
rect 271643 4320 271649 4384
rect 271333 4319 271649 4320
rect 150065 4314 150131 4317
rect 173801 4314 173867 4317
rect 150065 4312 173867 4314
rect 150065 4256 150070 4312
rect 150126 4256 173806 4312
rect 173862 4256 173867 4312
rect 150065 4254 173867 4256
rect 150065 4251 150131 4254
rect 173801 4251 173867 4254
rect 219065 4314 219131 4317
rect 223113 4314 223179 4317
rect 227713 4314 227779 4317
rect 219065 4312 227779 4314
rect 219065 4256 219070 4312
rect 219126 4256 223118 4312
rect 223174 4256 227718 4312
rect 227774 4256 227779 4312
rect 219065 4254 227779 4256
rect 219065 4251 219131 4254
rect 223113 4251 223179 4254
rect 227713 4251 227779 4254
rect 237281 4314 237347 4317
rect 248873 4314 248939 4317
rect 237281 4312 248939 4314
rect 237281 4256 237286 4312
rect 237342 4256 248878 4312
rect 248934 4256 248939 4312
rect 237281 4254 248939 4256
rect 237281 4251 237347 4254
rect 248873 4251 248939 4254
rect 249057 4314 249123 4317
rect 250161 4314 250227 4317
rect 249057 4312 250227 4314
rect 249057 4256 249062 4312
rect 249118 4256 250166 4312
rect 250222 4256 250227 4312
rect 249057 4254 250227 4256
rect 249057 4251 249123 4254
rect 250161 4251 250227 4254
rect 252645 4314 252711 4317
rect 271781 4314 271847 4317
rect 252645 4312 271154 4314
rect 252645 4256 252650 4312
rect 252706 4256 271154 4312
rect 252645 4254 271154 4256
rect 252645 4251 252711 4254
rect 141509 4178 141575 4181
rect 108990 4176 141575 4178
rect 108990 4120 141514 4176
rect 141570 4120 141575 4176
rect 108990 4118 141575 4120
rect 96540 4116 96546 4118
rect 102225 4115 102291 4118
rect 141509 4115 141575 4118
rect 145557 4178 145623 4181
rect 154021 4178 154087 4181
rect 145557 4176 154087 4178
rect 145557 4120 145562 4176
rect 145618 4120 154026 4176
rect 154082 4120 154087 4176
rect 145557 4118 154087 4120
rect 145557 4115 145623 4118
rect 154021 4115 154087 4118
rect 169569 4178 169635 4181
rect 219249 4178 219315 4181
rect 229001 4178 229067 4181
rect 169569 4176 219315 4178
rect 169569 4120 169574 4176
rect 169630 4120 219254 4176
rect 219310 4120 219315 4176
rect 169569 4118 219315 4120
rect 169569 4115 169635 4118
rect 219249 4115 219315 4118
rect 224726 4176 229067 4178
rect 224726 4120 229006 4176
rect 229062 4120 229067 4176
rect 224726 4118 229067 4120
rect 224726 4045 224786 4118
rect 229001 4115 229067 4118
rect 243077 4178 243143 4181
rect 248781 4178 248847 4181
rect 243077 4176 248847 4178
rect 243077 4120 243082 4176
rect 243138 4120 248786 4176
rect 248842 4120 248847 4176
rect 243077 4118 248847 4120
rect 243077 4115 243143 4118
rect 248781 4115 248847 4118
rect 260833 4178 260899 4181
rect 271094 4178 271154 4254
rect 271781 4312 272504 4314
rect 271781 4256 271786 4312
rect 271842 4256 272504 4312
rect 271781 4254 272504 4256
rect 271781 4251 271847 4254
rect 271689 4178 271755 4181
rect 260833 4176 270970 4178
rect 260833 4120 260838 4176
rect 260894 4120 270970 4176
rect 260833 4118 270970 4120
rect 271094 4176 271755 4178
rect 271094 4120 271694 4176
rect 271750 4120 271755 4176
rect 271094 4118 271755 4120
rect 260833 4115 260899 4118
rect 38929 4042 38995 4045
rect 92933 4042 92999 4045
rect 97625 4042 97691 4045
rect 38929 4040 80070 4042
rect 38929 3984 38934 4040
rect 38990 3984 80070 4040
rect 38929 3982 80070 3984
rect 38929 3979 38995 3982
rect 80010 3906 80070 3982
rect 92933 4040 97691 4042
rect 92933 3984 92938 4040
rect 92994 3984 97630 4040
rect 97686 3984 97691 4040
rect 92933 3982 97691 3984
rect 92933 3979 92999 3982
rect 97625 3979 97691 3982
rect 100293 4042 100359 4045
rect 100293 4040 102794 4042
rect 100293 3984 100298 4040
rect 100354 3984 102794 4040
rect 100293 3982 102794 3984
rect 100293 3979 100359 3982
rect 96613 3906 96679 3909
rect 80010 3904 96679 3906
rect 80010 3848 96618 3904
rect 96674 3848 96679 3904
rect 80010 3846 96679 3848
rect 102734 3906 102794 3982
rect 103278 3980 103284 4044
rect 103348 4042 103354 4044
rect 103421 4042 103487 4045
rect 103348 4040 103487 4042
rect 103348 3984 103426 4040
rect 103482 3984 103487 4040
rect 103348 3982 103487 3984
rect 103348 3980 103354 3982
rect 103421 3979 103487 3982
rect 104525 4044 104591 4045
rect 104525 4040 104572 4044
rect 104636 4042 104642 4044
rect 104525 3984 104530 4040
rect 104525 3980 104572 3984
rect 104636 3982 104682 4042
rect 104636 3980 104642 3982
rect 105486 3980 105492 4044
rect 105556 4042 105562 4044
rect 105629 4042 105695 4045
rect 105556 4040 105695 4042
rect 105556 3984 105634 4040
rect 105690 3984 105695 4040
rect 105556 3982 105695 3984
rect 105556 3980 105562 3982
rect 104525 3979 104591 3980
rect 105629 3979 105695 3982
rect 106958 3980 106964 4044
rect 107028 4042 107034 4044
rect 107101 4042 107167 4045
rect 107028 4040 107167 4042
rect 107028 3984 107106 4040
rect 107162 3984 107167 4040
rect 107028 3982 107167 3984
rect 107028 3980 107034 3982
rect 107101 3979 107167 3982
rect 107561 4042 107627 4045
rect 107694 4042 107700 4044
rect 107561 4040 107700 4042
rect 107561 3984 107566 4040
rect 107622 3984 107700 4040
rect 107561 3982 107700 3984
rect 107561 3979 107627 3982
rect 107694 3980 107700 3982
rect 107764 3980 107770 4044
rect 108021 4042 108087 4045
rect 109217 4044 109283 4045
rect 108246 4042 108252 4044
rect 108021 4040 108252 4042
rect 108021 3984 108026 4040
rect 108082 3984 108252 4040
rect 108021 3982 108252 3984
rect 108021 3979 108087 3982
rect 108246 3980 108252 3982
rect 108316 3980 108322 4044
rect 109166 3980 109172 4044
rect 109236 4042 109283 4044
rect 109236 4040 109328 4042
rect 109278 3984 109328 4040
rect 109236 3982 109328 3984
rect 109236 3980 109283 3982
rect 109902 3980 109908 4044
rect 109972 4042 109978 4044
rect 110045 4042 110111 4045
rect 110689 4044 110755 4045
rect 111241 4044 111307 4045
rect 110638 4042 110644 4044
rect 109972 4040 110111 4042
rect 109972 3984 110050 4040
rect 110106 3984 110111 4040
rect 109972 3982 110111 3984
rect 110598 3982 110644 4042
rect 110708 4040 110755 4044
rect 111190 4042 111196 4044
rect 110750 3984 110755 4040
rect 109972 3980 109978 3982
rect 109217 3979 109283 3980
rect 110045 3979 110111 3982
rect 110638 3980 110644 3982
rect 110708 3980 110755 3984
rect 111150 3982 111196 4042
rect 111260 4040 111307 4044
rect 111302 3984 111307 4040
rect 111190 3980 111196 3982
rect 111260 3980 111307 3984
rect 112110 3980 112116 4044
rect 112180 4042 112186 4044
rect 112345 4042 112411 4045
rect 112180 4040 112411 4042
rect 112180 3984 112350 4040
rect 112406 3984 112411 4040
rect 112180 3982 112411 3984
rect 112180 3980 112186 3982
rect 110689 3979 110755 3980
rect 111241 3979 111307 3980
rect 112345 3979 112411 3982
rect 112846 3980 112852 4044
rect 112916 4042 112922 4044
rect 112989 4042 113055 4045
rect 112916 4040 113055 4042
rect 112916 3984 112994 4040
rect 113050 3984 113055 4040
rect 112916 3982 113055 3984
rect 112916 3980 112922 3982
rect 112989 3979 113055 3982
rect 113214 3980 113220 4044
rect 113284 4042 113290 4044
rect 140957 4042 141023 4045
rect 141785 4042 141851 4045
rect 113284 4040 141851 4042
rect 113284 3984 140962 4040
rect 141018 3984 141790 4040
rect 141846 3984 141851 4040
rect 113284 3982 141851 3984
rect 113284 3980 113290 3982
rect 140957 3979 141023 3982
rect 141785 3979 141851 3982
rect 151997 4042 152063 4045
rect 215201 4044 215267 4045
rect 153142 4042 153148 4044
rect 151997 4040 153148 4042
rect 151997 3984 152002 4040
rect 152058 3984 153148 4040
rect 151997 3982 153148 3984
rect 151997 3979 152063 3982
rect 153142 3980 153148 3982
rect 153212 3980 153218 4044
rect 215150 4042 215156 4044
rect 215110 3982 215156 4042
rect 215220 4040 215267 4044
rect 215262 3984 215267 4040
rect 215150 3980 215156 3982
rect 215220 3980 215267 3984
rect 215201 3979 215267 3980
rect 218237 4042 218303 4045
rect 221733 4042 221799 4045
rect 218237 4040 221799 4042
rect 218237 3984 218242 4040
rect 218298 3984 221738 4040
rect 221794 3984 221799 4040
rect 218237 3982 221799 3984
rect 218237 3979 218303 3982
rect 221733 3979 221799 3982
rect 222193 4042 222259 4045
rect 223982 4042 223988 4044
rect 222193 4040 223988 4042
rect 222193 3984 222198 4040
rect 222254 3984 223988 4040
rect 222193 3982 223988 3984
rect 222193 3979 222259 3982
rect 223982 3980 223988 3982
rect 224052 3980 224058 4044
rect 224677 4040 224786 4045
rect 266261 4042 266327 4045
rect 270769 4042 270835 4045
rect 224677 3984 224682 4040
rect 224738 3984 224786 4040
rect 224677 3982 224786 3984
rect 224910 3982 244290 4042
rect 224677 3979 224743 3982
rect 102734 3846 103898 3906
rect 96613 3843 96679 3846
rect 34744 3840 35060 3841
rect 34744 3776 34750 3840
rect 34814 3776 34830 3840
rect 34894 3776 34910 3840
rect 34974 3776 34990 3840
rect 35054 3776 35060 3840
rect 34744 3775 35060 3776
rect 102341 3840 102657 3841
rect 102341 3776 102347 3840
rect 102411 3776 102427 3840
rect 102491 3776 102507 3840
rect 102571 3776 102587 3840
rect 102651 3776 102657 3840
rect 102341 3775 102657 3776
rect 92565 3770 92631 3773
rect 95233 3770 95299 3773
rect 92565 3768 95299 3770
rect 92565 3712 92570 3768
rect 92626 3712 95238 3768
rect 95294 3712 95299 3768
rect 92565 3710 95299 3712
rect 92565 3707 92631 3710
rect 95233 3707 95299 3710
rect 97533 3770 97599 3773
rect 97758 3770 97764 3772
rect 97533 3768 97764 3770
rect 97533 3712 97538 3768
rect 97594 3712 97764 3768
rect 97533 3710 97764 3712
rect 97533 3707 97599 3710
rect 97758 3708 97764 3710
rect 97828 3708 97834 3772
rect 48773 3634 48839 3637
rect 51625 3634 51691 3637
rect 48773 3632 51691 3634
rect 48773 3576 48778 3632
rect 48834 3576 51630 3632
rect 51686 3576 51691 3632
rect 48773 3574 51691 3576
rect 48773 3571 48839 3574
rect 51625 3571 51691 3574
rect 78581 3634 78647 3637
rect 103697 3634 103763 3637
rect 78581 3632 103763 3634
rect 78581 3576 78586 3632
rect 78642 3576 103702 3632
rect 103758 3576 103763 3632
rect 78581 3574 103763 3576
rect 103838 3634 103898 3846
rect 104014 3844 104020 3908
rect 104084 3906 104090 3908
rect 104617 3906 104683 3909
rect 104084 3904 104683 3906
rect 104084 3848 104622 3904
rect 104678 3848 104683 3904
rect 104084 3846 104683 3848
rect 104084 3844 104090 3846
rect 104617 3843 104683 3846
rect 104893 3906 104959 3909
rect 143533 3906 143599 3909
rect 104893 3904 143599 3906
rect 104893 3848 104898 3904
rect 104954 3848 143538 3904
rect 143594 3848 143599 3904
rect 104893 3846 143599 3848
rect 104893 3843 104959 3846
rect 143533 3843 143599 3846
rect 152365 3906 152431 3909
rect 161289 3906 161355 3909
rect 152365 3904 161355 3906
rect 152365 3848 152370 3904
rect 152426 3848 161294 3904
rect 161350 3848 161355 3904
rect 152365 3846 161355 3848
rect 152365 3843 152431 3846
rect 161289 3843 161355 3846
rect 209313 3906 209379 3909
rect 224910 3906 224970 3982
rect 209313 3904 224970 3906
rect 209313 3848 209318 3904
rect 209374 3848 224970 3904
rect 209313 3846 224970 3848
rect 209313 3843 209379 3846
rect 226006 3844 226012 3908
rect 226076 3906 226082 3908
rect 228541 3906 228607 3909
rect 226076 3904 228607 3906
rect 226076 3848 228546 3904
rect 228602 3848 228607 3904
rect 226076 3846 228607 3848
rect 244230 3906 244290 3982
rect 266261 4040 270835 4042
rect 266261 3984 266266 4040
rect 266322 3984 270774 4040
rect 270830 3984 270835 4040
rect 266261 3982 270835 3984
rect 270910 4042 270970 4118
rect 271689 4115 271755 4118
rect 271830 4118 272504 4178
rect 271830 4042 271890 4118
rect 270910 3982 271890 4042
rect 272014 3982 272504 4042
rect 266261 3979 266327 3982
rect 270769 3979 270835 3982
rect 248689 3906 248755 3909
rect 272014 3906 272074 3982
rect 244230 3904 248755 3906
rect 244230 3848 248694 3904
rect 248750 3848 248755 3904
rect 244230 3846 248755 3848
rect 226076 3844 226082 3846
rect 228541 3843 228607 3846
rect 248689 3843 248755 3846
rect 267782 3846 272074 3906
rect 272149 3906 272215 3909
rect 272149 3904 272504 3906
rect 272149 3848 272154 3904
rect 272210 3848 272504 3904
rect 272149 3846 272504 3848
rect 169938 3840 170254 3841
rect 169938 3776 169944 3840
rect 170008 3776 170024 3840
rect 170088 3776 170104 3840
rect 170168 3776 170184 3840
rect 170248 3776 170254 3840
rect 169938 3775 170254 3776
rect 237535 3840 237851 3841
rect 237535 3776 237541 3840
rect 237605 3776 237621 3840
rect 237685 3776 237701 3840
rect 237765 3776 237781 3840
rect 237845 3776 237851 3840
rect 237535 3775 237851 3776
rect 267782 3773 267842 3846
rect 272149 3843 272215 3846
rect 104433 3770 104499 3773
rect 104985 3770 105051 3773
rect 104433 3768 105051 3770
rect 104433 3712 104438 3768
rect 104494 3712 104990 3768
rect 105046 3712 105051 3768
rect 104433 3710 105051 3712
rect 104433 3707 104499 3710
rect 104985 3707 105051 3710
rect 105813 3770 105879 3773
rect 107142 3770 107148 3772
rect 105813 3768 107148 3770
rect 105813 3712 105818 3768
rect 105874 3712 107148 3768
rect 105813 3710 107148 3712
rect 105813 3707 105879 3710
rect 107142 3708 107148 3710
rect 107212 3708 107218 3772
rect 108849 3770 108915 3773
rect 146661 3770 146727 3773
rect 156137 3770 156203 3773
rect 157241 3770 157307 3773
rect 218881 3772 218947 3773
rect 218830 3770 218836 3772
rect 108849 3768 118710 3770
rect 108849 3712 108854 3768
rect 108910 3712 118710 3768
rect 108849 3710 118710 3712
rect 108849 3707 108915 3710
rect 115013 3634 115079 3637
rect 103838 3632 115079 3634
rect 103838 3576 115018 3632
rect 115074 3576 115079 3632
rect 103838 3574 115079 3576
rect 118650 3634 118710 3710
rect 146661 3768 157307 3770
rect 146661 3712 146666 3768
rect 146722 3712 156142 3768
rect 156198 3712 157246 3768
rect 157302 3712 157307 3768
rect 146661 3710 157307 3712
rect 218790 3710 218836 3770
rect 218900 3768 218947 3772
rect 218942 3712 218947 3768
rect 146661 3707 146727 3710
rect 156137 3707 156203 3710
rect 157241 3707 157307 3710
rect 218830 3708 218836 3710
rect 218900 3708 218947 3712
rect 218881 3707 218947 3708
rect 220813 3770 220879 3773
rect 222101 3770 222167 3773
rect 220813 3768 222167 3770
rect 220813 3712 220818 3768
rect 220874 3712 222106 3768
rect 222162 3712 222167 3768
rect 220813 3710 222167 3712
rect 220813 3707 220879 3710
rect 222101 3707 222167 3710
rect 223246 3708 223252 3772
rect 223316 3770 223322 3772
rect 223481 3770 223547 3773
rect 224953 3770 225019 3773
rect 223316 3768 223547 3770
rect 223316 3712 223486 3768
rect 223542 3712 223547 3768
rect 223316 3710 223547 3712
rect 223316 3708 223322 3710
rect 223481 3707 223547 3710
rect 223806 3768 225019 3770
rect 223806 3712 224958 3768
rect 225014 3712 225019 3768
rect 223806 3710 225019 3712
rect 146385 3634 146451 3637
rect 118650 3632 146451 3634
rect 118650 3576 146390 3632
rect 146446 3576 146451 3632
rect 118650 3574 146451 3576
rect 78581 3571 78647 3574
rect 103697 3571 103763 3574
rect 115013 3571 115079 3574
rect 146385 3571 146451 3574
rect 150341 3634 150407 3637
rect 160001 3634 160067 3637
rect 222009 3634 222075 3637
rect 223806 3634 223866 3710
rect 224953 3707 225019 3710
rect 227294 3708 227300 3772
rect 227364 3770 227370 3772
rect 227621 3770 227687 3773
rect 227364 3768 227687 3770
rect 227364 3712 227626 3768
rect 227682 3712 227687 3768
rect 227364 3710 227687 3712
rect 227364 3708 227370 3710
rect 227621 3707 227687 3710
rect 239397 3770 239463 3773
rect 259269 3770 259335 3773
rect 239397 3768 259335 3770
rect 239397 3712 239402 3768
rect 239458 3712 259274 3768
rect 259330 3712 259335 3768
rect 239397 3710 259335 3712
rect 239397 3707 239463 3710
rect 259269 3707 259335 3710
rect 267733 3768 267842 3773
rect 267733 3712 267738 3768
rect 267794 3712 267842 3768
rect 267733 3710 267842 3712
rect 268009 3770 268075 3773
rect 268009 3768 272504 3770
rect 268009 3712 268014 3768
rect 268070 3712 272504 3768
rect 268009 3710 272504 3712
rect 267733 3707 267799 3710
rect 268009 3707 268075 3710
rect 150341 3632 222075 3634
rect 150341 3576 150346 3632
rect 150402 3576 160006 3632
rect 160062 3576 222014 3632
rect 222070 3576 222075 3632
rect 150341 3574 222075 3576
rect 150341 3571 150407 3574
rect 160001 3571 160067 3574
rect 222009 3571 222075 3574
rect 222150 3574 223866 3634
rect 15101 3498 15167 3501
rect 49325 3498 49391 3501
rect 15101 3496 49391 3498
rect 15101 3440 15106 3496
rect 15162 3440 49330 3496
rect 49386 3440 49391 3496
rect 15101 3438 49391 3440
rect 15101 3435 15167 3438
rect 49325 3435 49391 3438
rect 51809 3498 51875 3501
rect 100293 3498 100359 3501
rect 51809 3496 100359 3498
rect 51809 3440 51814 3496
rect 51870 3440 100298 3496
rect 100354 3440 100359 3496
rect 51809 3438 100359 3440
rect 51809 3435 51875 3438
rect 100293 3435 100359 3438
rect 100477 3498 100543 3501
rect 103145 3498 103211 3501
rect 100477 3496 103211 3498
rect 100477 3440 100482 3496
rect 100538 3440 103150 3496
rect 103206 3440 103211 3496
rect 100477 3438 103211 3440
rect 100477 3435 100543 3438
rect 103145 3435 103211 3438
rect 106181 3498 106247 3501
rect 107377 3498 107443 3501
rect 106181 3496 107443 3498
rect 106181 3440 106186 3496
rect 106242 3440 107382 3496
rect 107438 3440 107443 3496
rect 106181 3438 107443 3440
rect 106181 3435 106247 3438
rect 107377 3435 107443 3438
rect 108113 3498 108179 3501
rect 113357 3498 113423 3501
rect 108113 3496 113423 3498
rect 108113 3440 108118 3496
rect 108174 3440 113362 3496
rect 113418 3440 113423 3496
rect 108113 3438 113423 3440
rect 108113 3435 108179 3438
rect 113357 3435 113423 3438
rect 139945 3498 140011 3501
rect 146477 3498 146543 3501
rect 139945 3496 146543 3498
rect 139945 3440 139950 3496
rect 140006 3440 146482 3496
rect 146538 3440 146543 3496
rect 139945 3438 146543 3440
rect 139945 3435 140011 3438
rect 146477 3435 146543 3438
rect 147213 3498 147279 3501
rect 217041 3498 217107 3501
rect 222150 3498 222210 3574
rect 223982 3572 223988 3636
rect 224052 3634 224058 3636
rect 227713 3634 227779 3637
rect 224052 3632 227779 3634
rect 224052 3576 227718 3632
rect 227774 3576 227779 3632
rect 224052 3574 227779 3576
rect 224052 3572 224058 3574
rect 227713 3571 227779 3574
rect 228725 3634 228791 3637
rect 229921 3634 229987 3637
rect 228725 3632 229987 3634
rect 228725 3576 228730 3632
rect 228786 3576 229926 3632
rect 229982 3576 229987 3632
rect 228725 3574 229987 3576
rect 228725 3571 228791 3574
rect 229921 3571 229987 3574
rect 231853 3634 231919 3637
rect 254025 3634 254091 3637
rect 231853 3632 254091 3634
rect 231853 3576 231858 3632
rect 231914 3576 254030 3632
rect 254086 3576 254091 3632
rect 231853 3574 254091 3576
rect 231853 3571 231919 3574
rect 254025 3571 254091 3574
rect 268837 3634 268903 3637
rect 272149 3634 272215 3637
rect 268837 3632 272074 3634
rect 268837 3576 268842 3632
rect 268898 3576 272074 3632
rect 268837 3574 272074 3576
rect 268837 3571 268903 3574
rect 147213 3496 222210 3498
rect 147213 3440 147218 3496
rect 147274 3440 217046 3496
rect 217102 3440 222210 3496
rect 147213 3438 222210 3440
rect 223573 3498 223639 3501
rect 248137 3498 248203 3501
rect 223573 3496 248203 3498
rect 223573 3440 223578 3496
rect 223634 3440 248142 3496
rect 248198 3440 248203 3496
rect 223573 3438 248203 3440
rect 147213 3435 147279 3438
rect 217041 3435 217107 3438
rect 223573 3435 223639 3438
rect 248137 3435 248203 3438
rect 258441 3498 258507 3501
rect 267549 3498 267615 3501
rect 258441 3496 267615 3498
rect 258441 3440 258446 3496
rect 258502 3440 267554 3496
rect 267610 3440 267615 3496
rect 258441 3438 267615 3440
rect 258441 3435 258507 3438
rect 267549 3435 267615 3438
rect 268009 3498 268075 3501
rect 272014 3498 272074 3574
rect 272149 3632 272504 3634
rect 272149 3576 272154 3632
rect 272210 3576 272504 3632
rect 272149 3574 272504 3576
rect 272149 3571 272215 3574
rect 268009 3496 271890 3498
rect 268009 3440 268014 3496
rect 268070 3440 271890 3496
rect 268009 3438 271890 3440
rect 272014 3438 272504 3498
rect 268009 3435 268075 3438
rect 47577 3362 47643 3365
rect 48221 3362 48287 3365
rect 47577 3360 48287 3362
rect 47577 3304 47582 3360
rect 47638 3304 48226 3360
rect 48282 3304 48287 3360
rect 47577 3302 48287 3304
rect 47577 3299 47643 3302
rect 48221 3299 48287 3302
rect 84101 3362 84167 3365
rect 117221 3362 117287 3365
rect 84101 3360 117287 3362
rect 84101 3304 84106 3360
rect 84162 3304 117226 3360
rect 117282 3304 117287 3360
rect 84101 3302 117287 3304
rect 84101 3299 84167 3302
rect 117221 3299 117287 3302
rect 144821 3362 144887 3365
rect 152917 3362 152983 3365
rect 154297 3364 154363 3365
rect 154246 3362 154252 3364
rect 144821 3360 152983 3362
rect 144821 3304 144826 3360
rect 144882 3304 152922 3360
rect 152978 3304 152983 3360
rect 144821 3302 152983 3304
rect 154206 3302 154252 3362
rect 154316 3360 154363 3364
rect 154358 3304 154363 3360
rect 144821 3299 144887 3302
rect 152917 3299 152983 3302
rect 154246 3300 154252 3302
rect 154316 3300 154363 3304
rect 154297 3299 154363 3300
rect 219157 3362 219223 3365
rect 227621 3362 227687 3365
rect 245469 3362 245535 3365
rect 259729 3362 259795 3365
rect 219157 3360 227687 3362
rect 219157 3304 219162 3360
rect 219218 3304 227626 3360
rect 227682 3304 227687 3360
rect 219157 3302 227687 3304
rect 219157 3299 219223 3302
rect 227621 3299 227687 3302
rect 229694 3360 245535 3362
rect 229694 3304 245474 3360
rect 245530 3304 245535 3360
rect 229694 3302 245535 3304
rect 68542 3296 68858 3297
rect 68542 3232 68548 3296
rect 68612 3232 68628 3296
rect 68692 3232 68708 3296
rect 68772 3232 68788 3296
rect 68852 3232 68858 3296
rect 68542 3231 68858 3232
rect 136139 3296 136455 3297
rect 136139 3232 136145 3296
rect 136209 3232 136225 3296
rect 136289 3232 136305 3296
rect 136369 3232 136385 3296
rect 136449 3232 136455 3296
rect 136139 3231 136455 3232
rect 203736 3296 204052 3297
rect 203736 3232 203742 3296
rect 203806 3232 203822 3296
rect 203886 3232 203902 3296
rect 203966 3232 203982 3296
rect 204046 3232 204052 3296
rect 203736 3231 204052 3232
rect 14365 3226 14431 3229
rect 49049 3226 49115 3229
rect 14365 3224 49115 3226
rect 14365 3168 14370 3224
rect 14426 3168 49054 3224
rect 49110 3168 49115 3224
rect 14365 3166 49115 3168
rect 14365 3163 14431 3166
rect 49049 3163 49115 3166
rect 93894 3164 93900 3228
rect 93964 3226 93970 3228
rect 94865 3226 94931 3229
rect 93964 3224 94931 3226
rect 93964 3168 94870 3224
rect 94926 3168 94931 3224
rect 93964 3166 94931 3168
rect 93964 3164 93970 3166
rect 94865 3163 94931 3166
rect 95233 3226 95299 3229
rect 96286 3226 96292 3228
rect 95233 3224 96292 3226
rect 95233 3168 95238 3224
rect 95294 3168 96292 3224
rect 95233 3166 96292 3168
rect 95233 3163 95299 3166
rect 96286 3164 96292 3166
rect 96356 3164 96362 3228
rect 96838 3164 96844 3228
rect 96908 3226 96914 3228
rect 100477 3226 100543 3229
rect 100753 3228 100819 3229
rect 100702 3226 100708 3228
rect 96908 3224 100543 3226
rect 96908 3168 100482 3224
rect 100538 3168 100543 3224
rect 96908 3166 100543 3168
rect 100662 3166 100708 3226
rect 100772 3224 100819 3228
rect 100814 3168 100819 3224
rect 96908 3164 96914 3166
rect 100477 3163 100543 3166
rect 100702 3164 100708 3166
rect 100772 3164 100819 3168
rect 100753 3163 100819 3164
rect 101029 3226 101095 3229
rect 101213 3226 101279 3229
rect 104893 3226 104959 3229
rect 101029 3224 104959 3226
rect 101029 3168 101034 3224
rect 101090 3168 101218 3224
rect 101274 3168 104898 3224
rect 104954 3168 104959 3224
rect 101029 3166 104959 3168
rect 101029 3163 101095 3166
rect 101213 3163 101279 3166
rect 104893 3163 104959 3166
rect 108941 3226 109007 3229
rect 144729 3228 144795 3229
rect 110270 3226 110276 3228
rect 108941 3224 110276 3226
rect 108941 3168 108946 3224
rect 109002 3168 110276 3224
rect 108941 3166 110276 3168
rect 108941 3163 109007 3166
rect 110270 3164 110276 3166
rect 110340 3164 110346 3228
rect 144678 3226 144684 3228
rect 144638 3166 144684 3226
rect 144748 3224 144795 3228
rect 144790 3168 144795 3224
rect 144678 3164 144684 3166
rect 144748 3164 144795 3168
rect 144729 3163 144795 3164
rect 149605 3226 149671 3229
rect 151997 3226 152063 3229
rect 149605 3224 152063 3226
rect 149605 3168 149610 3224
rect 149666 3168 152002 3224
rect 152058 3168 152063 3224
rect 149605 3166 152063 3168
rect 149605 3163 149671 3166
rect 151997 3163 152063 3166
rect 154113 3226 154179 3229
rect 186405 3226 186471 3229
rect 154113 3224 186471 3226
rect 154113 3168 154118 3224
rect 154174 3168 186410 3224
rect 186466 3168 186471 3224
rect 154113 3166 186471 3168
rect 154113 3163 154179 3166
rect 186405 3163 186471 3166
rect 209957 3226 210023 3229
rect 209957 3224 215310 3226
rect 209957 3168 209962 3224
rect 210018 3168 215310 3224
rect 209957 3166 215310 3168
rect 209957 3163 210023 3166
rect 32765 3090 32831 3093
rect 67633 3090 67699 3093
rect 32765 3088 67699 3090
rect 32765 3032 32770 3088
rect 32826 3032 67638 3088
rect 67694 3032 67699 3088
rect 32765 3030 67699 3032
rect 32765 3027 32831 3030
rect 67633 3027 67699 3030
rect 93945 3090 94011 3093
rect 94078 3090 94084 3092
rect 93945 3088 94084 3090
rect 93945 3032 93950 3088
rect 94006 3032 94084 3088
rect 93945 3030 94084 3032
rect 93945 3027 94011 3030
rect 94078 3028 94084 3030
rect 94148 3028 94154 3092
rect 96153 3090 96219 3093
rect 142061 3090 142127 3093
rect 176653 3090 176719 3093
rect 211521 3092 211587 3093
rect 211470 3090 211476 3092
rect 96153 3088 176719 3090
rect 96153 3032 96158 3088
rect 96214 3032 142066 3088
rect 142122 3032 176658 3088
rect 176714 3032 176719 3088
rect 96153 3030 176719 3032
rect 211430 3030 211476 3090
rect 211540 3088 211587 3092
rect 211582 3032 211587 3088
rect 96153 3027 96219 3030
rect 142061 3027 142127 3030
rect 176653 3027 176719 3030
rect 211470 3028 211476 3030
rect 211540 3028 211587 3032
rect 215250 3090 215310 3166
rect 217358 3164 217364 3228
rect 217428 3226 217434 3228
rect 217685 3226 217751 3229
rect 217428 3224 217751 3226
rect 217428 3168 217690 3224
rect 217746 3168 217751 3224
rect 217428 3166 217751 3168
rect 217428 3164 217434 3166
rect 217685 3163 217751 3166
rect 221038 3164 221044 3228
rect 221108 3226 221114 3228
rect 221457 3226 221523 3229
rect 221108 3224 221523 3226
rect 221108 3168 221462 3224
rect 221518 3168 221523 3224
rect 221108 3166 221523 3168
rect 221108 3164 221114 3166
rect 221457 3163 221523 3166
rect 222561 3226 222627 3229
rect 229694 3226 229754 3302
rect 245469 3299 245535 3302
rect 253890 3360 259795 3362
rect 253890 3304 259734 3360
rect 259790 3304 259795 3360
rect 253890 3302 259795 3304
rect 222561 3224 229754 3226
rect 222561 3168 222566 3224
rect 222622 3168 229754 3224
rect 222561 3166 229754 3168
rect 229921 3226 229987 3229
rect 239397 3226 239463 3229
rect 229921 3224 239463 3226
rect 229921 3168 229926 3224
rect 229982 3168 239402 3224
rect 239458 3168 239463 3224
rect 229921 3166 239463 3168
rect 222561 3163 222627 3166
rect 229921 3163 229987 3166
rect 239397 3163 239463 3166
rect 242893 3226 242959 3229
rect 253890 3226 253950 3302
rect 259729 3299 259795 3302
rect 268561 3362 268627 3365
rect 271137 3362 271203 3365
rect 268561 3360 271203 3362
rect 268561 3304 268566 3360
rect 268622 3304 271142 3360
rect 271198 3304 271203 3360
rect 268561 3302 271203 3304
rect 271830 3362 271890 3438
rect 271830 3302 272504 3362
rect 268561 3299 268627 3302
rect 271137 3299 271203 3302
rect 271333 3296 271649 3297
rect 271333 3232 271339 3296
rect 271403 3232 271419 3296
rect 271483 3232 271499 3296
rect 271563 3232 271579 3296
rect 271643 3232 271649 3296
rect 271333 3231 271649 3232
rect 258993 3228 259059 3229
rect 258942 3226 258948 3228
rect 242893 3224 253950 3226
rect 242893 3168 242898 3224
rect 242954 3168 253950 3224
rect 242893 3166 253950 3168
rect 258902 3166 258948 3226
rect 259012 3224 259059 3228
rect 271137 3226 271203 3229
rect 259054 3168 259059 3224
rect 242893 3163 242959 3166
rect 258942 3164 258948 3166
rect 259012 3164 259059 3168
rect 258993 3163 259059 3164
rect 263550 3224 271203 3226
rect 263550 3168 271142 3224
rect 271198 3168 271203 3224
rect 263550 3166 271203 3168
rect 237005 3090 237071 3093
rect 249057 3090 249123 3093
rect 215250 3088 237071 3090
rect 215250 3032 237010 3088
rect 237066 3032 237071 3088
rect 215250 3030 237071 3032
rect 211521 3027 211587 3028
rect 237005 3027 237071 3030
rect 244230 3088 249123 3090
rect 244230 3032 249062 3088
rect 249118 3032 249123 3088
rect 244230 3030 249123 3032
rect 42057 2954 42123 2957
rect 49233 2954 49299 2957
rect 114921 2954 114987 2957
rect 42057 2952 46950 2954
rect 42057 2896 42062 2952
rect 42118 2896 46950 2952
rect 42057 2894 46950 2896
rect 42057 2891 42123 2894
rect 841 2820 907 2821
rect 19241 2820 19307 2821
rect 790 2818 796 2820
rect 750 2758 796 2818
rect 860 2816 907 2820
rect 19190 2818 19196 2820
rect 902 2760 907 2816
rect 790 2756 796 2758
rect 860 2756 907 2760
rect 19150 2758 19196 2818
rect 19260 2816 19307 2820
rect 22829 2820 22895 2821
rect 25037 2820 25103 2821
rect 22829 2818 22876 2820
rect 19302 2760 19307 2816
rect 19190 2756 19196 2758
rect 19260 2756 19307 2760
rect 22784 2816 22876 2818
rect 22784 2760 22834 2816
rect 22784 2758 22876 2760
rect 841 2755 907 2756
rect 19241 2755 19307 2756
rect 22829 2756 22876 2758
rect 22940 2756 22946 2820
rect 25037 2818 25084 2820
rect 24992 2816 25084 2818
rect 24992 2760 25042 2816
rect 24992 2758 25084 2760
rect 25037 2756 25084 2758
rect 25148 2756 25154 2820
rect 27286 2756 27292 2820
rect 27356 2818 27362 2820
rect 27521 2818 27587 2821
rect 27356 2816 27587 2818
rect 27356 2760 27526 2816
rect 27582 2760 27587 2816
rect 27356 2758 27587 2760
rect 46890 2818 46950 2894
rect 49233 2952 114987 2954
rect 49233 2896 49238 2952
rect 49294 2896 114926 2952
rect 114982 2896 114987 2952
rect 49233 2894 114987 2896
rect 49233 2891 49299 2894
rect 114921 2891 114987 2894
rect 143901 2954 143967 2957
rect 143901 2952 147690 2954
rect 143901 2896 143906 2952
rect 143962 2896 147690 2952
rect 143901 2894 147690 2896
rect 143901 2891 143967 2894
rect 52085 2818 52151 2821
rect 46890 2816 52151 2818
rect 46890 2760 52090 2816
rect 52146 2760 52151 2816
rect 46890 2758 52151 2760
rect 27356 2756 27362 2758
rect 22829 2755 22895 2756
rect 25037 2755 25103 2756
rect 27521 2755 27587 2758
rect 52085 2755 52151 2758
rect 54886 2756 54892 2820
rect 54956 2818 54962 2820
rect 55121 2818 55187 2821
rect 54956 2816 55187 2818
rect 54956 2760 55126 2816
rect 55182 2760 55187 2816
rect 54956 2758 55187 2760
rect 54956 2756 54962 2758
rect 55121 2755 55187 2758
rect 95417 2818 95483 2821
rect 96981 2820 97047 2821
rect 95550 2818 95556 2820
rect 95417 2816 95556 2818
rect 95417 2760 95422 2816
rect 95478 2760 95556 2816
rect 95417 2758 95556 2760
rect 95417 2755 95483 2758
rect 95550 2756 95556 2758
rect 95620 2756 95626 2820
rect 96981 2816 97028 2820
rect 97092 2818 97098 2820
rect 104249 2818 104315 2821
rect 105721 2818 105787 2821
rect 96981 2760 96986 2816
rect 96981 2756 97028 2760
rect 97092 2758 97138 2818
rect 104249 2816 105787 2818
rect 104249 2760 104254 2816
rect 104310 2760 105726 2816
rect 105782 2760 105787 2816
rect 104249 2758 105787 2760
rect 97092 2756 97098 2758
rect 96981 2755 97047 2756
rect 104249 2755 104315 2758
rect 105721 2755 105787 2758
rect 109585 2818 109651 2821
rect 111701 2818 111767 2821
rect 109585 2816 111767 2818
rect 109585 2760 109590 2816
rect 109646 2760 111706 2816
rect 111762 2760 111767 2816
rect 109585 2758 111767 2760
rect 109585 2755 109651 2758
rect 111701 2755 111767 2758
rect 116526 2756 116532 2820
rect 116596 2818 116602 2820
rect 117221 2818 117287 2821
rect 116596 2816 117287 2818
rect 116596 2760 117226 2816
rect 117282 2760 117287 2816
rect 116596 2758 117287 2760
rect 116596 2756 116602 2758
rect 117221 2755 117287 2758
rect 123886 2756 123892 2820
rect 123956 2818 123962 2820
rect 124121 2818 124187 2821
rect 123956 2816 124187 2818
rect 123956 2760 124126 2816
rect 124182 2760 124187 2816
rect 123956 2758 124187 2760
rect 123956 2756 123962 2758
rect 124121 2755 124187 2758
rect 133454 2756 133460 2820
rect 133524 2818 133530 2820
rect 133781 2818 133847 2821
rect 133524 2816 133847 2818
rect 133524 2760 133786 2816
rect 133842 2760 133847 2816
rect 133524 2758 133847 2760
rect 133524 2756 133530 2758
rect 133781 2755 133847 2758
rect 140037 2818 140103 2821
rect 140865 2818 140931 2821
rect 145465 2820 145531 2821
rect 145414 2818 145420 2820
rect 140037 2816 140931 2818
rect 140037 2760 140042 2816
rect 140098 2760 140870 2816
rect 140926 2760 140931 2816
rect 140037 2758 140931 2760
rect 145374 2758 145420 2818
rect 145484 2816 145531 2820
rect 145526 2760 145531 2816
rect 140037 2755 140103 2758
rect 140865 2755 140931 2758
rect 145414 2756 145420 2758
rect 145484 2756 145531 2760
rect 147630 2818 147690 2894
rect 149094 2892 149100 2956
rect 149164 2954 149170 2956
rect 150341 2954 150407 2957
rect 149164 2952 150407 2954
rect 149164 2896 150346 2952
rect 150402 2896 150407 2952
rect 149164 2894 150407 2896
rect 149164 2892 149170 2894
rect 150341 2891 150407 2894
rect 153510 2892 153516 2956
rect 153580 2954 153586 2956
rect 153653 2954 153719 2957
rect 155033 2956 155099 2957
rect 154982 2954 154988 2956
rect 153580 2952 153719 2954
rect 153580 2896 153658 2952
rect 153714 2896 153719 2952
rect 153580 2894 153719 2896
rect 154942 2894 154988 2954
rect 155052 2952 155099 2956
rect 155094 2896 155099 2952
rect 153580 2892 153586 2894
rect 153653 2891 153719 2894
rect 154982 2892 154988 2894
rect 155052 2892 155099 2896
rect 155033 2891 155099 2892
rect 155861 2954 155927 2957
rect 157057 2954 157123 2957
rect 155861 2952 215310 2954
rect 155861 2896 155866 2952
rect 155922 2896 157062 2952
rect 157118 2896 215310 2952
rect 155861 2894 215310 2896
rect 155861 2891 155927 2894
rect 157057 2891 157123 2894
rect 154389 2818 154455 2821
rect 156413 2820 156479 2821
rect 156413 2818 156460 2820
rect 147630 2816 154455 2818
rect 147630 2760 154394 2816
rect 154450 2760 154455 2816
rect 147630 2758 154455 2760
rect 156368 2816 156460 2818
rect 156368 2760 156418 2816
rect 156368 2758 156460 2760
rect 145465 2755 145531 2756
rect 154389 2755 154455 2758
rect 156413 2756 156460 2758
rect 156524 2756 156530 2820
rect 189942 2756 189948 2820
rect 190012 2818 190018 2820
rect 190361 2818 190427 2821
rect 190012 2816 190427 2818
rect 190012 2760 190366 2816
rect 190422 2760 190427 2816
rect 190012 2758 190427 2760
rect 190012 2756 190018 2758
rect 156413 2755 156479 2756
rect 190361 2755 190427 2758
rect 191414 2756 191420 2820
rect 191484 2818 191490 2820
rect 191741 2818 191807 2821
rect 191484 2816 191807 2818
rect 191484 2760 191746 2816
rect 191802 2760 191807 2816
rect 191484 2758 191807 2760
rect 191484 2756 191490 2758
rect 191741 2755 191807 2758
rect 198038 2756 198044 2820
rect 198108 2818 198114 2820
rect 198641 2818 198707 2821
rect 198108 2816 198707 2818
rect 198108 2760 198646 2816
rect 198702 2760 198707 2816
rect 198108 2758 198707 2760
rect 198108 2756 198114 2758
rect 198641 2755 198707 2758
rect 199510 2756 199516 2820
rect 199580 2818 199586 2820
rect 200021 2818 200087 2821
rect 199580 2816 200087 2818
rect 199580 2760 200026 2816
rect 200082 2760 200087 2816
rect 199580 2758 200087 2760
rect 199580 2756 199586 2758
rect 200021 2755 200087 2758
rect 200982 2756 200988 2820
rect 201052 2818 201058 2820
rect 201401 2818 201467 2821
rect 201052 2816 201467 2818
rect 201052 2760 201406 2816
rect 201462 2760 201467 2816
rect 201052 2758 201467 2760
rect 201052 2756 201058 2758
rect 201401 2755 201467 2758
rect 209681 2818 209747 2821
rect 210734 2818 210740 2820
rect 209681 2816 210740 2818
rect 209681 2760 209686 2816
rect 209742 2760 210740 2816
rect 209681 2758 210740 2760
rect 209681 2755 209747 2758
rect 210734 2756 210740 2758
rect 210804 2756 210810 2820
rect 215250 2818 215310 2894
rect 216622 2892 216628 2956
rect 216692 2954 216698 2956
rect 217133 2954 217199 2957
rect 216692 2952 217199 2954
rect 216692 2896 217138 2952
rect 217194 2896 217199 2952
rect 216692 2894 217199 2896
rect 216692 2892 216698 2894
rect 217133 2891 217199 2894
rect 220997 2954 221063 2957
rect 224861 2954 224927 2957
rect 226190 2954 226196 2956
rect 220997 2952 224786 2954
rect 220997 2896 221002 2952
rect 221058 2896 224786 2952
rect 220997 2894 224786 2896
rect 220997 2891 221063 2894
rect 222561 2818 222627 2821
rect 215250 2816 222627 2818
rect 215250 2760 222566 2816
rect 222622 2760 222627 2816
rect 215250 2758 222627 2760
rect 222561 2755 222627 2758
rect 224350 2756 224356 2820
rect 224420 2818 224426 2820
rect 224493 2818 224559 2821
rect 224420 2816 224559 2818
rect 224420 2760 224498 2816
rect 224554 2760 224559 2816
rect 224420 2758 224559 2760
rect 224726 2818 224786 2894
rect 224861 2952 226196 2954
rect 224861 2896 224866 2952
rect 224922 2896 226196 2952
rect 224861 2894 226196 2896
rect 224861 2891 224927 2894
rect 226190 2892 226196 2894
rect 226260 2892 226266 2956
rect 244230 2954 244290 3030
rect 249057 3027 249123 3030
rect 250846 3028 250852 3092
rect 250916 3090 250922 3092
rect 250989 3090 251055 3093
rect 263550 3090 263610 3166
rect 271137 3163 271203 3166
rect 271781 3226 271847 3229
rect 271781 3224 272504 3226
rect 271781 3168 271786 3224
rect 271842 3168 272504 3224
rect 271781 3166 272504 3168
rect 271781 3163 271847 3166
rect 250916 3088 251055 3090
rect 250916 3032 250994 3088
rect 251050 3032 251055 3088
rect 250916 3030 251055 3032
rect 250916 3028 250922 3030
rect 250989 3027 251055 3030
rect 252234 3030 263610 3090
rect 267917 3090 267983 3093
rect 267917 3088 272504 3090
rect 267917 3032 267922 3088
rect 267978 3032 272504 3088
rect 267917 3030 272504 3032
rect 234570 2894 244290 2954
rect 234570 2818 234630 2894
rect 246430 2892 246436 2956
rect 246500 2954 246506 2956
rect 246849 2954 246915 2957
rect 246500 2952 246915 2954
rect 246500 2896 246854 2952
rect 246910 2896 246915 2952
rect 246500 2894 246915 2896
rect 246500 2892 246506 2894
rect 246849 2891 246915 2894
rect 250529 2954 250595 2957
rect 252234 2954 252294 3030
rect 267917 3027 267983 3030
rect 250529 2952 252294 2954
rect 250529 2896 250534 2952
rect 250590 2896 252294 2952
rect 250529 2894 252294 2896
rect 250529 2891 250595 2894
rect 255998 2892 256004 2956
rect 256068 2954 256074 2956
rect 256509 2954 256575 2957
rect 256068 2952 256575 2954
rect 256068 2896 256514 2952
rect 256570 2896 256575 2952
rect 256068 2894 256575 2896
rect 256068 2892 256074 2894
rect 256509 2891 256575 2894
rect 258766 2894 272504 2954
rect 224726 2758 234630 2818
rect 249609 2818 249675 2821
rect 258766 2818 258826 2894
rect 249609 2816 258826 2818
rect 249609 2760 249614 2816
rect 249670 2760 258826 2816
rect 249609 2758 258826 2760
rect 224420 2756 224426 2758
rect 224493 2755 224559 2758
rect 249609 2755 249675 2758
rect 259678 2756 259684 2820
rect 259748 2818 259754 2820
rect 259821 2818 259887 2821
rect 260465 2820 260531 2821
rect 260414 2818 260420 2820
rect 259748 2816 259887 2818
rect 259748 2760 259826 2816
rect 259882 2760 259887 2816
rect 259748 2758 259887 2760
rect 260374 2758 260420 2818
rect 260484 2816 260531 2820
rect 260526 2760 260531 2816
rect 259748 2756 259754 2758
rect 259821 2755 259887 2758
rect 260414 2756 260420 2758
rect 260484 2756 260531 2760
rect 261886 2756 261892 2820
rect 261956 2818 261962 2820
rect 262121 2818 262187 2821
rect 261956 2816 262187 2818
rect 261956 2760 262126 2816
rect 262182 2760 262187 2816
rect 261956 2758 262187 2760
rect 261956 2756 261962 2758
rect 260465 2755 260531 2756
rect 262121 2755 262187 2758
rect 262581 2818 262647 2821
rect 267917 2818 267983 2821
rect 262581 2816 267983 2818
rect 262581 2760 262586 2816
rect 262642 2760 267922 2816
rect 267978 2760 267983 2816
rect 262581 2758 267983 2760
rect 262581 2755 262647 2758
rect 267917 2755 267983 2758
rect 270677 2818 270743 2821
rect 271086 2818 271092 2820
rect 270677 2816 271092 2818
rect 270677 2760 270682 2816
rect 270738 2760 271092 2816
rect 270677 2758 271092 2760
rect 270677 2755 270743 2758
rect 271086 2756 271092 2758
rect 271156 2756 271162 2820
rect 271229 2818 271295 2821
rect 271229 2816 272504 2818
rect 271229 2760 271234 2816
rect 271290 2760 272504 2816
rect 271229 2758 272504 2760
rect 271229 2755 271295 2758
rect 34744 2752 35060 2753
rect 34744 2688 34750 2752
rect 34814 2688 34830 2752
rect 34894 2688 34910 2752
rect 34974 2688 34990 2752
rect 35054 2688 35060 2752
rect 34744 2687 35060 2688
rect 102341 2752 102657 2753
rect 102341 2688 102347 2752
rect 102411 2688 102427 2752
rect 102491 2688 102507 2752
rect 102571 2688 102587 2752
rect 102651 2688 102657 2752
rect 102341 2687 102657 2688
rect 169938 2752 170254 2753
rect 169938 2688 169944 2752
rect 170008 2688 170024 2752
rect 170088 2688 170104 2752
rect 170168 2688 170184 2752
rect 170248 2688 170254 2752
rect 169938 2687 170254 2688
rect 237535 2752 237851 2753
rect 237535 2688 237541 2752
rect 237605 2688 237621 2752
rect 237685 2688 237701 2752
rect 237765 2688 237781 2752
rect 237845 2688 237851 2752
rect 237535 2687 237851 2688
rect 94405 2682 94471 2685
rect 97717 2682 97783 2685
rect 120809 2682 120875 2685
rect 121085 2682 121151 2685
rect 94405 2680 97783 2682
rect 94405 2624 94410 2680
rect 94466 2624 97722 2680
rect 97778 2624 97783 2680
rect 94405 2622 97783 2624
rect 94405 2619 94471 2622
rect 97717 2619 97783 2622
rect 104206 2680 121151 2682
rect 104206 2624 120814 2680
rect 120870 2624 121090 2680
rect 121146 2624 121151 2680
rect 104206 2622 121151 2624
rect 4797 2546 4863 2549
rect 38745 2546 38811 2549
rect 4797 2544 38811 2546
rect 4797 2488 4802 2544
rect 4858 2488 38750 2544
rect 38806 2488 38811 2544
rect 4797 2486 38811 2488
rect 4797 2483 4863 2486
rect 38745 2483 38811 2486
rect 88977 2546 89043 2549
rect 104206 2546 104266 2622
rect 120809 2619 120875 2622
rect 121085 2619 121151 2622
rect 124121 2682 124187 2685
rect 156965 2682 157031 2685
rect 124121 2680 157031 2682
rect 124121 2624 124126 2680
rect 124182 2624 156970 2680
rect 157026 2624 157031 2680
rect 124121 2622 157031 2624
rect 124121 2619 124187 2622
rect 156965 2619 157031 2622
rect 219893 2682 219959 2685
rect 225413 2682 225479 2685
rect 251081 2682 251147 2685
rect 219893 2680 225479 2682
rect 219893 2624 219898 2680
rect 219954 2624 225418 2680
rect 225474 2624 225479 2680
rect 219893 2622 225479 2624
rect 219893 2619 219959 2622
rect 225413 2619 225479 2622
rect 238710 2680 251147 2682
rect 238710 2624 251086 2680
rect 251142 2624 251147 2680
rect 238710 2622 251147 2624
rect 88977 2544 104266 2546
rect 88977 2488 88982 2544
rect 89038 2488 104266 2544
rect 88977 2486 104266 2488
rect 105997 2546 106063 2549
rect 110137 2546 110203 2549
rect 105997 2544 110203 2546
rect 105997 2488 106002 2544
rect 106058 2488 110142 2544
rect 110198 2488 110203 2544
rect 105997 2486 110203 2488
rect 88977 2483 89043 2486
rect 105997 2483 106063 2486
rect 110137 2483 110203 2486
rect 110321 2546 110387 2549
rect 119429 2546 119495 2549
rect 110321 2544 119495 2546
rect 110321 2488 110326 2544
rect 110382 2488 119434 2544
rect 119490 2488 119495 2544
rect 110321 2486 119495 2488
rect 110321 2483 110387 2486
rect 119429 2483 119495 2486
rect 134149 2546 134215 2549
rect 156229 2546 156295 2549
rect 134149 2544 156295 2546
rect 134149 2488 134154 2544
rect 134210 2488 156234 2544
rect 156290 2488 156295 2544
rect 134149 2486 156295 2488
rect 134149 2483 134215 2486
rect 156229 2483 156295 2486
rect 156597 2546 156663 2549
rect 214557 2546 214623 2549
rect 156597 2544 214623 2546
rect 156597 2488 156602 2544
rect 156658 2488 214562 2544
rect 214618 2488 214623 2544
rect 156597 2486 214623 2488
rect 156597 2483 156663 2486
rect 214557 2483 214623 2486
rect 216857 2546 216923 2549
rect 221089 2546 221155 2549
rect 216857 2544 221155 2546
rect 216857 2488 216862 2544
rect 216918 2488 221094 2544
rect 221150 2488 221155 2544
rect 216857 2486 221155 2488
rect 216857 2483 216923 2486
rect 221089 2483 221155 2486
rect 223573 2546 223639 2549
rect 238710 2546 238770 2622
rect 251081 2619 251147 2622
rect 267917 2682 267983 2685
rect 267917 2680 272504 2682
rect 267917 2624 267922 2680
rect 267978 2624 272504 2680
rect 267917 2622 272504 2624
rect 267917 2619 267983 2622
rect 249701 2546 249767 2549
rect 223573 2544 238770 2546
rect 223573 2488 223578 2544
rect 223634 2488 238770 2544
rect 223573 2486 238770 2488
rect 243494 2544 249767 2546
rect 243494 2488 249706 2544
rect 249762 2488 249767 2544
rect 243494 2486 249767 2488
rect 223573 2483 223639 2486
rect 65057 2410 65123 2413
rect 91185 2410 91251 2413
rect 96429 2410 96495 2413
rect 65057 2408 80070 2410
rect 65057 2352 65062 2408
rect 65118 2352 80070 2408
rect 65057 2350 80070 2352
rect 65057 2347 65123 2350
rect 80010 2274 80070 2350
rect 91185 2408 96495 2410
rect 91185 2352 91190 2408
rect 91246 2352 96434 2408
rect 96490 2352 96495 2408
rect 91185 2350 96495 2352
rect 91185 2347 91251 2350
rect 96429 2347 96495 2350
rect 96654 2348 96660 2412
rect 96724 2410 96730 2412
rect 96889 2410 96955 2413
rect 96724 2408 96955 2410
rect 96724 2352 96894 2408
rect 96950 2352 96955 2408
rect 96724 2350 96955 2352
rect 96724 2348 96730 2350
rect 96889 2347 96955 2350
rect 101305 2410 101371 2413
rect 146293 2410 146359 2413
rect 151721 2412 151787 2413
rect 151670 2410 151676 2412
rect 101305 2408 147690 2410
rect 101305 2352 101310 2408
rect 101366 2352 146298 2408
rect 146354 2352 147690 2408
rect 101305 2350 147690 2352
rect 151630 2350 151676 2410
rect 151740 2408 151787 2412
rect 214373 2410 214439 2413
rect 151782 2352 151787 2408
rect 101305 2347 101371 2350
rect 146293 2347 146359 2350
rect 93669 2274 93735 2277
rect 95969 2274 96035 2277
rect 80010 2272 93735 2274
rect 80010 2216 93674 2272
rect 93730 2216 93735 2272
rect 80010 2214 93735 2216
rect 93669 2211 93735 2214
rect 93902 2272 96035 2274
rect 93902 2216 95974 2272
rect 96030 2216 96035 2272
rect 93902 2214 96035 2216
rect 68542 2208 68858 2209
rect 68542 2144 68548 2208
rect 68612 2144 68628 2208
rect 68692 2144 68708 2208
rect 68772 2144 68788 2208
rect 68852 2144 68858 2208
rect 68542 2143 68858 2144
rect 23105 2138 23171 2141
rect 53281 2138 53347 2141
rect 23105 2136 53347 2138
rect 23105 2080 23110 2136
rect 23166 2080 53286 2136
rect 53342 2080 53347 2136
rect 23105 2078 53347 2080
rect 23105 2075 23171 2078
rect 53281 2075 53347 2078
rect 89621 2138 89687 2141
rect 93902 2138 93962 2214
rect 95969 2211 96035 2214
rect 96110 2214 109050 2274
rect 94221 2140 94287 2141
rect 94221 2138 94268 2140
rect 89621 2136 93962 2138
rect 89621 2080 89626 2136
rect 89682 2080 93962 2136
rect 89621 2078 93962 2080
rect 94176 2136 94268 2138
rect 94176 2080 94226 2136
rect 94176 2078 94268 2080
rect 89621 2075 89687 2078
rect 94221 2076 94268 2078
rect 94332 2076 94338 2140
rect 95325 2138 95391 2141
rect 96110 2138 96170 2214
rect 96429 2140 96495 2141
rect 96429 2138 96476 2140
rect 95325 2136 96170 2138
rect 95325 2080 95330 2136
rect 95386 2080 96170 2136
rect 95325 2078 96170 2080
rect 96384 2136 96476 2138
rect 96384 2080 96434 2136
rect 96384 2078 96476 2080
rect 94221 2075 94287 2076
rect 95325 2075 95391 2078
rect 96429 2076 96476 2078
rect 96540 2076 96546 2140
rect 97809 2138 97875 2141
rect 104065 2138 104131 2141
rect 97809 2136 104131 2138
rect 97809 2080 97814 2136
rect 97870 2080 104070 2136
rect 104126 2080 104131 2136
rect 97809 2078 104131 2080
rect 108990 2138 109050 2214
rect 114318 2212 114324 2276
rect 114388 2274 114394 2276
rect 114553 2274 114619 2277
rect 114388 2272 114619 2274
rect 114388 2216 114558 2272
rect 114614 2216 114619 2272
rect 114388 2214 114619 2216
rect 147630 2274 147690 2350
rect 151670 2348 151676 2350
rect 151740 2348 151787 2352
rect 151721 2347 151787 2348
rect 151862 2408 214439 2410
rect 151862 2352 214378 2408
rect 214434 2352 214439 2408
rect 151862 2350 214439 2352
rect 151862 2274 151922 2350
rect 214373 2347 214439 2350
rect 215937 2410 216003 2413
rect 227069 2410 227135 2413
rect 215937 2408 227135 2410
rect 215937 2352 215942 2408
rect 215998 2352 227074 2408
rect 227130 2352 227135 2408
rect 215937 2350 227135 2352
rect 215937 2347 216003 2350
rect 227069 2347 227135 2350
rect 227897 2410 227963 2413
rect 243494 2410 243554 2486
rect 249701 2483 249767 2486
rect 268377 2546 268443 2549
rect 268377 2544 272504 2546
rect 268377 2488 268382 2544
rect 268438 2488 272504 2544
rect 268377 2486 272504 2488
rect 268377 2483 268443 2486
rect 227897 2408 243554 2410
rect 227897 2352 227902 2408
rect 227958 2352 243554 2408
rect 227897 2350 243554 2352
rect 248413 2410 248479 2413
rect 248413 2408 272504 2410
rect 248413 2352 248418 2408
rect 248474 2352 272504 2408
rect 248413 2350 272504 2352
rect 227897 2347 227963 2350
rect 248413 2347 248479 2350
rect 147630 2214 151922 2274
rect 154389 2274 154455 2277
rect 176837 2274 176903 2277
rect 154389 2272 176903 2274
rect 154389 2216 154394 2272
rect 154450 2216 176842 2272
rect 176898 2216 176903 2272
rect 154389 2214 176903 2216
rect 114388 2212 114394 2214
rect 114553 2211 114619 2214
rect 154389 2211 154455 2214
rect 176837 2211 176903 2214
rect 213637 2274 213703 2277
rect 245009 2274 245075 2277
rect 247401 2274 247467 2277
rect 213637 2272 245075 2274
rect 213637 2216 213642 2272
rect 213698 2216 245014 2272
rect 245070 2216 245075 2272
rect 213637 2214 245075 2216
rect 213637 2211 213703 2214
rect 245009 2211 245075 2214
rect 245334 2272 247467 2274
rect 245334 2216 247406 2272
rect 247462 2216 247467 2272
rect 245334 2214 247467 2216
rect 136139 2208 136455 2209
rect 136139 2144 136145 2208
rect 136209 2144 136225 2208
rect 136289 2144 136305 2208
rect 136369 2144 136385 2208
rect 136449 2144 136455 2208
rect 136139 2143 136455 2144
rect 203736 2208 204052 2209
rect 203736 2144 203742 2208
rect 203806 2144 203822 2208
rect 203886 2144 203902 2208
rect 203966 2144 203982 2208
rect 204046 2144 204052 2208
rect 203736 2143 204052 2144
rect 123477 2138 123543 2141
rect 124121 2138 124187 2141
rect 108990 2136 124187 2138
rect 108990 2080 123482 2136
rect 123538 2080 124126 2136
rect 124182 2080 124187 2136
rect 108990 2078 124187 2080
rect 96429 2075 96495 2076
rect 97809 2075 97875 2078
rect 104065 2075 104131 2078
rect 123477 2075 123543 2078
rect 124121 2075 124187 2078
rect 147581 2138 147647 2141
rect 151261 2138 151327 2141
rect 179413 2138 179479 2141
rect 147581 2136 151327 2138
rect 147581 2080 147586 2136
rect 147642 2080 151266 2136
rect 151322 2080 151327 2136
rect 147581 2078 151327 2080
rect 147581 2075 147647 2078
rect 151261 2075 151327 2078
rect 157290 2136 179479 2138
rect 157290 2080 179418 2136
rect 179474 2080 179479 2136
rect 157290 2078 179479 2080
rect 8661 2002 8727 2005
rect 43345 2002 43411 2005
rect 8661 2000 43411 2002
rect 8661 1944 8666 2000
rect 8722 1944 43350 2000
rect 43406 1944 43411 2000
rect 8661 1942 43411 1944
rect 8661 1939 8727 1942
rect 43345 1939 43411 1942
rect 84837 2002 84903 2005
rect 117681 2002 117747 2005
rect 149605 2002 149671 2005
rect 84837 2000 117747 2002
rect 84837 1944 84842 2000
rect 84898 1944 117686 2000
rect 117742 1944 117747 2000
rect 84837 1942 117747 1944
rect 84837 1939 84903 1942
rect 117681 1939 117747 1942
rect 122790 2000 149671 2002
rect 122790 1944 149610 2000
rect 149666 1944 149671 2000
rect 122790 1942 149671 1944
rect 72049 1866 72115 1869
rect 74625 1866 74691 1869
rect 93669 1866 93735 1869
rect 95049 1866 95115 1869
rect 72049 1864 74691 1866
rect 72049 1808 72054 1864
rect 72110 1808 74630 1864
rect 74686 1808 74691 1864
rect 72049 1806 74691 1808
rect 72049 1803 72115 1806
rect 74625 1803 74691 1806
rect 80010 1806 92674 1866
rect 22001 1730 22067 1733
rect 22134 1730 22140 1732
rect 22001 1728 22140 1730
rect 22001 1672 22006 1728
rect 22062 1672 22140 1728
rect 22001 1670 22140 1672
rect 22001 1667 22067 1670
rect 22134 1668 22140 1670
rect 22204 1668 22210 1732
rect 40401 1730 40467 1733
rect 80010 1730 80070 1806
rect 92381 1730 92447 1733
rect 40401 1728 80070 1730
rect 40401 1672 40406 1728
rect 40462 1672 80070 1728
rect 40401 1670 80070 1672
rect 90958 1728 92447 1730
rect 90958 1672 92386 1728
rect 92442 1672 92447 1728
rect 90958 1670 92447 1672
rect 92614 1730 92674 1806
rect 93669 1864 95115 1866
rect 93669 1808 93674 1864
rect 93730 1808 95054 1864
rect 95110 1808 95115 1864
rect 93669 1806 95115 1808
rect 93669 1803 93735 1806
rect 95049 1803 95115 1806
rect 95233 1866 95299 1869
rect 105077 1866 105143 1869
rect 121821 1866 121887 1869
rect 122097 1866 122163 1869
rect 122790 1866 122850 1942
rect 149605 1939 149671 1942
rect 149973 2002 150039 2005
rect 157290 2002 157350 2078
rect 179413 2075 179479 2078
rect 216029 2138 216095 2141
rect 245334 2138 245394 2214
rect 247401 2211 247467 2214
rect 254117 2274 254183 2277
rect 271137 2274 271203 2277
rect 254117 2272 271203 2274
rect 254117 2216 254122 2272
rect 254178 2216 271142 2272
rect 271198 2216 271203 2272
rect 254117 2214 271203 2216
rect 254117 2211 254183 2214
rect 271137 2211 271203 2214
rect 271830 2214 272504 2274
rect 271333 2208 271649 2209
rect 271333 2144 271339 2208
rect 271403 2144 271419 2208
rect 271483 2144 271499 2208
rect 271563 2144 271579 2208
rect 271643 2144 271649 2208
rect 271333 2143 271649 2144
rect 260281 2138 260347 2141
rect 216029 2136 245394 2138
rect 216029 2080 216034 2136
rect 216090 2080 245394 2136
rect 216029 2078 245394 2080
rect 245610 2136 260347 2138
rect 245610 2080 260286 2136
rect 260342 2080 260347 2136
rect 245610 2078 260347 2080
rect 216029 2075 216095 2078
rect 149973 2000 157350 2002
rect 149973 1944 149978 2000
rect 150034 1944 157350 2000
rect 149973 1942 157350 1944
rect 191833 2002 191899 2005
rect 192109 2002 192175 2005
rect 219893 2002 219959 2005
rect 191833 2000 219959 2002
rect 191833 1944 191838 2000
rect 191894 1944 192114 2000
rect 192170 1944 219898 2000
rect 219954 1944 219959 2000
rect 191833 1942 219959 1944
rect 149973 1939 150039 1942
rect 191833 1939 191899 1942
rect 192109 1939 192175 1942
rect 219893 1939 219959 1942
rect 220077 2002 220143 2005
rect 224861 2002 224927 2005
rect 220077 2000 224927 2002
rect 220077 1944 220082 2000
rect 220138 1944 224866 2000
rect 224922 1944 224927 2000
rect 220077 1942 224927 1944
rect 220077 1939 220143 1942
rect 224861 1939 224927 1942
rect 226425 2002 226491 2005
rect 245610 2002 245670 2078
rect 260281 2075 260347 2078
rect 267590 2076 267596 2140
rect 267660 2138 267666 2140
rect 267733 2138 267799 2141
rect 267660 2136 267799 2138
rect 267660 2080 267738 2136
rect 267794 2080 267799 2136
rect 267660 2078 267799 2080
rect 267660 2076 267666 2078
rect 267733 2075 267799 2078
rect 226425 2000 245670 2002
rect 226425 1944 226430 2000
rect 226486 1944 245670 2000
rect 226425 1942 245670 1944
rect 250805 2002 250871 2005
rect 258717 2002 258783 2005
rect 271830 2002 271890 2214
rect 271965 2138 272031 2141
rect 271965 2136 272504 2138
rect 271965 2080 271970 2136
rect 272026 2080 272504 2136
rect 271965 2078 272504 2080
rect 271965 2075 272031 2078
rect 250805 2000 258783 2002
rect 250805 1944 250810 2000
rect 250866 1944 258722 2000
rect 258778 1944 258783 2000
rect 250805 1942 258783 1944
rect 226425 1939 226491 1942
rect 250805 1939 250871 1942
rect 258717 1939 258783 1942
rect 263550 1942 271890 2002
rect 272057 2002 272123 2005
rect 272057 2000 272504 2002
rect 272057 1944 272062 2000
rect 272118 1944 272504 2000
rect 272057 1942 272504 1944
rect 95233 1864 105143 1866
rect 95233 1808 95238 1864
rect 95294 1808 105082 1864
rect 105138 1808 105143 1864
rect 95233 1806 105143 1808
rect 95233 1803 95299 1806
rect 105077 1803 105143 1806
rect 108990 1864 122850 1866
rect 108990 1808 121826 1864
rect 121882 1808 122102 1864
rect 122158 1808 122850 1864
rect 108990 1806 122850 1808
rect 140221 1868 140287 1869
rect 140221 1864 140268 1868
rect 140332 1866 140338 1868
rect 141601 1866 141667 1869
rect 174721 1866 174787 1869
rect 140221 1808 140226 1864
rect 96797 1730 96863 1733
rect 92614 1728 96863 1730
rect 92614 1672 96802 1728
rect 96858 1672 96863 1728
rect 92614 1670 96863 1672
rect 40401 1667 40467 1670
rect 34744 1664 35060 1665
rect 34744 1600 34750 1664
rect 34814 1600 34830 1664
rect 34894 1600 34910 1664
rect 34974 1600 34990 1664
rect 35054 1600 35060 1664
rect 34744 1599 35060 1600
rect 19926 1532 19932 1596
rect 19996 1594 20002 1596
rect 20713 1594 20779 1597
rect 19996 1592 20779 1594
rect 19996 1536 20718 1592
rect 20774 1536 20779 1592
rect 19996 1534 20779 1536
rect 19996 1532 20002 1534
rect 20713 1531 20779 1534
rect 32438 1532 32444 1596
rect 32508 1594 32514 1596
rect 33133 1594 33199 1597
rect 32508 1592 33199 1594
rect 32508 1536 33138 1592
rect 33194 1536 33199 1592
rect 32508 1534 33199 1536
rect 32508 1532 32514 1534
rect 33133 1531 33199 1534
rect 57830 1532 57836 1596
rect 57900 1594 57906 1596
rect 57973 1594 58039 1597
rect 59353 1596 59419 1597
rect 59302 1594 59308 1596
rect 57900 1592 58039 1594
rect 57900 1536 57978 1592
rect 58034 1536 58039 1592
rect 57900 1534 58039 1536
rect 59262 1534 59308 1594
rect 59372 1592 59419 1596
rect 59414 1536 59419 1592
rect 57900 1532 57906 1534
rect 57973 1531 58039 1534
rect 59302 1532 59308 1534
rect 59372 1532 59419 1536
rect 59353 1531 59419 1532
rect 59537 1594 59603 1597
rect 90958 1594 91018 1670
rect 92381 1667 92447 1670
rect 96797 1667 96863 1670
rect 96981 1730 97047 1733
rect 97993 1730 98059 1733
rect 100845 1730 100911 1733
rect 96981 1728 100911 1730
rect 96981 1672 96986 1728
rect 97042 1672 97998 1728
rect 98054 1672 100850 1728
rect 100906 1672 100911 1728
rect 96981 1670 100911 1672
rect 96981 1667 97047 1670
rect 97993 1667 98059 1670
rect 100845 1667 100911 1670
rect 102341 1664 102657 1665
rect 102341 1600 102347 1664
rect 102411 1600 102427 1664
rect 102491 1600 102507 1664
rect 102571 1600 102587 1664
rect 102651 1600 102657 1664
rect 102341 1599 102657 1600
rect 91185 1596 91251 1597
rect 91134 1594 91140 1596
rect 59537 1592 91018 1594
rect 59537 1536 59542 1592
rect 59598 1536 91018 1592
rect 59537 1534 91018 1536
rect 91094 1534 91140 1594
rect 91204 1592 91251 1596
rect 91246 1536 91251 1592
rect 59537 1531 59603 1534
rect 91134 1532 91140 1534
rect 91204 1532 91251 1536
rect 91185 1531 91251 1532
rect 91369 1594 91435 1597
rect 95325 1594 95391 1597
rect 91369 1592 95391 1594
rect 91369 1536 91374 1592
rect 91430 1536 95330 1592
rect 95386 1536 95391 1592
rect 91369 1534 95391 1536
rect 91369 1531 91435 1534
rect 95325 1531 95391 1534
rect 96245 1596 96311 1597
rect 96245 1592 96292 1596
rect 96356 1594 96362 1596
rect 97901 1594 97967 1597
rect 98494 1594 98500 1596
rect 96245 1536 96250 1592
rect 96245 1532 96292 1536
rect 96356 1534 96402 1594
rect 97901 1592 98500 1594
rect 97901 1536 97906 1592
rect 97962 1536 98500 1592
rect 97901 1534 98500 1536
rect 96356 1532 96362 1534
rect 96245 1531 96311 1532
rect 97901 1531 97967 1534
rect 98494 1532 98500 1534
rect 98564 1532 98570 1596
rect 20662 1396 20668 1460
rect 20732 1458 20738 1460
rect 22369 1458 22435 1461
rect 20732 1456 22435 1458
rect 20732 1400 22374 1456
rect 22430 1400 22435 1456
rect 20732 1398 22435 1400
rect 20732 1396 20738 1398
rect 22369 1395 22435 1398
rect 23749 1458 23815 1461
rect 54293 1458 54359 1461
rect 23749 1456 88074 1458
rect 23749 1400 23754 1456
rect 23810 1400 54298 1456
rect 54354 1400 88074 1456
rect 23749 1398 88074 1400
rect 23749 1395 23815 1398
rect 54293 1395 54359 1398
rect 4521 1324 4587 1325
rect 6729 1324 6795 1325
rect 14825 1324 14891 1325
rect 4470 1322 4476 1324
rect 4430 1262 4476 1322
rect 4540 1320 4587 1324
rect 6678 1322 6684 1324
rect 4582 1264 4587 1320
rect 4470 1260 4476 1262
rect 4540 1260 4587 1264
rect 6638 1262 6684 1322
rect 6748 1320 6795 1324
rect 14774 1322 14780 1324
rect 6790 1264 6795 1320
rect 6678 1260 6684 1262
rect 6748 1260 6795 1264
rect 14734 1262 14780 1322
rect 14844 1320 14891 1324
rect 14886 1264 14891 1320
rect 14774 1260 14780 1262
rect 14844 1260 14891 1264
rect 4521 1259 4587 1260
rect 6729 1259 6795 1260
rect 14825 1259 14891 1260
rect 23565 1324 23631 1325
rect 23565 1320 23612 1324
rect 23676 1322 23682 1324
rect 23841 1322 23907 1325
rect 25773 1324 25839 1325
rect 26509 1324 26575 1325
rect 76465 1324 76531 1325
rect 78673 1324 78739 1325
rect 81617 1324 81683 1325
rect 83825 1324 83891 1325
rect 24342 1322 24348 1324
rect 23565 1264 23570 1320
rect 23565 1260 23612 1264
rect 23676 1262 23722 1322
rect 23841 1320 24348 1322
rect 23841 1264 23846 1320
rect 23902 1264 24348 1320
rect 23841 1262 24348 1264
rect 23676 1260 23682 1262
rect 23565 1259 23631 1260
rect 23841 1259 23907 1262
rect 24342 1260 24348 1262
rect 24412 1260 24418 1324
rect 25773 1320 25820 1324
rect 25884 1322 25890 1324
rect 25773 1264 25778 1320
rect 25773 1260 25820 1264
rect 25884 1262 25930 1322
rect 26509 1320 26556 1324
rect 26620 1322 26626 1324
rect 76414 1322 76420 1324
rect 26509 1264 26514 1320
rect 25884 1260 25890 1262
rect 26509 1260 26556 1264
rect 26620 1262 26666 1322
rect 76374 1262 76420 1322
rect 76484 1320 76531 1324
rect 78622 1322 78628 1324
rect 76526 1264 76531 1320
rect 26620 1260 26626 1262
rect 76414 1260 76420 1262
rect 76484 1260 76531 1264
rect 78582 1262 78628 1322
rect 78692 1320 78739 1324
rect 81566 1322 81572 1324
rect 78734 1264 78739 1320
rect 78622 1260 78628 1262
rect 78692 1260 78739 1264
rect 81526 1262 81572 1322
rect 81636 1320 81683 1324
rect 83774 1322 83780 1324
rect 81678 1264 81683 1320
rect 81566 1260 81572 1262
rect 81636 1260 81683 1264
rect 83734 1262 83780 1322
rect 83844 1320 83891 1324
rect 83886 1264 83891 1320
rect 83774 1260 83780 1262
rect 83844 1260 83891 1264
rect 88014 1322 88074 1398
rect 88190 1396 88196 1460
rect 88260 1458 88266 1460
rect 88333 1458 88399 1461
rect 89069 1458 89135 1461
rect 108990 1458 109050 1806
rect 121821 1803 121887 1806
rect 122097 1803 122163 1806
rect 140221 1804 140268 1808
rect 140332 1806 140378 1866
rect 141601 1864 174787 1866
rect 141601 1808 141606 1864
rect 141662 1808 174726 1864
rect 174782 1808 174787 1864
rect 141601 1806 174787 1808
rect 140332 1804 140338 1806
rect 140221 1803 140287 1804
rect 141601 1803 141667 1806
rect 174721 1803 174787 1806
rect 194358 1804 194364 1868
rect 194428 1866 194434 1868
rect 194593 1866 194659 1869
rect 194428 1864 194659 1866
rect 194428 1808 194598 1864
rect 194654 1808 194659 1864
rect 194428 1806 194659 1808
rect 194428 1804 194434 1806
rect 194593 1803 194659 1806
rect 195830 1804 195836 1868
rect 195900 1866 195906 1868
rect 196065 1866 196131 1869
rect 195900 1864 196131 1866
rect 195900 1808 196070 1864
rect 196126 1808 196131 1864
rect 195900 1806 196131 1808
rect 195900 1804 195906 1806
rect 196065 1803 196131 1806
rect 212206 1804 212212 1868
rect 212276 1866 212282 1868
rect 214005 1866 214071 1869
rect 212276 1864 214071 1866
rect 212276 1808 214010 1864
rect 214066 1808 214071 1864
rect 212276 1806 214071 1808
rect 212276 1804 212282 1806
rect 214005 1803 214071 1806
rect 216121 1866 216187 1869
rect 216397 1866 216463 1869
rect 218881 1866 218947 1869
rect 216121 1864 218947 1866
rect 216121 1808 216126 1864
rect 216182 1808 216402 1864
rect 216458 1808 218886 1864
rect 218942 1808 218947 1864
rect 216121 1806 218947 1808
rect 216121 1803 216187 1806
rect 216397 1803 216463 1806
rect 218881 1803 218947 1806
rect 219341 1866 219407 1869
rect 251265 1866 251331 1869
rect 219341 1864 251331 1866
rect 219341 1808 219346 1864
rect 219402 1808 251270 1864
rect 251326 1808 251331 1864
rect 219341 1806 251331 1808
rect 219341 1803 219407 1806
rect 251265 1803 251331 1806
rect 146845 1730 146911 1733
rect 149329 1730 149395 1733
rect 146845 1728 149395 1730
rect 146845 1672 146850 1728
rect 146906 1672 149334 1728
rect 149390 1672 149395 1728
rect 146845 1670 149395 1672
rect 146845 1667 146911 1670
rect 149329 1667 149395 1670
rect 149605 1730 149671 1733
rect 156597 1730 156663 1733
rect 149605 1728 156663 1730
rect 149605 1672 149610 1728
rect 149666 1672 156602 1728
rect 156658 1672 156663 1728
rect 149605 1670 156663 1672
rect 149605 1667 149671 1670
rect 156597 1667 156663 1670
rect 156781 1730 156847 1733
rect 162945 1730 163011 1733
rect 156781 1728 163011 1730
rect 156781 1672 156786 1728
rect 156842 1672 162950 1728
rect 163006 1672 163011 1728
rect 156781 1670 163011 1672
rect 156781 1667 156847 1670
rect 162945 1667 163011 1670
rect 214557 1730 214623 1733
rect 220077 1730 220143 1733
rect 214557 1728 220143 1730
rect 214557 1672 214562 1728
rect 214618 1672 220082 1728
rect 220138 1672 220143 1728
rect 214557 1670 220143 1672
rect 214557 1667 214623 1670
rect 220077 1667 220143 1670
rect 221733 1730 221799 1733
rect 226517 1730 226583 1733
rect 230381 1730 230447 1733
rect 221733 1728 226583 1730
rect 221733 1672 221738 1728
rect 221794 1672 226522 1728
rect 226578 1672 226583 1728
rect 221733 1670 226583 1672
rect 221733 1667 221799 1670
rect 226517 1667 226583 1670
rect 229050 1728 230447 1730
rect 229050 1672 230386 1728
rect 230442 1672 230447 1728
rect 229050 1670 230447 1672
rect 169938 1664 170254 1665
rect 169938 1600 169944 1664
rect 170008 1600 170024 1664
rect 170088 1600 170104 1664
rect 170168 1600 170184 1664
rect 170248 1600 170254 1664
rect 169938 1599 170254 1600
rect 150249 1594 150315 1597
rect 153101 1594 153167 1597
rect 150249 1592 153167 1594
rect 150249 1536 150254 1592
rect 150310 1536 153106 1592
rect 153162 1536 153167 1592
rect 150249 1534 153167 1536
rect 150249 1531 150315 1534
rect 153101 1531 153167 1534
rect 208577 1594 208643 1597
rect 229050 1594 229110 1670
rect 230381 1667 230447 1670
rect 246665 1730 246731 1733
rect 263550 1730 263610 1942
rect 272057 1939 272123 1942
rect 268837 1866 268903 1869
rect 268837 1864 272504 1866
rect 268837 1808 268842 1864
rect 268898 1808 272504 1864
rect 268837 1806 272504 1808
rect 268837 1803 268903 1806
rect 246665 1728 263610 1730
rect 246665 1672 246670 1728
rect 246726 1672 263610 1728
rect 246665 1670 263610 1672
rect 269622 1670 272504 1730
rect 246665 1667 246731 1670
rect 237535 1664 237851 1665
rect 237535 1600 237541 1664
rect 237605 1600 237621 1664
rect 237685 1600 237701 1664
rect 237765 1600 237781 1664
rect 237845 1600 237851 1664
rect 237535 1599 237851 1600
rect 208577 1592 229110 1594
rect 208577 1536 208582 1592
rect 208638 1536 229110 1592
rect 208577 1534 229110 1536
rect 208577 1531 208643 1534
rect 237230 1532 237236 1596
rect 237300 1594 237306 1596
rect 237373 1594 237439 1597
rect 246941 1594 247007 1597
rect 237300 1592 237439 1594
rect 237300 1536 237378 1592
rect 237434 1536 237439 1592
rect 237300 1534 237439 1536
rect 237300 1532 237306 1534
rect 237373 1531 237439 1534
rect 238710 1592 247007 1594
rect 238710 1536 246946 1592
rect 247002 1536 247007 1592
rect 238710 1534 247007 1536
rect 88260 1456 88399 1458
rect 88260 1400 88338 1456
rect 88394 1400 88399 1456
rect 88260 1398 88399 1400
rect 88260 1396 88266 1398
rect 88333 1395 88399 1398
rect 88566 1456 109050 1458
rect 88566 1400 89074 1456
rect 89130 1400 109050 1456
rect 88566 1398 109050 1400
rect 109217 1458 109283 1461
rect 111333 1458 111399 1461
rect 109217 1456 111399 1458
rect 109217 1400 109222 1456
rect 109278 1400 111338 1456
rect 111394 1400 111399 1456
rect 109217 1398 111399 1400
rect 88566 1322 88626 1398
rect 89069 1395 89135 1398
rect 109217 1395 109283 1398
rect 111333 1395 111399 1398
rect 113582 1396 113588 1460
rect 113652 1458 113658 1460
rect 114553 1458 114619 1461
rect 113652 1456 114619 1458
rect 113652 1400 114558 1456
rect 114614 1400 114619 1456
rect 113652 1398 114619 1400
rect 113652 1396 113658 1398
rect 114553 1395 114619 1398
rect 114829 1460 114895 1461
rect 115565 1460 115631 1461
rect 117313 1460 117379 1461
rect 114829 1456 114876 1460
rect 114940 1458 114946 1460
rect 114829 1400 114834 1456
rect 114829 1396 114876 1400
rect 114940 1398 114986 1458
rect 115565 1456 115612 1460
rect 115676 1458 115682 1460
rect 117262 1458 117268 1460
rect 115565 1400 115570 1456
rect 114940 1396 114946 1398
rect 115565 1396 115612 1400
rect 115676 1398 115722 1458
rect 117222 1398 117268 1458
rect 117332 1456 117379 1460
rect 117374 1400 117379 1456
rect 115676 1396 115682 1398
rect 117262 1396 117268 1398
rect 117332 1396 117379 1400
rect 126830 1396 126836 1460
rect 126900 1458 126906 1460
rect 126973 1458 127039 1461
rect 126900 1456 127039 1458
rect 126900 1400 126978 1456
rect 127034 1400 127039 1456
rect 126900 1398 127039 1400
rect 126900 1396 126906 1398
rect 114829 1395 114895 1396
rect 115565 1395 115631 1396
rect 117313 1395 117379 1396
rect 126973 1395 127039 1398
rect 128302 1396 128308 1460
rect 128372 1458 128378 1460
rect 128445 1458 128511 1461
rect 128372 1456 128511 1458
rect 128372 1400 128450 1456
rect 128506 1400 128511 1456
rect 128372 1398 128511 1400
rect 128372 1396 128378 1398
rect 128445 1395 128511 1398
rect 134926 1396 134932 1460
rect 134996 1458 135002 1460
rect 135253 1458 135319 1461
rect 134996 1456 135319 1458
rect 134996 1400 135258 1456
rect 135314 1400 135319 1456
rect 134996 1398 135319 1400
rect 134996 1396 135002 1398
rect 135253 1395 135319 1398
rect 137318 1396 137324 1460
rect 137388 1458 137394 1460
rect 138013 1458 138079 1461
rect 137388 1456 138079 1458
rect 137388 1400 138018 1456
rect 138074 1400 138079 1456
rect 137388 1398 138079 1400
rect 137388 1396 137394 1398
rect 138013 1395 138079 1398
rect 140681 1458 140747 1461
rect 150617 1460 150683 1461
rect 152089 1460 152155 1461
rect 140998 1458 141004 1460
rect 140681 1456 141004 1458
rect 140681 1400 140686 1456
rect 140742 1400 141004 1456
rect 140681 1398 141004 1400
rect 140681 1395 140747 1398
rect 140998 1396 141004 1398
rect 141068 1396 141074 1460
rect 150566 1458 150572 1460
rect 150526 1398 150572 1458
rect 150636 1456 150683 1460
rect 152038 1458 152044 1460
rect 150678 1400 150683 1456
rect 150566 1396 150572 1398
rect 150636 1396 150683 1400
rect 151998 1398 152044 1458
rect 152108 1456 152155 1460
rect 152150 1400 152155 1456
rect 152038 1396 152044 1398
rect 152108 1396 152155 1400
rect 155718 1396 155724 1460
rect 155788 1458 155794 1460
rect 155953 1458 156019 1461
rect 157241 1460 157307 1461
rect 157190 1458 157196 1460
rect 155788 1456 156019 1458
rect 155788 1400 155958 1456
rect 156014 1400 156019 1456
rect 155788 1398 156019 1400
rect 157150 1398 157196 1458
rect 157260 1456 157307 1460
rect 157302 1400 157307 1456
rect 155788 1396 155794 1398
rect 150617 1395 150683 1396
rect 152089 1395 152155 1396
rect 155953 1395 156019 1398
rect 157190 1396 157196 1398
rect 157260 1396 157307 1400
rect 168230 1396 168236 1460
rect 168300 1458 168306 1460
rect 168373 1458 168439 1461
rect 186313 1460 186379 1461
rect 197353 1460 197419 1461
rect 186262 1458 186268 1460
rect 168300 1456 168439 1458
rect 168300 1400 168378 1456
rect 168434 1400 168439 1456
rect 168300 1398 168439 1400
rect 186222 1398 186268 1458
rect 186332 1456 186379 1460
rect 197302 1458 197308 1460
rect 186374 1400 186379 1456
rect 168300 1396 168306 1398
rect 157241 1395 157307 1396
rect 168373 1395 168439 1398
rect 186262 1396 186268 1398
rect 186332 1396 186379 1400
rect 197262 1398 197308 1458
rect 197372 1456 197419 1460
rect 197414 1400 197419 1456
rect 197302 1396 197308 1398
rect 197372 1396 197419 1400
rect 201718 1396 201724 1460
rect 201788 1458 201794 1460
rect 202873 1458 202939 1461
rect 201788 1456 202939 1458
rect 201788 1400 202878 1456
rect 202934 1400 202939 1456
rect 201788 1398 202939 1400
rect 201788 1396 201794 1398
rect 186313 1395 186379 1396
rect 197353 1395 197419 1396
rect 202873 1395 202939 1398
rect 209681 1458 209747 1461
rect 209998 1458 210004 1460
rect 209681 1456 210004 1458
rect 209681 1400 209686 1456
rect 209742 1400 210004 1456
rect 209681 1398 210004 1400
rect 209681 1395 209747 1398
rect 209998 1396 210004 1398
rect 210068 1396 210074 1460
rect 218094 1396 218100 1460
rect 218164 1458 218170 1460
rect 218329 1458 218395 1461
rect 218164 1456 218395 1458
rect 218164 1400 218334 1456
rect 218390 1400 218395 1456
rect 218164 1398 218395 1400
rect 218164 1396 218170 1398
rect 218329 1395 218395 1398
rect 219566 1396 219572 1460
rect 219636 1458 219642 1460
rect 219709 1458 219775 1461
rect 222561 1460 222627 1461
rect 222510 1458 222516 1460
rect 219636 1456 219775 1458
rect 219636 1400 219714 1456
rect 219770 1400 219775 1456
rect 219636 1398 219775 1400
rect 222470 1398 222516 1458
rect 222580 1456 222627 1460
rect 222622 1400 222627 1456
rect 219636 1396 219642 1398
rect 219709 1395 219775 1398
rect 222510 1396 222516 1398
rect 222580 1396 222627 1400
rect 226190 1396 226196 1460
rect 226260 1458 226266 1460
rect 226333 1458 226399 1461
rect 226260 1456 226399 1458
rect 226260 1400 226338 1456
rect 226394 1400 226399 1456
rect 226260 1398 226399 1400
rect 226260 1396 226266 1398
rect 222561 1395 222627 1396
rect 226333 1395 226399 1398
rect 226517 1458 226583 1461
rect 238710 1458 238770 1534
rect 246941 1531 247007 1534
rect 249374 1532 249380 1596
rect 249444 1594 249450 1596
rect 251357 1594 251423 1597
rect 249444 1592 251423 1594
rect 249444 1536 251362 1592
rect 251418 1536 251423 1592
rect 249444 1534 251423 1536
rect 249444 1532 249450 1534
rect 251357 1531 251423 1534
rect 251582 1532 251588 1596
rect 251652 1594 251658 1596
rect 252553 1594 252619 1597
rect 251652 1592 252619 1594
rect 251652 1536 252558 1592
rect 252614 1536 252619 1592
rect 251652 1534 252619 1536
rect 251652 1532 251658 1534
rect 252553 1531 252619 1534
rect 256734 1532 256740 1596
rect 256804 1594 256810 1596
rect 258165 1594 258231 1597
rect 269622 1594 269682 1670
rect 256804 1592 258231 1594
rect 256804 1536 258170 1592
rect 258226 1536 258231 1592
rect 256804 1534 258231 1536
rect 256804 1532 256810 1534
rect 258165 1531 258231 1534
rect 258398 1534 269682 1594
rect 269849 1594 269915 1597
rect 271965 1594 272031 1597
rect 269849 1592 272031 1594
rect 269849 1536 269854 1592
rect 269910 1536 271970 1592
rect 272026 1536 272031 1592
rect 269849 1534 272031 1536
rect 242801 1460 242867 1461
rect 245745 1460 245811 1461
rect 242750 1458 242756 1460
rect 226517 1456 238770 1458
rect 226517 1400 226522 1456
rect 226578 1400 238770 1456
rect 226517 1398 238770 1400
rect 242710 1398 242756 1458
rect 242820 1456 242867 1460
rect 245694 1458 245700 1460
rect 242862 1400 242867 1456
rect 226517 1395 226583 1398
rect 242750 1396 242756 1398
rect 242820 1396 242867 1400
rect 245654 1398 245700 1458
rect 245764 1456 245811 1460
rect 245806 1400 245811 1456
rect 245694 1396 245700 1398
rect 245764 1396 245811 1400
rect 248638 1396 248644 1460
rect 248708 1458 248714 1460
rect 249793 1458 249859 1461
rect 248708 1456 249859 1458
rect 248708 1400 249798 1456
rect 249854 1400 249859 1456
rect 248708 1398 249859 1400
rect 248708 1396 248714 1398
rect 242801 1395 242867 1396
rect 245745 1395 245811 1396
rect 249793 1395 249859 1398
rect 252318 1396 252324 1460
rect 252388 1458 252394 1460
rect 252645 1458 252711 1461
rect 252388 1456 252711 1458
rect 252388 1400 252650 1456
rect 252706 1400 252711 1456
rect 252388 1398 252711 1400
rect 252388 1396 252394 1398
rect 252645 1395 252711 1398
rect 255221 1458 255287 1461
rect 257521 1460 257587 1461
rect 257470 1458 257476 1460
rect 255221 1456 257354 1458
rect 255221 1400 255226 1456
rect 255282 1400 257354 1456
rect 255221 1398 257354 1400
rect 257430 1398 257476 1458
rect 257540 1456 257587 1460
rect 258398 1458 258458 1534
rect 269849 1531 269915 1534
rect 271965 1531 272031 1534
rect 272149 1594 272215 1597
rect 272149 1592 272504 1594
rect 272149 1536 272154 1592
rect 272210 1536 272504 1592
rect 272149 1534 272504 1536
rect 272149 1531 272215 1534
rect 257582 1400 257587 1456
rect 255221 1395 255287 1398
rect 88014 1262 88626 1322
rect 88926 1260 88932 1324
rect 88996 1322 89002 1324
rect 89529 1322 89595 1325
rect 88996 1320 89595 1322
rect 88996 1264 89534 1320
rect 89590 1264 89595 1320
rect 88996 1262 89595 1264
rect 88996 1260 89002 1262
rect 25773 1259 25839 1260
rect 26509 1259 26575 1260
rect 76465 1259 76531 1260
rect 78673 1259 78739 1260
rect 81617 1259 81683 1260
rect 83825 1259 83891 1260
rect 89529 1259 89595 1262
rect 89846 1260 89852 1324
rect 89916 1322 89922 1324
rect 90173 1322 90239 1325
rect 89916 1320 90239 1322
rect 89916 1264 90178 1320
rect 90234 1264 90239 1320
rect 89916 1262 90239 1264
rect 89916 1260 89922 1262
rect 90173 1259 90239 1262
rect 90398 1260 90404 1324
rect 90468 1322 90474 1324
rect 90817 1322 90883 1325
rect 90468 1320 90883 1322
rect 90468 1264 90822 1320
rect 90878 1264 90883 1320
rect 90468 1262 90883 1264
rect 90468 1260 90474 1262
rect 90817 1259 90883 1262
rect 91870 1260 91876 1324
rect 91940 1322 91946 1324
rect 92013 1322 92079 1325
rect 91940 1320 92079 1322
rect 91940 1264 92018 1320
rect 92074 1264 92079 1320
rect 91940 1262 92079 1264
rect 91940 1260 91946 1262
rect 92013 1259 92079 1262
rect 92749 1322 92815 1325
rect 93342 1322 93348 1324
rect 92749 1320 93348 1322
rect 92749 1264 92754 1320
rect 92810 1264 93348 1320
rect 92749 1262 93348 1264
rect 92749 1259 92815 1262
rect 93342 1260 93348 1262
rect 93412 1260 93418 1324
rect 99189 1322 99255 1325
rect 104065 1322 104131 1325
rect 99189 1320 104131 1322
rect 99189 1264 99194 1320
rect 99250 1264 104070 1320
rect 104126 1264 104131 1320
rect 99189 1262 104131 1264
rect 99189 1259 99255 1262
rect 104065 1259 104131 1262
rect 144545 1322 144611 1325
rect 152457 1322 152523 1325
rect 144545 1320 152523 1322
rect 144545 1264 144550 1320
rect 144606 1264 152462 1320
rect 152518 1264 152523 1320
rect 144545 1262 152523 1264
rect 144545 1259 144611 1262
rect 152457 1259 152523 1262
rect 152774 1260 152780 1324
rect 152844 1322 152850 1324
rect 154481 1322 154547 1325
rect 152844 1320 154547 1322
rect 152844 1264 154486 1320
rect 154542 1264 154547 1320
rect 152844 1262 154547 1264
rect 152844 1260 152850 1262
rect 154481 1259 154547 1262
rect 157926 1260 157932 1324
rect 157996 1322 158002 1324
rect 158621 1322 158687 1325
rect 157996 1320 158687 1322
rect 157996 1264 158626 1320
rect 158682 1264 158687 1320
rect 157996 1262 158687 1264
rect 157996 1260 158002 1262
rect 158621 1259 158687 1262
rect 160369 1322 160435 1325
rect 166993 1322 167059 1325
rect 160369 1320 167059 1322
rect 160369 1264 160374 1320
rect 160430 1264 166998 1320
rect 167054 1264 167059 1320
rect 160369 1262 167059 1264
rect 160369 1259 160435 1262
rect 166993 1259 167059 1262
rect 218053 1322 218119 1325
rect 220813 1322 220879 1325
rect 218053 1320 220879 1322
rect 218053 1264 218058 1320
rect 218114 1264 220818 1320
rect 220874 1264 220879 1320
rect 218053 1262 220879 1264
rect 218053 1259 218119 1262
rect 220813 1259 220879 1262
rect 222193 1322 222259 1325
rect 226241 1322 226307 1325
rect 222193 1320 226307 1322
rect 222193 1264 222198 1320
rect 222254 1264 226246 1320
rect 226302 1264 226307 1320
rect 222193 1262 226307 1264
rect 222193 1259 222259 1262
rect 226241 1259 226307 1262
rect 228633 1322 228699 1325
rect 243537 1322 243603 1325
rect 257294 1322 257354 1398
rect 257470 1396 257476 1398
rect 257540 1396 257587 1400
rect 257521 1395 257587 1396
rect 257662 1398 258458 1458
rect 258717 1458 258783 1461
rect 258717 1456 272504 1458
rect 258717 1400 258722 1456
rect 258778 1400 272504 1456
rect 258717 1398 272504 1400
rect 257662 1322 257722 1398
rect 258717 1395 258783 1398
rect 228633 1320 238770 1322
rect 228633 1264 228638 1320
rect 228694 1264 238770 1320
rect 228633 1262 238770 1264
rect 228633 1259 228699 1262
rect 29494 1124 29500 1188
rect 29564 1186 29570 1188
rect 29913 1186 29979 1189
rect 29564 1184 29979 1186
rect 29564 1128 29918 1184
rect 29974 1128 29979 1184
rect 29564 1126 29979 1128
rect 29564 1124 29570 1126
rect 29913 1123 29979 1126
rect 88517 1186 88583 1189
rect 112345 1186 112411 1189
rect 88517 1184 112411 1186
rect 88517 1128 88522 1184
rect 88578 1128 112350 1184
rect 112406 1128 112411 1184
rect 88517 1126 112411 1128
rect 88517 1123 88583 1126
rect 112345 1123 112411 1126
rect 149513 1186 149579 1189
rect 155769 1186 155835 1189
rect 149513 1184 155835 1186
rect 149513 1128 149518 1184
rect 149574 1128 155774 1184
rect 155830 1128 155835 1184
rect 149513 1126 155835 1128
rect 149513 1123 149579 1126
rect 155769 1123 155835 1126
rect 158662 1124 158668 1188
rect 158732 1186 158738 1188
rect 159357 1186 159423 1189
rect 158732 1184 159423 1186
rect 158732 1128 159362 1184
rect 159418 1128 159423 1184
rect 158732 1126 159423 1128
rect 158732 1124 158738 1126
rect 159357 1123 159423 1126
rect 160134 1124 160140 1188
rect 160204 1186 160210 1188
rect 160829 1186 160895 1189
rect 161657 1188 161723 1189
rect 163865 1188 163931 1189
rect 161606 1186 161612 1188
rect 160204 1184 160895 1186
rect 160204 1128 160834 1184
rect 160890 1128 160895 1184
rect 160204 1126 160895 1128
rect 161566 1126 161612 1186
rect 161676 1184 161723 1188
rect 163814 1186 163820 1188
rect 161718 1128 161723 1184
rect 160204 1124 160210 1126
rect 160829 1123 160895 1126
rect 161606 1124 161612 1126
rect 161676 1124 161723 1128
rect 163774 1126 163820 1186
rect 163884 1184 163931 1188
rect 163926 1128 163931 1184
rect 163814 1124 163820 1126
rect 163884 1124 163931 1128
rect 161657 1123 161723 1124
rect 163865 1123 163931 1124
rect 165245 1188 165311 1189
rect 165981 1188 166047 1189
rect 166809 1188 166875 1189
rect 165245 1184 165292 1188
rect 165356 1186 165362 1188
rect 165245 1128 165250 1184
rect 165245 1124 165292 1128
rect 165356 1126 165402 1186
rect 165981 1184 166028 1188
rect 166092 1186 166098 1188
rect 166758 1186 166764 1188
rect 165981 1128 165986 1184
rect 165356 1124 165362 1126
rect 165981 1124 166028 1128
rect 166092 1126 166138 1186
rect 166718 1126 166764 1186
rect 166828 1184 166875 1188
rect 166870 1128 166875 1184
rect 166092 1124 166098 1126
rect 166758 1124 166764 1126
rect 166828 1124 166875 1128
rect 165245 1123 165311 1124
rect 165981 1123 166047 1124
rect 166809 1123 166875 1124
rect 211797 1186 211863 1189
rect 223481 1186 223547 1189
rect 211797 1184 223547 1186
rect 211797 1128 211802 1184
rect 211858 1128 223486 1184
rect 223542 1128 223547 1184
rect 211797 1126 223547 1128
rect 211797 1123 211863 1126
rect 223481 1123 223547 1126
rect 223982 1124 223988 1188
rect 224052 1186 224058 1188
rect 224217 1186 224283 1189
rect 224052 1184 224283 1186
rect 224052 1128 224222 1184
rect 224278 1128 224283 1184
rect 224052 1126 224283 1128
rect 224052 1124 224058 1126
rect 224217 1123 224283 1126
rect 225454 1124 225460 1188
rect 225524 1186 225530 1188
rect 225689 1186 225755 1189
rect 225524 1184 225755 1186
rect 225524 1128 225694 1184
rect 225750 1128 225755 1184
rect 225524 1126 225755 1128
rect 225524 1124 225530 1126
rect 225689 1123 225755 1126
rect 227662 1124 227668 1188
rect 227732 1186 227738 1188
rect 227989 1186 228055 1189
rect 227732 1184 228055 1186
rect 227732 1128 227994 1184
rect 228050 1128 228055 1184
rect 227732 1126 228055 1128
rect 227732 1124 227738 1126
rect 227989 1123 228055 1126
rect 229870 1124 229876 1188
rect 229940 1186 229946 1188
rect 230013 1186 230079 1189
rect 229940 1184 230079 1186
rect 229940 1128 230018 1184
rect 230074 1128 230079 1184
rect 229940 1126 230079 1128
rect 229940 1124 229946 1126
rect 230013 1123 230079 1126
rect 230606 1124 230612 1188
rect 230676 1186 230682 1188
rect 231577 1186 231643 1189
rect 230676 1184 231643 1186
rect 230676 1128 231582 1184
rect 231638 1128 231643 1184
rect 230676 1126 231643 1128
rect 230676 1124 230682 1126
rect 231577 1123 231643 1126
rect 232078 1124 232084 1188
rect 232148 1186 232154 1188
rect 232405 1186 232471 1189
rect 232148 1184 232471 1186
rect 232148 1128 232410 1184
rect 232466 1128 232471 1184
rect 232148 1126 232471 1128
rect 232148 1124 232154 1126
rect 232405 1123 232471 1126
rect 232814 1124 232820 1188
rect 232884 1186 232890 1188
rect 233141 1186 233207 1189
rect 232884 1184 233207 1186
rect 232884 1128 233146 1184
rect 233202 1128 233207 1184
rect 232884 1126 233207 1128
rect 232884 1124 232890 1126
rect 233141 1123 233207 1126
rect 235022 1124 235028 1188
rect 235092 1186 235098 1188
rect 235165 1186 235231 1189
rect 235092 1184 235231 1186
rect 235092 1128 235170 1184
rect 235226 1128 235231 1184
rect 235092 1126 235231 1128
rect 235092 1124 235098 1126
rect 235165 1123 235231 1126
rect 236494 1124 236500 1188
rect 236564 1186 236570 1188
rect 236821 1186 236887 1189
rect 236564 1184 236887 1186
rect 236564 1128 236826 1184
rect 236882 1128 236887 1184
rect 236564 1126 236887 1128
rect 238710 1186 238770 1262
rect 243537 1320 255882 1322
rect 243537 1264 243542 1320
rect 243598 1264 255882 1320
rect 243537 1262 255882 1264
rect 257294 1262 257722 1322
rect 268009 1322 268075 1325
rect 271965 1322 272031 1325
rect 268009 1320 271890 1322
rect 268009 1264 268014 1320
rect 268070 1264 271890 1320
rect 268009 1262 271890 1264
rect 243537 1259 243603 1262
rect 255681 1186 255747 1189
rect 238710 1184 255747 1186
rect 238710 1128 255686 1184
rect 255742 1128 255747 1184
rect 238710 1126 255747 1128
rect 255822 1186 255882 1262
rect 268009 1259 268075 1262
rect 257797 1186 257863 1189
rect 255822 1184 257863 1186
rect 255822 1128 257802 1184
rect 257858 1128 257863 1184
rect 255822 1126 257863 1128
rect 271830 1186 271890 1262
rect 271965 1320 272504 1322
rect 271965 1264 271970 1320
rect 272026 1264 272504 1320
rect 271965 1262 272504 1264
rect 271965 1259 272031 1262
rect 271830 1126 272504 1186
rect 236564 1124 236570 1126
rect 236821 1123 236887 1126
rect 255681 1123 255747 1126
rect 257797 1123 257863 1126
rect 68542 1120 68858 1121
rect 68542 1056 68548 1120
rect 68612 1056 68628 1120
rect 68692 1056 68708 1120
rect 68772 1056 68788 1120
rect 68852 1056 68858 1120
rect 68542 1055 68858 1056
rect 136139 1120 136455 1121
rect 136139 1056 136145 1120
rect 136209 1056 136225 1120
rect 136289 1056 136305 1120
rect 136369 1056 136385 1120
rect 136449 1056 136455 1120
rect 136139 1055 136455 1056
rect 203736 1120 204052 1121
rect 203736 1056 203742 1120
rect 203806 1056 203822 1120
rect 203886 1056 203902 1120
rect 203966 1056 203982 1120
rect 204046 1056 204052 1120
rect 203736 1055 204052 1056
rect 271333 1120 271649 1121
rect 271333 1056 271339 1120
rect 271403 1056 271419 1120
rect 271483 1056 271499 1120
rect 271563 1056 271579 1120
rect 271643 1056 271649 1120
rect 271333 1055 271649 1056
rect 1526 988 1532 1052
rect 1596 1050 1602 1052
rect 1669 1050 1735 1053
rect 3785 1052 3851 1053
rect 3734 1050 3740 1052
rect 1596 1048 1735 1050
rect 1596 992 1674 1048
rect 1730 992 1735 1048
rect 1596 990 1735 992
rect 3694 990 3740 1050
rect 3804 1048 3851 1052
rect 3846 992 3851 1048
rect 1596 988 1602 990
rect 1669 987 1735 990
rect 3734 988 3740 990
rect 3804 988 3851 992
rect 3785 987 3851 988
rect 5165 1052 5231 1053
rect 5165 1048 5212 1052
rect 5276 1050 5282 1052
rect 7097 1050 7163 1053
rect 9673 1052 9739 1053
rect 7414 1050 7420 1052
rect 5165 992 5170 1048
rect 5165 988 5212 992
rect 5276 990 5322 1050
rect 7097 1048 7420 1050
rect 7097 992 7102 1048
rect 7158 992 7420 1048
rect 7097 990 7420 992
rect 5276 988 5282 990
rect 5165 987 5231 988
rect 7097 987 7163 990
rect 7414 988 7420 990
rect 7484 988 7490 1052
rect 9622 1050 9628 1052
rect 9582 990 9628 1050
rect 9692 1048 9739 1052
rect 9734 992 9739 1048
rect 9622 988 9628 990
rect 9692 988 9739 992
rect 11830 988 11836 1052
rect 11900 1050 11906 1052
rect 11973 1050 12039 1053
rect 11900 1048 12039 1050
rect 11900 992 11978 1048
rect 12034 992 12039 1048
rect 11900 990 12039 992
rect 11900 988 11906 990
rect 9673 987 9739 988
rect 11973 987 12039 990
rect 12566 988 12572 1052
rect 12636 1050 12642 1052
rect 12709 1050 12775 1053
rect 14089 1052 14155 1053
rect 14038 1050 14044 1052
rect 12636 1048 12775 1050
rect 12636 992 12714 1048
rect 12770 992 12775 1048
rect 12636 990 12775 992
rect 13998 990 14044 1050
rect 14108 1048 14155 1052
rect 14150 992 14155 1048
rect 12636 988 12642 990
rect 12709 987 12775 990
rect 14038 988 14044 990
rect 14108 988 14155 992
rect 14089 987 14155 988
rect 15469 1052 15535 1053
rect 15469 1048 15516 1052
rect 15580 1050 15586 1052
rect 15469 992 15474 1048
rect 15469 988 15516 992
rect 15580 990 15626 1050
rect 15580 988 15586 990
rect 17718 988 17724 1052
rect 17788 1050 17794 1052
rect 17861 1050 17927 1053
rect 17788 1048 17927 1050
rect 17788 992 17866 1048
rect 17922 992 17927 1048
rect 17788 990 17927 992
rect 17788 988 17794 990
rect 15469 987 15535 988
rect 17861 987 17927 990
rect 71262 988 71268 1052
rect 71332 1050 71338 1052
rect 71497 1050 71563 1053
rect 71332 1048 71563 1050
rect 71332 992 71502 1048
rect 71558 992 71563 1048
rect 71332 990 71563 992
rect 71332 988 71338 990
rect 71497 987 71563 990
rect 71998 988 72004 1052
rect 72068 1050 72074 1052
rect 72233 1050 72299 1053
rect 72068 1048 72299 1050
rect 72068 992 72238 1048
rect 72294 992 72299 1048
rect 72068 990 72299 992
rect 72068 988 72074 990
rect 72233 987 72299 990
rect 73470 988 73476 1052
rect 73540 1050 73546 1052
rect 73705 1050 73771 1053
rect 75729 1052 75795 1053
rect 77201 1052 77267 1053
rect 79409 1052 79475 1053
rect 80881 1052 80947 1053
rect 82353 1052 82419 1053
rect 84561 1052 84627 1053
rect 86033 1052 86099 1053
rect 75678 1050 75684 1052
rect 73540 1048 73771 1050
rect 73540 992 73710 1048
rect 73766 992 73771 1048
rect 73540 990 73771 992
rect 75638 990 75684 1050
rect 75748 1048 75795 1052
rect 77150 1050 77156 1052
rect 75790 992 75795 1048
rect 73540 988 73546 990
rect 73705 987 73771 990
rect 75678 988 75684 990
rect 75748 988 75795 992
rect 77110 990 77156 1050
rect 77220 1048 77267 1052
rect 79358 1050 79364 1052
rect 77262 992 77267 1048
rect 77150 988 77156 990
rect 77220 988 77267 992
rect 79318 990 79364 1050
rect 79428 1048 79475 1052
rect 80830 1050 80836 1052
rect 79470 992 79475 1048
rect 79358 988 79364 990
rect 79428 988 79475 992
rect 80790 990 80836 1050
rect 80900 1048 80947 1052
rect 82302 1050 82308 1052
rect 80942 992 80947 1048
rect 80830 988 80836 990
rect 80900 988 80947 992
rect 82262 990 82308 1050
rect 82372 1048 82419 1052
rect 84510 1050 84516 1052
rect 82414 992 82419 1048
rect 82302 988 82308 990
rect 82372 988 82419 992
rect 84470 990 84516 1050
rect 84580 1048 84627 1052
rect 85982 1050 85988 1052
rect 84622 992 84627 1048
rect 84510 988 84516 990
rect 84580 988 84627 992
rect 85942 990 85988 1050
rect 86052 1048 86099 1052
rect 86094 992 86099 1048
rect 85982 988 85988 990
rect 86052 988 86099 992
rect 75729 987 75795 988
rect 77201 987 77267 988
rect 79409 987 79475 988
rect 80881 987 80947 988
rect 82353 987 82419 988
rect 84561 987 84627 988
rect 86033 987 86099 988
rect 93025 1050 93091 1053
rect 94589 1050 94655 1053
rect 115105 1050 115171 1053
rect 93025 1048 94655 1050
rect 93025 992 93030 1048
rect 93086 992 94594 1048
rect 94650 992 94655 1048
rect 93025 990 94655 992
rect 93025 987 93091 990
rect 94589 987 94655 990
rect 94822 1048 115171 1050
rect 94822 992 115110 1048
rect 115166 992 115171 1048
rect 94822 990 115171 992
rect 69105 916 69171 917
rect 69054 914 69060 916
rect 69014 854 69060 914
rect 69124 912 69171 916
rect 69166 856 69171 912
rect 69054 852 69060 854
rect 69124 852 69171 856
rect 69105 851 69171 852
rect 69565 914 69631 917
rect 69790 914 69796 916
rect 69565 912 69796 914
rect 69565 856 69570 912
rect 69626 856 69796 912
rect 69565 854 69796 856
rect 69565 851 69631 854
rect 69790 852 69796 854
rect 69860 852 69866 916
rect 70526 852 70532 916
rect 70596 914 70602 916
rect 70945 914 71011 917
rect 70596 912 71011 914
rect 70596 856 70950 912
rect 71006 856 71011 912
rect 70596 854 71011 856
rect 70596 852 70602 854
rect 70945 851 71011 854
rect 72734 852 72740 916
rect 72804 914 72810 916
rect 72969 914 73035 917
rect 74257 916 74323 917
rect 74206 914 74212 916
rect 72804 912 73035 914
rect 72804 856 72974 912
rect 73030 856 73035 912
rect 72804 854 73035 856
rect 74166 854 74212 914
rect 74276 912 74323 916
rect 74318 856 74323 912
rect 72804 852 72810 854
rect 72969 851 73035 854
rect 74206 852 74212 854
rect 74276 852 74323 856
rect 74257 851 74323 852
rect 74717 914 74783 917
rect 74942 914 74948 916
rect 74717 912 74948 914
rect 74717 856 74722 912
rect 74778 856 74948 912
rect 74717 854 74948 856
rect 74717 851 74783 854
rect 74942 852 74948 854
rect 75012 852 75018 916
rect 77293 914 77359 917
rect 77886 914 77892 916
rect 77293 912 77892 914
rect 77293 856 77298 912
rect 77354 856 77892 912
rect 77293 854 77892 856
rect 77293 851 77359 854
rect 77886 852 77892 854
rect 77956 852 77962 916
rect 79961 914 80027 917
rect 80094 914 80100 916
rect 79961 912 80100 914
rect 79961 856 79966 912
rect 80022 856 80100 912
rect 79961 854 80100 856
rect 79961 851 80027 854
rect 80094 852 80100 854
rect 80164 852 80170 916
rect 82629 914 82695 917
rect 86769 916 86835 917
rect 83038 914 83044 916
rect 82629 912 83044 914
rect 82629 856 82634 912
rect 82690 856 83044 912
rect 82629 854 83044 856
rect 82629 851 82695 854
rect 83038 852 83044 854
rect 83108 852 83114 916
rect 86718 914 86724 916
rect 86678 854 86724 914
rect 86788 912 86835 916
rect 86830 856 86835 912
rect 86718 852 86724 854
rect 86788 852 86835 856
rect 86769 851 86835 852
rect 92381 914 92447 917
rect 94822 914 94882 990
rect 115105 987 115171 990
rect 139526 988 139532 1052
rect 139596 1050 139602 1052
rect 139761 1050 139827 1053
rect 139596 1048 139827 1050
rect 139596 992 139766 1048
rect 139822 992 139827 1048
rect 139596 990 139827 992
rect 139596 988 139602 990
rect 139761 987 139827 990
rect 148317 1050 148383 1053
rect 151353 1050 151419 1053
rect 152365 1050 152431 1053
rect 148317 1048 152431 1050
rect 148317 992 148322 1048
rect 148378 992 151358 1048
rect 151414 992 152370 1048
rect 152426 992 152431 1048
rect 148317 990 152431 992
rect 148317 987 148383 990
rect 151353 987 151419 990
rect 152365 987 152431 990
rect 158437 1050 158503 1053
rect 168373 1050 168439 1053
rect 158437 1048 168439 1050
rect 158437 992 158442 1048
rect 158498 992 168378 1048
rect 168434 992 168439 1048
rect 158437 990 168439 992
rect 158437 987 158503 990
rect 168373 987 168439 990
rect 170305 1050 170371 1053
rect 180517 1050 180583 1053
rect 209773 1050 209839 1053
rect 170305 1048 180583 1050
rect 170305 992 170310 1048
rect 170366 992 180522 1048
rect 180578 992 180583 1048
rect 170305 990 180583 992
rect 170305 987 170371 990
rect 180517 987 180583 990
rect 205406 1048 209839 1050
rect 205406 992 209778 1048
rect 209834 992 209839 1048
rect 205406 990 209839 992
rect 92381 912 94882 914
rect 92381 856 92386 912
rect 92442 856 94882 912
rect 92381 854 94882 856
rect 92381 851 92447 854
rect 99230 852 99236 916
rect 99300 914 99306 916
rect 100753 914 100819 917
rect 99300 912 100819 914
rect 99300 856 100758 912
rect 100814 856 100819 912
rect 99300 854 100819 856
rect 99300 852 99306 854
rect 100753 851 100819 854
rect 104157 914 104223 917
rect 114921 914 114987 917
rect 143625 914 143691 917
rect 104157 912 114987 914
rect 104157 856 104162 912
rect 104218 856 114926 912
rect 114982 856 114987 912
rect 104157 854 114987 856
rect 104157 851 104223 854
rect 114921 851 114987 854
rect 122790 912 143691 914
rect 122790 856 143630 912
rect 143686 856 143691 912
rect 122790 854 143691 856
rect 2957 780 3023 781
rect 2957 776 3004 780
rect 3068 778 3074 780
rect 5349 778 5415 781
rect 10317 780 10383 781
rect 5942 778 5948 780
rect 2957 720 2962 776
rect 2957 716 3004 720
rect 3068 718 3114 778
rect 5349 776 5948 778
rect 5349 720 5354 776
rect 5410 720 5948 776
rect 5349 718 5948 720
rect 3068 716 3074 718
rect 2957 715 3023 716
rect 5349 715 5415 718
rect 5942 716 5948 718
rect 6012 716 6018 780
rect 10317 776 10364 780
rect 10428 778 10434 780
rect 10317 720 10322 776
rect 10317 716 10364 720
rect 10428 718 10474 778
rect 10428 716 10434 718
rect 11094 716 11100 780
rect 11164 778 11170 780
rect 11697 778 11763 781
rect 11164 776 11763 778
rect 11164 720 11702 776
rect 11758 720 11763 776
rect 11164 718 11763 720
rect 11164 716 11170 718
rect 10317 715 10383 716
rect 11697 715 11763 718
rect 15653 778 15719 781
rect 17033 780 17099 781
rect 16246 778 16252 780
rect 15653 776 16252 778
rect 15653 720 15658 776
rect 15714 720 16252 776
rect 15653 718 16252 720
rect 15653 715 15719 718
rect 16246 716 16252 718
rect 16316 716 16322 780
rect 16982 778 16988 780
rect 16942 718 16988 778
rect 17052 776 17099 780
rect 17094 720 17099 776
rect 16982 716 16988 718
rect 17052 716 17099 720
rect 17033 715 17099 716
rect 45737 778 45803 781
rect 108481 778 108547 781
rect 45737 776 108547 778
rect 45737 720 45742 776
rect 45798 720 108486 776
rect 108542 720 108547 776
rect 45737 718 108547 720
rect 45737 715 45803 718
rect 108481 715 108547 718
rect 1945 642 2011 645
rect 2262 642 2268 644
rect 1945 640 2268 642
rect 1945 584 1950 640
rect 2006 584 2268 640
rect 1945 582 2268 584
rect 1945 579 2011 582
rect 2262 580 2268 582
rect 2332 580 2338 644
rect 13302 580 13308 644
rect 13372 642 13378 644
rect 13445 642 13511 645
rect 21449 644 21515 645
rect 21398 642 21404 644
rect 13372 640 13511 642
rect 13372 584 13450 640
rect 13506 584 13511 640
rect 13372 582 13511 584
rect 21358 582 21404 642
rect 21468 640 21515 644
rect 21510 584 21515 640
rect 13372 580 13378 582
rect 13445 579 13511 582
rect 21398 580 21404 582
rect 21468 580 21515 584
rect 28022 580 28028 644
rect 28092 642 28098 644
rect 28165 642 28231 645
rect 30281 644 30347 645
rect 30230 642 30236 644
rect 28092 640 28231 642
rect 28092 584 28170 640
rect 28226 584 28231 640
rect 28092 582 28231 584
rect 30190 582 30236 642
rect 30300 640 30347 644
rect 30342 584 30347 640
rect 28092 580 28098 582
rect 21449 579 21515 580
rect 28165 579 28231 582
rect 30230 580 30236 582
rect 30300 580 30347 584
rect 30966 580 30972 644
rect 31036 642 31042 644
rect 31201 642 31267 645
rect 31036 640 31267 642
rect 31036 584 31206 640
rect 31262 584 31267 640
rect 31036 582 31267 584
rect 31036 580 31042 582
rect 30281 579 30347 580
rect 31201 579 31267 582
rect 31702 580 31708 644
rect 31772 642 31778 644
rect 32489 642 32555 645
rect 31772 640 32555 642
rect 31772 584 32494 640
rect 32550 584 32555 640
rect 31772 582 32555 584
rect 31772 580 31778 582
rect 32489 579 32555 582
rect 34922 580 34928 644
rect 34992 642 34998 644
rect 35157 642 35223 645
rect 34992 640 35223 642
rect 34992 584 35162 640
rect 35218 584 35223 640
rect 34992 582 35223 584
rect 34992 580 34998 582
rect 35157 579 35223 582
rect 35617 644 35683 645
rect 35617 640 35664 644
rect 35728 642 35734 644
rect 36261 642 36327 645
rect 36394 642 36400 644
rect 35617 584 35622 640
rect 35617 580 35664 584
rect 35728 582 35774 642
rect 36261 640 36400 642
rect 36261 584 36266 640
rect 36322 584 36400 640
rect 36261 582 36400 584
rect 35728 580 35734 582
rect 35617 579 35683 580
rect 36261 579 36327 582
rect 36394 580 36400 582
rect 36464 580 36470 644
rect 36905 642 36971 645
rect 37130 642 37136 644
rect 36905 640 37136 642
rect 36905 584 36910 640
rect 36966 584 37136 640
rect 36905 582 37136 584
rect 36905 579 36971 582
rect 37130 580 37136 582
rect 37200 580 37206 644
rect 37866 580 37872 644
rect 37936 642 37942 644
rect 38101 642 38167 645
rect 37936 640 38167 642
rect 37936 584 38106 640
rect 38162 584 38167 640
rect 37936 582 38167 584
rect 37936 580 37942 582
rect 38101 579 38167 582
rect 38561 644 38627 645
rect 38561 640 38608 644
rect 38672 642 38678 644
rect 39941 642 40007 645
rect 40769 644 40835 645
rect 40074 642 40080 644
rect 38561 584 38566 640
rect 38561 580 38608 584
rect 38672 582 38718 642
rect 39941 640 40080 642
rect 39941 584 39946 640
rect 40002 584 40080 640
rect 39941 582 40080 584
rect 38672 580 38678 582
rect 38561 579 38627 580
rect 39941 579 40007 582
rect 40074 580 40080 582
rect 40144 580 40150 644
rect 40769 640 40816 644
rect 40880 642 40886 644
rect 41413 642 41479 645
rect 41546 642 41552 644
rect 40769 584 40774 640
rect 40769 580 40816 584
rect 40880 582 40926 642
rect 41413 640 41552 642
rect 41413 584 41418 640
rect 41474 584 41552 640
rect 41413 582 41552 584
rect 40880 580 40886 582
rect 40769 579 40835 580
rect 41413 579 41479 582
rect 41546 580 41552 582
rect 41616 580 41622 644
rect 42057 642 42123 645
rect 42282 642 42288 644
rect 42057 640 42288 642
rect 42057 584 42062 640
rect 42118 584 42288 640
rect 42057 582 42288 584
rect 42057 579 42123 582
rect 42282 580 42288 582
rect 42352 580 42358 644
rect 43018 580 43024 644
rect 43088 642 43094 644
rect 43253 642 43319 645
rect 43088 640 43319 642
rect 43088 584 43258 640
rect 43314 584 43319 640
rect 43088 582 43319 584
rect 43088 580 43094 582
rect 43253 579 43319 582
rect 43754 580 43760 644
rect 43824 642 43830 644
rect 43989 642 44055 645
rect 43824 640 44055 642
rect 43824 584 43994 640
rect 44050 584 44055 640
rect 43824 582 44055 584
rect 43824 580 43830 582
rect 43989 579 44055 582
rect 44490 580 44496 644
rect 44560 642 44566 644
rect 44633 642 44699 645
rect 44560 640 44699 642
rect 44560 584 44638 640
rect 44694 584 44699 640
rect 44560 582 44699 584
rect 44560 580 44566 582
rect 44633 579 44699 582
rect 45226 580 45232 644
rect 45296 642 45302 644
rect 45461 642 45527 645
rect 45296 640 45527 642
rect 45296 584 45466 640
rect 45522 584 45527 640
rect 45296 582 45527 584
rect 45296 580 45302 582
rect 45461 579 45527 582
rect 45921 644 45987 645
rect 45921 640 45968 644
rect 46032 642 46038 644
rect 46565 642 46631 645
rect 46698 642 46704 644
rect 45921 584 45926 640
rect 45921 580 45968 584
rect 46032 582 46078 642
rect 46565 640 46704 642
rect 46565 584 46570 640
rect 46626 584 46704 640
rect 46565 582 46704 584
rect 46032 580 46038 582
rect 45921 579 45987 580
rect 46565 579 46631 582
rect 46698 580 46704 582
rect 46768 580 46774 644
rect 47209 642 47275 645
rect 48221 644 48287 645
rect 47434 642 47440 644
rect 47209 640 47440 642
rect 47209 584 47214 640
rect 47270 584 47440 640
rect 47209 582 47440 584
rect 47209 579 47275 582
rect 47434 580 47440 582
rect 47504 580 47510 644
rect 48170 642 48176 644
rect 48130 582 48176 642
rect 48240 640 48287 644
rect 48282 584 48287 640
rect 48170 580 48176 582
rect 48240 580 48287 584
rect 48906 580 48912 644
rect 48976 642 48982 644
rect 49141 642 49207 645
rect 48976 640 49207 642
rect 48976 584 49146 640
rect 49202 584 49207 640
rect 48976 582 49207 584
rect 48976 580 48982 582
rect 48221 579 48287 580
rect 49141 579 49207 582
rect 49642 580 49648 644
rect 49712 642 49718 644
rect 49785 642 49851 645
rect 49712 640 49851 642
rect 49712 584 49790 640
rect 49846 584 49851 640
rect 49712 582 49851 584
rect 49712 580 49718 582
rect 49785 579 49851 582
rect 50378 580 50384 644
rect 50448 642 50454 644
rect 50613 642 50679 645
rect 50448 640 50679 642
rect 50448 584 50618 640
rect 50674 584 50679 640
rect 50448 582 50679 584
rect 50448 580 50454 582
rect 50613 579 50679 582
rect 51114 580 51120 644
rect 51184 642 51190 644
rect 51349 642 51415 645
rect 51184 640 51415 642
rect 51184 584 51354 640
rect 51410 584 51415 640
rect 51184 582 51415 584
rect 51184 580 51190 582
rect 51349 579 51415 582
rect 51850 580 51856 644
rect 51920 642 51926 644
rect 52085 642 52151 645
rect 51920 640 52151 642
rect 51920 584 52090 640
rect 52146 584 52151 640
rect 51920 582 52151 584
rect 51920 580 51926 582
rect 52085 579 52151 582
rect 52913 642 52979 645
rect 53322 642 53328 644
rect 52913 640 53328 642
rect 52913 584 52918 640
rect 52974 584 53328 640
rect 52913 582 53328 584
rect 52913 579 52979 582
rect 53322 580 53328 582
rect 53392 580 53398 644
rect 54058 580 54064 644
rect 54128 642 54134 644
rect 54477 642 54543 645
rect 92197 642 92263 645
rect 54128 640 54543 642
rect 54128 584 54482 640
rect 54538 584 54543 640
rect 54128 582 54543 584
rect 54128 580 54134 582
rect 54477 579 54543 582
rect 55170 640 92263 642
rect 55170 584 92202 640
rect 92258 584 92263 640
rect 55170 582 92263 584
rect 7741 506 7807 509
rect 8150 506 8156 508
rect 7741 504 8156 506
rect 7741 448 7746 504
rect 7802 448 8156 504
rect 7741 446 8156 448
rect 7741 443 7807 446
rect 8150 444 8156 446
rect 8220 444 8226 508
rect 39849 506 39915 509
rect 55170 506 55230 582
rect 92197 579 92263 582
rect 92473 642 92539 645
rect 94773 644 94839 645
rect 92606 642 92612 644
rect 92473 640 92612 642
rect 92473 584 92478 640
rect 92534 584 92612 640
rect 92473 582 92612 584
rect 92473 579 92539 582
rect 92606 580 92612 582
rect 92676 580 92682 644
rect 94773 640 94820 644
rect 94884 642 94890 644
rect 99281 642 99347 645
rect 99966 642 99972 644
rect 94773 584 94778 640
rect 94773 580 94820 584
rect 94884 582 94930 642
rect 99281 640 99972 642
rect 99281 584 99286 640
rect 99342 584 99972 640
rect 99281 582 99972 584
rect 94884 580 94890 582
rect 94773 579 94839 580
rect 99281 579 99347 582
rect 99966 580 99972 582
rect 100036 580 100042 644
rect 104065 642 104131 645
rect 122790 642 122850 854
rect 143625 851 143691 854
rect 144729 914 144795 917
rect 205406 914 205466 990
rect 209730 987 209839 990
rect 211889 1050 211955 1053
rect 243629 1050 243695 1053
rect 211889 1048 243695 1050
rect 211889 992 211894 1048
rect 211950 992 243634 1048
rect 243690 992 243695 1048
rect 211889 990 243695 992
rect 211889 987 211955 990
rect 243629 987 243695 990
rect 246941 1050 247007 1053
rect 266302 1050 266308 1052
rect 246941 1048 266308 1050
rect 246941 992 246946 1048
rect 247002 992 266308 1048
rect 246941 990 266308 992
rect 246941 987 247007 990
rect 266302 988 266308 990
rect 266372 988 266378 1052
rect 272198 990 272504 1050
rect 144729 912 205466 914
rect 144729 856 144734 912
rect 144790 856 205466 912
rect 144729 854 205466 856
rect 144729 851 144795 854
rect 205582 852 205588 916
rect 205652 914 205658 916
rect 205817 914 205883 917
rect 205652 912 205883 914
rect 205652 856 205822 912
rect 205878 856 205883 912
rect 205652 854 205883 856
rect 205652 852 205658 854
rect 205817 851 205883 854
rect 206318 852 206324 916
rect 206388 914 206394 916
rect 206553 914 206619 917
rect 206388 912 206619 914
rect 206388 856 206558 912
rect 206614 856 206619 912
rect 206388 854 206619 856
rect 206388 852 206394 854
rect 206553 851 206619 854
rect 207054 852 207060 916
rect 207124 914 207130 916
rect 207657 914 207723 917
rect 207124 912 207723 914
rect 207124 856 207662 912
rect 207718 856 207723 912
rect 207124 854 207723 856
rect 207124 852 207130 854
rect 207657 851 207723 854
rect 208526 852 208532 916
rect 208596 914 208602 916
rect 208945 914 209011 917
rect 208596 912 209011 914
rect 208596 856 208950 912
rect 209006 856 209011 912
rect 208596 854 209011 856
rect 209730 914 209790 987
rect 242893 914 242959 917
rect 209730 912 242959 914
rect 209730 856 242898 912
rect 242954 856 242959 912
rect 209730 854 242959 856
rect 208596 852 208602 854
rect 208945 851 209011 854
rect 242893 851 242959 854
rect 243537 914 243603 917
rect 260465 914 260531 917
rect 243537 912 260531 914
rect 243537 856 243542 912
rect 243598 856 260470 912
rect 260526 856 260531 912
rect 243537 854 260531 856
rect 243537 851 243603 854
rect 260465 851 260531 854
rect 267917 914 267983 917
rect 271965 914 272031 917
rect 267917 912 272031 914
rect 267917 856 267922 912
rect 267978 856 271970 912
rect 272026 856 272031 912
rect 267917 854 272031 856
rect 267917 851 267983 854
rect 271965 851 272031 854
rect 138841 780 138907 781
rect 141785 780 141851 781
rect 138790 778 138796 780
rect 138750 718 138796 778
rect 138860 776 138907 780
rect 141734 778 141740 780
rect 138902 720 138907 776
rect 138790 716 138796 718
rect 138860 716 138907 720
rect 141694 718 141740 778
rect 141804 776 141851 780
rect 141846 720 141851 776
rect 141734 716 141740 718
rect 141804 716 141851 720
rect 142470 716 142476 780
rect 142540 778 142546 780
rect 144913 778 144979 781
rect 142540 776 144979 778
rect 142540 720 144918 776
rect 144974 720 144979 776
rect 142540 718 144979 720
rect 142540 716 142546 718
rect 138841 715 138907 716
rect 141785 715 141851 716
rect 144913 715 144979 718
rect 146150 716 146156 780
rect 146220 778 146226 780
rect 147673 778 147739 781
rect 148409 780 148475 781
rect 148358 778 148364 780
rect 146220 776 147739 778
rect 146220 720 147678 776
rect 147734 720 147739 776
rect 146220 718 147739 720
rect 148318 718 148364 778
rect 148428 776 148475 780
rect 148470 720 148475 776
rect 146220 716 146226 718
rect 147673 715 147739 718
rect 148358 716 148364 718
rect 148428 716 148475 720
rect 149830 716 149836 780
rect 149900 778 149906 780
rect 150433 778 150499 781
rect 149900 776 150499 778
rect 149900 720 150438 776
rect 150494 720 150499 776
rect 149900 718 150499 720
rect 149900 716 149906 718
rect 148409 715 148475 716
rect 150433 715 150499 718
rect 151854 716 151860 780
rect 151924 778 151930 780
rect 160369 778 160435 781
rect 151924 776 160435 778
rect 151924 720 160374 776
rect 160430 720 160435 776
rect 151924 718 160435 720
rect 151924 716 151930 718
rect 160369 715 160435 718
rect 160553 778 160619 781
rect 160553 776 215770 778
rect 160553 720 160558 776
rect 160614 720 215770 776
rect 160553 718 215770 720
rect 160553 715 160619 718
rect 104065 640 122850 642
rect 104065 584 104070 640
rect 104126 584 122850 640
rect 104065 582 122850 584
rect 124397 642 124463 645
rect 125317 644 125383 645
rect 124530 642 124536 644
rect 124397 640 124536 642
rect 124397 584 124402 640
rect 124458 584 124536 640
rect 124397 582 124536 584
rect 104065 579 104131 582
rect 124397 579 124463 582
rect 124530 580 124536 582
rect 124600 580 124606 644
rect 125266 642 125272 644
rect 125226 582 125272 642
rect 125336 640 125383 644
rect 125378 584 125383 640
rect 125266 580 125272 582
rect 125336 580 125383 584
rect 126002 580 126008 644
rect 126072 642 126078 644
rect 126237 642 126303 645
rect 126072 640 126303 642
rect 126072 584 126242 640
rect 126298 584 126303 640
rect 126072 582 126303 584
rect 126072 580 126078 582
rect 125317 579 125383 580
rect 126237 579 126303 582
rect 128946 580 128952 644
rect 129016 642 129022 644
rect 129181 642 129247 645
rect 129016 640 129247 642
rect 129016 584 129186 640
rect 129242 584 129247 640
rect 129016 582 129247 584
rect 129016 580 129022 582
rect 129181 579 129247 582
rect 130418 580 130424 644
rect 130488 642 130494 644
rect 130837 642 130903 645
rect 130488 640 130903 642
rect 130488 584 130842 640
rect 130898 584 130903 640
rect 130488 582 130903 584
rect 130488 580 130494 582
rect 130837 579 130903 582
rect 131154 580 131160 644
rect 131224 642 131230 644
rect 131665 642 131731 645
rect 131224 640 131731 642
rect 131224 584 131670 640
rect 131726 584 131731 640
rect 131224 582 131731 584
rect 131224 580 131230 582
rect 131665 579 131731 582
rect 134098 580 134104 644
rect 134168 642 134174 644
rect 134517 642 134583 645
rect 134168 640 134583 642
rect 134168 584 134522 640
rect 134578 584 134583 640
rect 134168 582 134583 584
rect 134168 580 134174 582
rect 134517 579 134583 582
rect 138054 580 138060 644
rect 138124 642 138130 644
rect 138749 642 138815 645
rect 138124 640 138815 642
rect 138124 584 138754 640
rect 138810 584 138815 640
rect 138124 582 138815 584
rect 138124 580 138130 582
rect 138749 579 138815 582
rect 143206 580 143212 644
rect 143276 642 143282 644
rect 144913 642 144979 645
rect 143276 640 144979 642
rect 143276 584 144918 640
rect 144974 584 144979 640
rect 143276 582 144979 584
rect 143276 580 143282 582
rect 144913 579 144979 582
rect 147622 580 147628 644
rect 147692 642 147698 644
rect 147857 642 147923 645
rect 147692 640 147923 642
rect 147692 584 147862 640
rect 147918 584 147923 640
rect 147692 582 147923 584
rect 147692 580 147698 582
rect 147857 579 147923 582
rect 151302 580 151308 644
rect 151372 642 151378 644
rect 154113 642 154179 645
rect 151372 640 154179 642
rect 151372 584 154118 640
rect 154174 584 154179 640
rect 151372 582 154179 584
rect 151372 580 151378 582
rect 154113 579 154179 582
rect 159398 580 159404 644
rect 159468 642 159474 644
rect 160093 642 160159 645
rect 159468 640 160159 642
rect 159468 584 160098 640
rect 160154 584 160159 640
rect 159468 582 160159 584
rect 159468 580 159474 582
rect 160093 579 160159 582
rect 162117 642 162183 645
rect 162342 642 162348 644
rect 162117 640 162348 642
rect 162117 584 162122 640
rect 162178 584 162348 640
rect 162117 582 162348 584
rect 162117 579 162183 582
rect 162342 580 162348 582
rect 162412 580 162418 644
rect 163078 580 163084 644
rect 163148 642 163154 644
rect 163497 642 163563 645
rect 164601 644 164667 645
rect 169017 644 169083 645
rect 164550 642 164556 644
rect 163148 640 163563 642
rect 163148 584 163502 640
rect 163558 584 163563 640
rect 163148 582 163563 584
rect 164510 582 164556 642
rect 164620 640 164667 644
rect 168966 642 168972 644
rect 164662 584 164667 640
rect 163148 580 163154 582
rect 163497 579 163563 582
rect 164550 580 164556 582
rect 164620 580 164667 584
rect 168926 582 168972 642
rect 169036 640 169083 644
rect 169078 584 169083 640
rect 168966 580 168972 582
rect 169036 580 169083 584
rect 171450 580 171456 644
rect 171520 642 171526 644
rect 171685 642 171751 645
rect 172237 644 172303 645
rect 172973 644 173039 645
rect 172186 642 172192 644
rect 171520 640 171751 642
rect 171520 584 171690 640
rect 171746 584 171751 640
rect 171520 582 171751 584
rect 172146 582 172192 642
rect 172256 640 172303 644
rect 172922 642 172928 644
rect 172298 584 172303 640
rect 171520 580 171526 582
rect 164601 579 164667 580
rect 169017 579 169083 580
rect 171685 579 171751 582
rect 172186 580 172192 582
rect 172256 580 172303 584
rect 172882 582 172928 642
rect 172992 640 173039 644
rect 173034 584 173039 640
rect 172922 580 172928 582
rect 172992 580 173039 584
rect 173658 580 173664 644
rect 173728 642 173734 644
rect 173893 642 173959 645
rect 174445 644 174511 645
rect 174394 642 174400 644
rect 173728 640 173959 642
rect 173728 584 173898 640
rect 173954 584 173959 640
rect 173728 582 173959 584
rect 174354 582 174400 642
rect 174464 640 174511 644
rect 174506 584 174511 640
rect 173728 580 173734 582
rect 172237 579 172303 580
rect 172973 579 173039 580
rect 173893 579 173959 582
rect 174394 580 174400 582
rect 174464 580 174511 584
rect 175130 580 175136 644
rect 175200 642 175206 644
rect 175273 642 175339 645
rect 176653 644 176719 645
rect 176602 642 176608 644
rect 175200 640 175339 642
rect 175200 584 175278 640
rect 175334 584 175339 640
rect 175200 582 175339 584
rect 176562 582 176608 642
rect 176672 640 176719 644
rect 176714 584 176719 640
rect 175200 580 175206 582
rect 174445 579 174511 580
rect 175273 579 175339 582
rect 176602 580 176608 582
rect 176672 580 176719 584
rect 177338 580 177344 644
rect 177408 642 177414 644
rect 177849 642 177915 645
rect 177408 640 177915 642
rect 177408 584 177854 640
rect 177910 584 177915 640
rect 177408 582 177915 584
rect 177408 580 177414 582
rect 176653 579 176719 580
rect 177849 579 177915 582
rect 178074 580 178080 644
rect 178144 642 178150 644
rect 178493 642 178559 645
rect 178144 640 178559 642
rect 178144 584 178498 640
rect 178554 584 178559 640
rect 178144 582 178559 584
rect 178144 580 178150 582
rect 178493 579 178559 582
rect 178810 580 178816 644
rect 178880 642 178886 644
rect 179137 642 179203 645
rect 179597 644 179663 645
rect 180333 644 180399 645
rect 179546 642 179552 644
rect 178880 640 179203 642
rect 178880 584 179142 640
rect 179198 584 179203 640
rect 178880 582 179203 584
rect 179506 582 179552 642
rect 179616 640 179663 644
rect 180282 642 180288 644
rect 179658 584 179663 640
rect 178880 580 178886 582
rect 179137 579 179203 582
rect 179546 580 179552 582
rect 179616 580 179663 584
rect 180242 582 180288 642
rect 180352 640 180399 644
rect 180394 584 180399 640
rect 180282 580 180288 582
rect 180352 580 180399 584
rect 179597 579 179663 580
rect 180333 579 180399 580
rect 180517 642 180583 645
rect 215569 642 215635 645
rect 180517 640 215635 642
rect 180517 584 180522 640
rect 180578 584 215574 640
rect 215630 584 215635 640
rect 180517 582 215635 584
rect 215710 642 215770 718
rect 215886 716 215892 780
rect 215956 778 215962 780
rect 218053 778 218119 781
rect 223573 778 223639 781
rect 224769 780 224835 781
rect 224718 778 224724 780
rect 215956 776 218119 778
rect 215956 720 218058 776
rect 218114 720 218119 776
rect 215956 718 218119 720
rect 215956 716 215962 718
rect 218053 715 218119 718
rect 220126 776 223639 778
rect 220126 720 223578 776
rect 223634 720 223639 776
rect 220126 718 223639 720
rect 224678 718 224724 778
rect 224788 776 224835 780
rect 224830 720 224835 776
rect 219157 642 219223 645
rect 220126 642 220186 718
rect 223573 715 223639 718
rect 224718 716 224724 718
rect 224788 716 224835 720
rect 225086 716 225092 780
rect 225156 778 225162 780
rect 248505 778 248571 781
rect 260097 778 260163 781
rect 225156 776 248571 778
rect 225156 720 248510 776
rect 248566 720 248571 776
rect 225156 718 248571 720
rect 225156 716 225162 718
rect 224769 715 224835 716
rect 248505 715 248571 718
rect 249014 776 260163 778
rect 249014 720 260102 776
rect 260158 720 260163 776
rect 249014 718 260163 720
rect 215710 640 219223 642
rect 215710 584 219162 640
rect 219218 584 219223 640
rect 215710 582 219223 584
rect 180517 579 180583 582
rect 215569 579 215635 582
rect 219157 579 219223 582
rect 219390 582 220186 642
rect 39849 504 55230 506
rect 39849 448 39854 504
rect 39910 448 55230 504
rect 39849 446 55230 448
rect 39849 443 39915 446
rect 55530 444 55536 508
rect 55600 506 55606 508
rect 55673 506 55739 509
rect 55600 504 55739 506
rect 55600 448 55678 504
rect 55734 448 55739 504
rect 55600 446 55739 448
rect 55600 444 55606 446
rect 55673 443 55739 446
rect 56266 444 56272 508
rect 56336 506 56342 508
rect 56409 506 56475 509
rect 56336 504 56475 506
rect 56336 448 56414 504
rect 56470 448 56475 504
rect 56336 446 56475 448
rect 56336 444 56342 446
rect 56409 443 56475 446
rect 57002 444 57008 508
rect 57072 506 57078 508
rect 57145 506 57211 509
rect 57072 504 57211 506
rect 57072 448 57150 504
rect 57206 448 57211 504
rect 57072 446 57211 448
rect 57072 444 57078 446
rect 57145 443 57211 446
rect 58249 506 58315 509
rect 59997 508 60063 509
rect 58474 506 58480 508
rect 58249 504 58480 506
rect 58249 448 58254 504
rect 58310 448 58480 504
rect 58249 446 58480 448
rect 58249 443 58315 446
rect 58474 444 58480 446
rect 58544 444 58550 508
rect 59946 506 59952 508
rect 59906 446 59952 506
rect 60016 504 60063 508
rect 60058 448 60063 504
rect 59946 444 59952 446
rect 60016 444 60063 448
rect 60682 444 60688 508
rect 60752 506 60758 508
rect 60917 506 60983 509
rect 61469 508 61535 509
rect 61418 506 61424 508
rect 60752 504 60983 506
rect 60752 448 60922 504
rect 60978 448 60983 504
rect 60752 446 60983 448
rect 61378 446 61424 506
rect 61488 504 61535 508
rect 61530 448 61535 504
rect 60752 444 60758 446
rect 59997 443 60063 444
rect 60917 443 60983 446
rect 61418 444 61424 446
rect 61488 444 61535 448
rect 62154 444 62160 508
rect 62224 506 62230 508
rect 62389 506 62455 509
rect 62224 504 62455 506
rect 62224 448 62394 504
rect 62450 448 62455 504
rect 62224 446 62455 448
rect 62224 444 62230 446
rect 61469 443 61535 444
rect 62389 443 62455 446
rect 62890 444 62896 508
rect 62960 506 62966 508
rect 63125 506 63191 509
rect 65885 508 65951 509
rect 65834 506 65840 508
rect 62960 504 63191 506
rect 62960 448 63130 504
rect 63186 448 63191 504
rect 62960 446 63191 448
rect 65794 446 65840 506
rect 65904 504 65951 508
rect 65946 448 65951 504
rect 62960 444 62966 446
rect 63125 443 63191 446
rect 65834 444 65840 446
rect 65904 444 65951 448
rect 66570 444 66576 508
rect 66640 506 66646 508
rect 67265 506 67331 509
rect 87505 508 87571 509
rect 87454 506 87460 508
rect 66640 504 67331 506
rect 66640 448 67270 504
rect 67326 448 67331 504
rect 66640 446 67331 448
rect 87414 446 87460 506
rect 87524 504 87571 508
rect 117773 506 117839 509
rect 87566 448 87571 504
rect 66640 444 66646 446
rect 65885 443 65951 444
rect 67265 443 67331 446
rect 87454 444 87460 446
rect 87524 444 87571 448
rect 87505 443 87571 444
rect 89670 504 117839 506
rect 89670 448 117778 504
rect 117834 448 117839 504
rect 89670 446 117839 448
rect 8385 370 8451 373
rect 8886 370 8892 372
rect 8385 368 8892 370
rect 8385 312 8390 368
rect 8446 312 8892 368
rect 8385 310 8892 312
rect 8385 307 8451 310
rect 8886 308 8892 310
rect 8956 308 8962 372
rect 18454 308 18460 372
rect 18524 370 18530 372
rect 18597 370 18663 373
rect 28809 372 28875 373
rect 28758 370 28764 372
rect 18524 368 18663 370
rect 18524 312 18602 368
rect 18658 312 18663 368
rect 18524 310 18663 312
rect 28718 310 28764 370
rect 28828 368 28875 372
rect 28870 312 28875 368
rect 18524 308 18530 310
rect 18597 307 18663 310
rect 28758 308 28764 310
rect 28828 308 28875 312
rect 28809 307 28875 308
rect 38837 370 38903 373
rect 39338 370 39344 372
rect 38837 368 39344 370
rect 38837 312 38842 368
rect 38898 312 39344 368
rect 38837 310 39344 312
rect 38837 307 38903 310
rect 39338 308 39344 310
rect 39408 308 39414 372
rect 52586 308 52592 372
rect 52656 370 52662 372
rect 53097 370 53163 373
rect 52656 368 53163 370
rect 52656 312 53102 368
rect 53158 312 53163 368
rect 52656 310 53163 312
rect 52656 308 52662 310
rect 53097 307 53163 310
rect 63626 308 63632 372
rect 63696 370 63702 372
rect 63861 370 63927 373
rect 63696 368 63927 370
rect 63696 312 63866 368
rect 63922 312 63927 368
rect 63696 310 63927 312
rect 63696 308 63702 310
rect 63861 307 63927 310
rect 64362 308 64368 372
rect 64432 370 64438 372
rect 64597 370 64663 373
rect 64432 368 64663 370
rect 64432 312 64602 368
rect 64658 312 64663 368
rect 64432 310 64663 312
rect 64432 308 64438 310
rect 64597 307 64663 310
rect 65098 308 65104 372
rect 65168 370 65174 372
rect 65977 370 66043 373
rect 65168 368 66043 370
rect 65168 312 65982 368
rect 66038 312 66043 368
rect 65168 310 66043 312
rect 65168 308 65174 310
rect 65977 307 66043 310
rect 85021 370 85087 373
rect 85246 370 85252 372
rect 85021 368 85252 370
rect 85021 312 85026 368
rect 85082 312 85252 368
rect 85021 310 85252 312
rect 85021 307 85087 310
rect 85246 308 85252 310
rect 85316 308 85322 372
rect 85481 370 85547 373
rect 89670 370 89730 446
rect 117773 443 117839 446
rect 117906 444 117912 508
rect 117976 506 117982 508
rect 118049 506 118115 509
rect 118693 508 118759 509
rect 118642 506 118648 508
rect 117976 504 118115 506
rect 117976 448 118054 504
rect 118110 448 118115 504
rect 117976 446 118115 448
rect 118606 446 118648 506
rect 118712 504 118759 508
rect 118754 448 118759 504
rect 117976 444 117982 446
rect 118049 443 118115 446
rect 118642 444 118648 446
rect 118712 444 118759 448
rect 118693 443 118759 444
rect 119337 508 119403 509
rect 119337 504 119384 508
rect 119448 506 119454 508
rect 119337 448 119342 504
rect 119337 444 119384 448
rect 119448 446 119494 506
rect 119448 444 119454 446
rect 120114 444 120120 508
rect 120184 506 120190 508
rect 120349 506 120415 509
rect 120184 504 120415 506
rect 120184 448 120354 504
rect 120410 448 120415 504
rect 120184 446 120415 448
rect 120184 444 120190 446
rect 119337 443 119403 444
rect 120349 443 120415 446
rect 120850 444 120856 508
rect 120920 506 120926 508
rect 121085 506 121151 509
rect 120920 504 121151 506
rect 120920 448 121090 504
rect 121146 448 121151 504
rect 120920 446 121151 448
rect 120920 444 120926 446
rect 121085 443 121151 446
rect 121586 444 121592 508
rect 121656 506 121662 508
rect 121821 506 121887 509
rect 121656 504 121887 506
rect 121656 448 121826 504
rect 121882 448 121887 504
rect 121656 446 121887 448
rect 121656 444 121662 446
rect 121821 443 121887 446
rect 122322 444 122328 508
rect 122392 506 122398 508
rect 122649 506 122715 509
rect 122392 504 122715 506
rect 122392 448 122654 504
rect 122710 448 122715 504
rect 122392 446 122715 448
rect 122392 444 122398 446
rect 122649 443 122715 446
rect 123058 444 123064 508
rect 123128 506 123134 508
rect 123385 506 123451 509
rect 123128 504 123451 506
rect 123128 448 123390 504
rect 123446 448 123451 504
rect 123128 446 123451 448
rect 123128 444 123134 446
rect 123385 443 123451 446
rect 127474 444 127480 508
rect 127544 506 127550 508
rect 127801 506 127867 509
rect 143993 508 144059 509
rect 143942 506 143948 508
rect 127544 504 127867 506
rect 127544 448 127806 504
rect 127862 448 127867 504
rect 127544 446 127867 448
rect 143902 446 143948 506
rect 144012 504 144059 508
rect 144054 448 144059 504
rect 127544 444 127550 446
rect 127801 443 127867 446
rect 143942 444 143948 446
rect 144012 444 144059 448
rect 143993 443 144059 444
rect 144502 446 174002 506
rect 85481 368 89730 370
rect 85481 312 85486 368
rect 85542 312 89730 368
rect 85481 310 89730 312
rect 85481 307 85547 310
rect 95182 308 95188 372
rect 95252 370 95258 372
rect 103513 370 103579 373
rect 95252 368 103579 370
rect 95252 312 103518 368
rect 103574 312 103579 368
rect 95252 310 103579 312
rect 95252 308 95258 310
rect 103513 307 103579 310
rect 129682 308 129688 372
rect 129752 370 129758 372
rect 130745 370 130811 373
rect 129752 368 130811 370
rect 129752 312 130750 368
rect 130806 312 130811 368
rect 129752 310 130811 312
rect 129752 308 129758 310
rect 130745 307 130811 310
rect 131890 308 131896 372
rect 131960 370 131966 372
rect 132125 370 132191 373
rect 131960 368 132191 370
rect 131960 312 132130 368
rect 132186 312 132191 368
rect 131960 310 132191 312
rect 131960 308 131966 310
rect 132125 307 132191 310
rect 132626 308 132632 372
rect 132696 370 132702 372
rect 133229 370 133295 373
rect 132696 368 133295 370
rect 132696 312 133234 368
rect 133290 312 133295 368
rect 132696 310 133295 312
rect 132696 308 132702 310
rect 133229 307 133295 310
rect 141417 370 141483 373
rect 144502 370 144562 446
rect 146937 372 147003 373
rect 146886 370 146892 372
rect 141417 368 144562 370
rect 141417 312 141422 368
rect 141478 312 144562 368
rect 141417 310 144562 312
rect 146846 310 146892 370
rect 146956 368 147003 372
rect 146998 312 147003 368
rect 141417 307 141483 310
rect 146886 308 146892 310
rect 146956 308 147003 312
rect 146937 307 147003 308
rect 147630 310 160754 370
rect 94313 234 94379 237
rect 104157 234 104223 237
rect 94313 232 104223 234
rect 94313 176 94318 232
rect 94374 176 104162 232
rect 104218 176 104223 232
rect 94313 174 104223 176
rect 94313 171 94379 174
rect 104157 171 104223 174
rect 140313 234 140379 237
rect 147630 234 147690 310
rect 140313 232 147690 234
rect 140313 176 140318 232
rect 140374 176 147690 232
rect 140313 174 147690 176
rect 140313 171 140379 174
rect 153142 172 153148 236
rect 153212 234 153218 236
rect 160553 234 160619 237
rect 153212 232 160619 234
rect 153212 176 160558 232
rect 160614 176 160619 232
rect 153212 174 160619 176
rect 160694 234 160754 310
rect 160870 308 160876 372
rect 160940 370 160946 372
rect 161289 370 161355 373
rect 160940 368 161355 370
rect 160940 312 161294 368
rect 161350 312 161355 368
rect 160940 310 161355 312
rect 160940 308 160946 310
rect 161289 307 161355 310
rect 167494 308 167500 372
rect 167564 370 167570 372
rect 167913 370 167979 373
rect 167564 368 167979 370
rect 167564 312 167918 368
rect 167974 312 167979 368
rect 167564 310 167979 312
rect 173942 370 174002 446
rect 175866 444 175872 508
rect 175936 506 175942 508
rect 176561 506 176627 509
rect 181805 508 181871 509
rect 181754 506 181760 508
rect 175936 504 176627 506
rect 175936 448 176566 504
rect 176622 448 176627 504
rect 175936 446 176627 448
rect 181714 446 181760 506
rect 181824 504 181871 508
rect 181866 448 181871 504
rect 175936 444 175942 446
rect 176561 443 176627 446
rect 181754 444 181760 446
rect 181824 444 181871 448
rect 182490 444 182496 508
rect 182560 506 182566 508
rect 183001 506 183067 509
rect 183277 508 183343 509
rect 183226 506 183232 508
rect 182560 504 183067 506
rect 182560 448 183006 504
rect 183062 448 183067 504
rect 182560 446 183067 448
rect 183186 446 183232 506
rect 183296 504 183343 508
rect 183338 448 183343 504
rect 182560 444 182566 446
rect 181805 443 181871 444
rect 183001 443 183067 446
rect 183226 444 183232 446
rect 183296 444 183343 448
rect 183962 444 183968 508
rect 184032 506 184038 508
rect 184289 506 184355 509
rect 184749 508 184815 509
rect 185485 508 185551 509
rect 186957 508 187023 509
rect 184698 506 184704 508
rect 184032 504 184355 506
rect 184032 448 184294 504
rect 184350 448 184355 504
rect 184032 446 184355 448
rect 184658 446 184704 506
rect 184768 504 184815 508
rect 185434 506 185440 508
rect 184810 448 184815 504
rect 184032 444 184038 446
rect 183277 443 183343 444
rect 184289 443 184355 446
rect 184698 444 184704 446
rect 184768 444 184815 448
rect 185394 446 185440 506
rect 185504 504 185551 508
rect 186906 506 186912 508
rect 185546 448 185551 504
rect 185434 444 185440 446
rect 185504 444 185551 448
rect 186866 446 186912 506
rect 186976 504 187023 508
rect 187018 448 187023 504
rect 186906 444 186912 446
rect 186976 444 187023 448
rect 187642 444 187648 508
rect 187712 506 187718 508
rect 188153 506 188219 509
rect 187712 504 188219 506
rect 187712 448 188158 504
rect 188214 448 188219 504
rect 187712 446 188219 448
rect 187712 444 187718 446
rect 184749 443 184815 444
rect 185485 443 185551 444
rect 186957 443 187023 444
rect 188153 443 188219 446
rect 188378 444 188384 508
rect 188448 506 188454 508
rect 188613 506 188679 509
rect 188448 504 188679 506
rect 188448 448 188618 504
rect 188674 448 188679 504
rect 188448 446 188679 448
rect 188448 444 188454 446
rect 188613 443 188679 446
rect 189114 444 189120 508
rect 189184 506 189190 508
rect 189441 506 189507 509
rect 189184 504 189507 506
rect 189184 448 189446 504
rect 189502 448 189507 504
rect 189184 446 189507 448
rect 189184 444 189190 446
rect 189441 443 189507 446
rect 190586 444 190592 508
rect 190656 506 190662 508
rect 191097 506 191163 509
rect 192845 508 192911 509
rect 193581 508 193647 509
rect 192794 506 192800 508
rect 190656 504 191163 506
rect 190656 448 191102 504
rect 191158 448 191163 504
rect 190656 446 191163 448
rect 192754 446 192800 506
rect 192864 504 192911 508
rect 193530 506 193536 508
rect 192906 448 192911 504
rect 190656 444 190662 446
rect 191097 443 191163 446
rect 192794 444 192800 446
rect 192864 444 192911 448
rect 193490 446 193536 506
rect 193600 504 193647 508
rect 193642 448 193647 504
rect 193530 444 193536 446
rect 193600 444 193647 448
rect 195002 444 195008 508
rect 195072 506 195078 508
rect 195605 506 195671 509
rect 195072 504 195671 506
rect 195072 448 195610 504
rect 195666 448 195671 504
rect 195072 446 195671 448
rect 195072 444 195078 446
rect 192845 443 192911 444
rect 193581 443 193647 444
rect 195605 443 195671 446
rect 196474 444 196480 508
rect 196544 506 196550 508
rect 196617 506 196683 509
rect 196544 504 196683 506
rect 196544 448 196622 504
rect 196678 448 196683 504
rect 196544 446 196683 448
rect 196544 444 196550 446
rect 196617 443 196683 446
rect 198682 444 198688 508
rect 198752 506 198758 508
rect 199929 506 199995 509
rect 198752 504 199995 506
rect 198752 448 199934 504
rect 199990 448 199995 504
rect 198752 446 199995 448
rect 198752 444 198758 446
rect 199929 443 199995 446
rect 200154 444 200160 508
rect 200224 506 200230 508
rect 201217 506 201283 509
rect 202413 508 202479 509
rect 202362 506 202368 508
rect 200224 504 201283 506
rect 200224 448 201222 504
rect 201278 448 201283 504
rect 200224 446 201283 448
rect 202322 446 202368 506
rect 202432 504 202479 508
rect 202474 448 202479 504
rect 200224 444 200230 446
rect 201217 443 201283 446
rect 202362 444 202368 446
rect 202432 444 202479 448
rect 203098 444 203104 508
rect 203168 506 203174 508
rect 204069 506 204135 509
rect 203168 504 204135 506
rect 203168 448 204074 504
rect 204130 448 204135 504
rect 203168 446 204135 448
rect 203168 444 203174 446
rect 202413 443 202479 444
rect 204069 443 204135 446
rect 208485 506 208551 509
rect 209262 506 209268 508
rect 208485 504 209268 506
rect 208485 448 208490 504
rect 208546 448 209268 504
rect 208485 446 209268 448
rect 208485 443 208551 446
rect 209262 444 209268 446
rect 209332 444 209338 508
rect 213678 444 213684 508
rect 213748 506 213754 508
rect 216673 506 216739 509
rect 213748 504 216739 506
rect 213748 448 216678 504
rect 216734 448 216739 504
rect 213748 446 216739 448
rect 213748 444 213754 446
rect 216673 443 216739 446
rect 176837 370 176903 373
rect 173942 368 176903 370
rect 173942 312 176842 368
rect 176898 312 176903 368
rect 173942 310 176903 312
rect 167564 308 167570 310
rect 167913 307 167979 310
rect 176837 307 176903 310
rect 181018 308 181024 372
rect 181088 370 181094 372
rect 181713 370 181779 373
rect 181088 368 181779 370
rect 181088 312 181718 368
rect 181774 312 181779 368
rect 181088 310 181779 312
rect 181088 308 181094 310
rect 181713 307 181779 310
rect 192058 308 192064 372
rect 192128 370 192134 372
rect 192569 370 192635 373
rect 192128 368 192635 370
rect 192128 312 192574 368
rect 192630 312 192635 368
rect 192128 310 192635 312
rect 192128 308 192134 310
rect 192569 307 192635 310
rect 207790 308 207796 372
rect 207860 370 207866 372
rect 208301 370 208367 373
rect 212993 372 213059 373
rect 214465 372 214531 373
rect 212942 370 212948 372
rect 207860 368 208367 370
rect 207860 312 208306 368
rect 208362 312 208367 368
rect 207860 310 208367 312
rect 212902 310 212948 370
rect 213012 368 213059 372
rect 214414 370 214420 372
rect 213054 312 213059 368
rect 207860 308 207866 310
rect 208301 307 208367 310
rect 212942 308 212948 310
rect 213012 308 213059 312
rect 214374 310 214420 370
rect 214484 368 214531 372
rect 214526 312 214531 368
rect 214414 308 214420 310
rect 214484 308 214531 312
rect 212993 307 213059 308
rect 214465 307 214531 308
rect 215569 370 215635 373
rect 219390 370 219450 582
rect 221774 580 221780 644
rect 221844 642 221850 644
rect 225965 642 226031 645
rect 221844 640 226031 642
rect 221844 584 225970 640
rect 226026 584 226031 640
rect 221844 582 226031 584
rect 221844 580 221850 582
rect 225965 579 226031 582
rect 226926 580 226932 644
rect 226996 642 227002 644
rect 227437 642 227503 645
rect 226996 640 227503 642
rect 226996 584 227442 640
rect 227498 584 227503 640
rect 226996 582 227503 584
rect 226996 580 227002 582
rect 227437 579 227503 582
rect 228398 580 228404 644
rect 228468 642 228474 644
rect 228725 642 228791 645
rect 228468 640 228791 642
rect 228468 584 228730 640
rect 228786 584 228791 640
rect 228468 582 228791 584
rect 228468 580 228474 582
rect 228725 579 228791 582
rect 229134 580 229140 644
rect 229204 642 229210 644
rect 229461 642 229527 645
rect 229204 640 229527 642
rect 229204 584 229466 640
rect 229522 584 229527 640
rect 229204 582 229527 584
rect 229204 580 229210 582
rect 229461 579 229527 582
rect 231342 580 231348 644
rect 231412 642 231418 644
rect 231853 642 231919 645
rect 231412 640 231919 642
rect 231412 584 231858 640
rect 231914 584 231919 640
rect 231412 582 231919 584
rect 231412 580 231418 582
rect 231853 579 231919 582
rect 233550 580 233556 644
rect 233620 642 233626 644
rect 233877 642 233943 645
rect 233620 640 233943 642
rect 233620 584 233882 640
rect 233938 584 233943 640
rect 233620 582 233943 584
rect 233620 580 233626 582
rect 233877 579 233943 582
rect 234286 580 234292 644
rect 234356 642 234362 644
rect 234613 642 234679 645
rect 235809 644 235875 645
rect 235758 642 235764 644
rect 234356 640 234679 642
rect 234356 584 234618 640
rect 234674 584 234679 640
rect 234356 582 234679 584
rect 235718 582 235764 642
rect 235828 640 235875 644
rect 235870 584 235875 640
rect 234356 580 234362 582
rect 234613 579 234679 582
rect 235758 580 235764 582
rect 235828 580 235875 584
rect 239714 580 239720 644
rect 239784 642 239790 644
rect 239949 642 240015 645
rect 239784 640 240015 642
rect 239784 584 239954 640
rect 240010 584 240015 640
rect 239784 582 240015 584
rect 239784 580 239790 582
rect 235809 579 235875 580
rect 239949 579 240015 582
rect 240450 580 240456 644
rect 240520 642 240526 644
rect 240961 642 241027 645
rect 241237 644 241303 645
rect 241973 644 242039 645
rect 243445 644 243511 645
rect 244181 644 244247 645
rect 244917 644 244983 645
rect 241186 642 241192 644
rect 240520 640 241027 642
rect 240520 584 240966 640
rect 241022 584 241027 640
rect 240520 582 241027 584
rect 241146 582 241192 642
rect 241256 640 241303 644
rect 241922 642 241928 644
rect 241298 584 241303 640
rect 240520 580 240526 582
rect 240961 579 241027 582
rect 241186 580 241192 582
rect 241256 580 241303 584
rect 241882 582 241928 642
rect 241992 640 242039 644
rect 243394 642 243400 644
rect 242034 584 242039 640
rect 241922 580 241928 582
rect 241992 580 242039 584
rect 243354 582 243400 642
rect 243464 640 243511 644
rect 244130 642 244136 644
rect 243506 584 243511 640
rect 243394 580 243400 582
rect 243464 580 243511 584
rect 244090 582 244136 642
rect 244200 640 244247 644
rect 244866 642 244872 644
rect 244242 584 244247 640
rect 244130 580 244136 582
rect 244200 580 244247 584
rect 244826 582 244872 642
rect 244936 640 244983 644
rect 244978 584 244983 640
rect 244866 580 244872 582
rect 244936 580 244983 584
rect 241237 579 241303 580
rect 241973 579 242039 580
rect 243445 579 243511 580
rect 244181 579 244247 580
rect 244917 579 244983 580
rect 247033 644 247099 645
rect 247033 640 247080 644
rect 247144 642 247150 644
rect 247033 584 247038 640
rect 247033 580 247080 584
rect 247144 582 247190 642
rect 247144 580 247150 582
rect 247810 580 247816 644
rect 247880 642 247886 644
rect 248413 642 248479 645
rect 247880 640 248479 642
rect 247880 584 248418 640
rect 248474 584 248479 640
rect 247880 582 248479 584
rect 247880 580 247886 582
rect 247033 579 247099 580
rect 248413 579 248479 582
rect 230197 506 230263 509
rect 215569 368 219450 370
rect 215569 312 215574 368
rect 215630 312 219450 368
rect 215569 310 219450 312
rect 220126 504 230263 506
rect 220126 448 230202 504
rect 230258 448 230263 504
rect 220126 446 230263 448
rect 215569 307 215635 310
rect 174261 234 174327 237
rect 160694 232 174327 234
rect 160694 176 174266 232
rect 174322 176 174327 232
rect 160694 174 174327 176
rect 153212 172 153218 174
rect 160553 171 160619 174
rect 174261 171 174327 174
rect 210969 234 211035 237
rect 220126 234 220186 446
rect 230197 443 230263 446
rect 230381 506 230447 509
rect 249014 506 249074 718
rect 260097 715 260163 718
rect 267733 778 267799 781
rect 272198 778 272258 990
rect 267733 776 272258 778
rect 267733 720 267738 776
rect 267794 720 272258 776
rect 267733 718 272258 720
rect 267733 715 267799 718
rect 250069 644 250135 645
rect 250018 642 250024 644
rect 249978 582 250024 642
rect 250088 640 250135 644
rect 250130 584 250135 640
rect 250018 580 250024 582
rect 250088 580 250135 584
rect 254434 580 254440 644
rect 254504 642 254510 644
rect 254853 642 254919 645
rect 254504 640 254919 642
rect 254504 584 254858 640
rect 254914 584 254919 640
rect 254504 582 254919 584
rect 254504 580 254510 582
rect 250069 579 250135 580
rect 254853 579 254919 582
rect 255170 580 255176 644
rect 255240 642 255246 644
rect 256785 642 256851 645
rect 255240 640 256851 642
rect 255240 584 256790 640
rect 256846 584 256851 640
rect 255240 582 256851 584
rect 255240 580 255246 582
rect 256785 579 256851 582
rect 258073 644 258139 645
rect 261109 644 261175 645
rect 258073 640 258120 644
rect 258184 642 258190 644
rect 261058 642 261064 644
rect 258073 584 258078 640
rect 258073 580 258120 584
rect 258184 582 258230 642
rect 261018 582 261064 642
rect 261128 640 261175 644
rect 261170 584 261175 640
rect 258184 580 258190 582
rect 261058 580 261064 582
rect 261128 580 261175 584
rect 262530 580 262536 644
rect 262600 642 262606 644
rect 262857 642 262923 645
rect 263317 644 263383 645
rect 263266 642 263272 644
rect 262600 640 262923 642
rect 262600 584 262862 640
rect 262918 584 262923 640
rect 262600 582 262923 584
rect 263226 582 263272 642
rect 263336 640 263383 644
rect 263378 584 263383 640
rect 262600 580 262606 582
rect 258073 579 258139 580
rect 261109 579 261175 580
rect 262857 579 262923 582
rect 263266 580 263272 582
rect 263336 580 263383 584
rect 264002 580 264008 644
rect 264072 642 264078 644
rect 264329 642 264395 645
rect 264072 640 264395 642
rect 264072 584 264334 640
rect 264390 584 264395 640
rect 264072 582 264395 584
rect 264072 580 264078 582
rect 263317 579 263383 580
rect 264329 579 264395 582
rect 264738 580 264744 644
rect 264808 642 264814 644
rect 264973 642 265039 645
rect 264808 640 265039 642
rect 264808 584 264978 640
rect 265034 584 265039 640
rect 264808 582 265039 584
rect 264808 580 264814 582
rect 264973 579 265039 582
rect 265474 580 265480 644
rect 265544 642 265550 644
rect 265801 642 265867 645
rect 265544 640 265867 642
rect 265544 584 265806 640
rect 265862 584 265867 640
rect 265544 582 265867 584
rect 265544 580 265550 582
rect 265801 579 265867 582
rect 266210 580 266216 644
rect 266280 642 266286 644
rect 266353 642 266419 645
rect 266280 640 266419 642
rect 266280 584 266358 640
rect 266414 584 266419 640
rect 266280 582 266419 584
rect 266280 580 266286 582
rect 266353 579 266419 582
rect 266905 644 266971 645
rect 267641 644 267707 645
rect 268377 644 268443 645
rect 266905 640 266952 644
rect 267016 642 267022 644
rect 266905 584 266910 640
rect 266905 580 266952 584
rect 267016 582 267062 642
rect 267641 640 267688 644
rect 267752 642 267758 644
rect 267641 584 267646 640
rect 267016 580 267022 582
rect 267641 580 267688 584
rect 267752 582 267798 642
rect 268377 640 268424 644
rect 268488 642 268494 644
rect 268377 584 268382 640
rect 267752 580 267758 582
rect 268377 580 268424 584
rect 268488 582 268534 642
rect 268488 580 268494 582
rect 269154 580 269160 644
rect 269224 642 269230 644
rect 269757 642 269823 645
rect 269224 640 269823 642
rect 269224 584 269762 640
rect 269818 584 269823 640
rect 269224 582 269823 584
rect 269224 580 269230 582
rect 266905 579 266971 580
rect 267641 579 267707 580
rect 268377 579 268443 580
rect 269757 579 269823 582
rect 270626 580 270632 644
rect 270696 642 270702 644
rect 270769 642 270835 645
rect 270696 640 270835 642
rect 270696 584 270774 640
rect 270830 584 270835 640
rect 270696 582 270835 584
rect 270696 580 270702 582
rect 270769 579 270835 582
rect 230381 504 249074 506
rect 230381 448 230386 504
rect 230442 448 249074 504
rect 230381 446 249074 448
rect 230381 443 230447 446
rect 252962 444 252968 508
rect 253032 506 253038 508
rect 253841 506 253907 509
rect 253032 504 253907 506
rect 253032 448 253846 504
rect 253902 448 253907 504
rect 253032 446 253907 448
rect 253032 444 253038 446
rect 253841 443 253907 446
rect 220302 308 220308 372
rect 220372 370 220378 372
rect 220813 370 220879 373
rect 220372 368 220879 370
rect 220372 312 220818 368
rect 220874 312 220879 368
rect 220372 310 220879 312
rect 220372 308 220378 310
rect 220813 307 220879 310
rect 221089 370 221155 373
rect 230289 370 230355 373
rect 221089 368 230355 370
rect 221089 312 221094 368
rect 221150 312 230294 368
rect 230350 312 230355 368
rect 221089 310 230355 312
rect 221089 307 221155 310
rect 230289 307 230355 310
rect 253698 308 253704 372
rect 253768 370 253774 372
rect 255957 370 256023 373
rect 253768 368 256023 370
rect 253768 312 255962 368
rect 256018 312 256023 368
rect 253768 310 256023 312
rect 253768 308 253774 310
rect 255957 307 256023 310
rect 269890 308 269896 372
rect 269960 370 269966 372
rect 270309 370 270375 373
rect 269960 368 270375 370
rect 269960 312 270314 368
rect 270370 312 270375 368
rect 269960 310 270375 312
rect 269960 308 269966 310
rect 270309 307 270375 310
rect 210969 232 220186 234
rect 210969 176 210974 232
rect 211030 176 220186 232
rect 210969 174 220186 176
rect 230197 234 230263 237
rect 236269 234 236335 237
rect 230197 232 236335 234
rect 230197 176 230202 232
rect 230258 176 236274 232
rect 236330 176 236335 232
rect 230197 174 236335 176
rect 210969 171 211035 174
rect 230197 171 230263 174
rect 236269 171 236335 174
rect 92197 98 92263 101
rect 98269 98 98335 101
rect 92197 96 98335 98
rect 92197 40 92202 96
rect 92258 40 98274 96
rect 98330 40 98335 96
rect 92197 38 98335 40
rect 92197 35 92263 38
rect 98269 35 98335 38
rect 141233 98 141299 101
rect 160001 98 160067 101
rect 141233 96 160067 98
rect 141233 40 141238 96
rect 141294 40 160006 96
rect 160062 40 160067 96
rect 141233 38 160067 40
rect 141233 35 141299 38
rect 160001 35 160067 38
rect 213361 98 213427 101
rect 231393 98 231459 101
rect 213361 96 231459 98
rect 213361 40 213366 96
rect 213422 40 231398 96
rect 231454 40 231459 96
rect 213361 38 231459 40
rect 213361 35 213427 38
rect 231393 35 231459 38
<< via3 >>
rect 52592 10508 52656 10572
rect 81572 10568 81636 10572
rect 81572 10512 81622 10568
rect 81622 10512 81636 10568
rect 81572 10508 81636 10512
rect 82308 10508 82372 10572
rect 86724 10568 86788 10572
rect 86724 10512 86774 10568
rect 86774 10512 86788 10568
rect 86724 10508 86788 10512
rect 147628 10508 147692 10572
rect 172192 10568 172256 10572
rect 172192 10512 172242 10568
rect 172242 10512 172256 10568
rect 172192 10508 172256 10512
rect 179552 10508 179616 10572
rect 207796 10508 207860 10572
rect 212948 10508 213012 10572
rect 218100 10508 218164 10572
rect 72004 10432 72068 10436
rect 72004 10376 72054 10432
rect 72054 10376 72068 10432
rect 72004 10372 72068 10376
rect 96660 10432 96724 10436
rect 96660 10376 96674 10432
rect 96674 10376 96724 10432
rect 96660 10372 96724 10376
rect 125272 10372 125336 10436
rect 154252 10432 154316 10436
rect 154252 10376 154302 10432
rect 154302 10376 154316 10432
rect 154252 10372 154316 10376
rect 172928 10372 172992 10436
rect 181024 10372 181088 10436
rect 190592 10372 190656 10436
rect 192800 10432 192864 10436
rect 192800 10376 192850 10432
rect 192850 10376 192864 10432
rect 192800 10372 192864 10376
rect 202368 10432 202432 10436
rect 202368 10376 202418 10432
rect 202418 10376 202432 10432
rect 202368 10372 202432 10376
rect 210004 10372 210068 10436
rect 221044 10372 221108 10436
rect 245608 10372 245672 10436
rect 252968 10372 253032 10436
rect 261064 10372 261128 10436
rect 265480 10372 265544 10436
rect 31708 10236 31772 10300
rect 34928 10236 34992 10300
rect 35664 10296 35728 10300
rect 35664 10240 35678 10296
rect 35678 10240 35728 10296
rect 35664 10236 35728 10240
rect 36400 10236 36464 10300
rect 37136 10236 37200 10300
rect 37872 10236 37936 10300
rect 38608 10236 38672 10300
rect 39344 10236 39408 10300
rect 40080 10236 40144 10300
rect 40816 10296 40880 10300
rect 40816 10240 40830 10296
rect 40830 10240 40880 10296
rect 40816 10236 40880 10240
rect 41552 10236 41616 10300
rect 42288 10236 42352 10300
rect 43024 10236 43088 10300
rect 43760 10236 43824 10300
rect 44496 10236 44560 10300
rect 45232 10236 45296 10300
rect 45968 10296 46032 10300
rect 45968 10240 45982 10296
rect 45982 10240 46032 10296
rect 45968 10236 46032 10240
rect 46704 10236 46768 10300
rect 47440 10236 47504 10300
rect 48176 10296 48240 10300
rect 48176 10240 48226 10296
rect 48226 10240 48240 10296
rect 48176 10236 48240 10240
rect 48912 10236 48976 10300
rect 49648 10236 49712 10300
rect 50384 10236 50448 10300
rect 51120 10236 51184 10300
rect 51856 10236 51920 10300
rect 53328 10296 53392 10300
rect 53328 10240 53342 10296
rect 53342 10240 53392 10296
rect 53328 10236 53392 10240
rect 54064 10236 54128 10300
rect 54800 10296 54864 10300
rect 54800 10240 54850 10296
rect 54850 10240 54864 10296
rect 54800 10236 54864 10240
rect 55536 10236 55600 10300
rect 56272 10236 56336 10300
rect 57008 10236 57072 10300
rect 57744 10296 57808 10300
rect 57744 10240 57794 10296
rect 57794 10240 57808 10296
rect 57744 10236 57808 10240
rect 58480 10236 58544 10300
rect 59216 10296 59280 10300
rect 59216 10240 59266 10296
rect 59266 10240 59280 10296
rect 59216 10236 59280 10240
rect 59952 10236 60016 10300
rect 60688 10236 60752 10300
rect 61424 10236 61488 10300
rect 62160 10236 62224 10300
rect 62896 10236 62960 10300
rect 63632 10236 63696 10300
rect 64368 10236 64432 10300
rect 65104 10236 65168 10300
rect 65840 10296 65904 10300
rect 65840 10240 65890 10296
rect 65890 10240 65904 10296
rect 65840 10236 65904 10240
rect 66576 10236 66640 10300
rect 89668 10236 89732 10300
rect 103192 10296 103256 10300
rect 103192 10240 103242 10296
rect 103242 10240 103256 10296
rect 103192 10236 103256 10240
rect 103928 10296 103992 10300
rect 103928 10240 103942 10296
rect 103942 10240 103992 10296
rect 103928 10236 103992 10240
rect 104664 10296 104728 10300
rect 104664 10240 104714 10296
rect 104714 10240 104728 10296
rect 104664 10236 104728 10240
rect 105400 10236 105464 10300
rect 106136 10236 106200 10300
rect 106872 10236 106936 10300
rect 107608 10236 107672 10300
rect 108344 10296 108408 10300
rect 108344 10240 108394 10296
rect 108394 10240 108408 10296
rect 108344 10236 108408 10240
rect 109080 10296 109144 10300
rect 109080 10240 109094 10296
rect 109094 10240 109144 10296
rect 109080 10236 109144 10240
rect 109816 10236 109880 10300
rect 110552 10236 110616 10300
rect 111288 10236 111352 10300
rect 112024 10236 112088 10300
rect 112760 10236 112824 10300
rect 113496 10296 113560 10300
rect 113496 10240 113546 10296
rect 113546 10240 113560 10296
rect 113496 10236 113560 10240
rect 114232 10296 114296 10300
rect 114232 10240 114246 10296
rect 114246 10240 114296 10296
rect 114232 10236 114296 10240
rect 114968 10236 115032 10300
rect 115704 10296 115768 10300
rect 115704 10240 115754 10296
rect 115754 10240 115768 10296
rect 115704 10236 115768 10240
rect 116440 10236 116504 10300
rect 117176 10296 117240 10300
rect 117176 10240 117226 10296
rect 117226 10240 117240 10296
rect 117176 10236 117240 10240
rect 117912 10236 117976 10300
rect 118648 10296 118712 10300
rect 118648 10240 118698 10296
rect 118698 10240 118712 10296
rect 118648 10236 118712 10240
rect 119384 10296 119448 10300
rect 119384 10240 119398 10296
rect 119398 10240 119448 10296
rect 119384 10236 119448 10240
rect 120120 10236 120184 10300
rect 120856 10236 120920 10300
rect 121592 10236 121656 10300
rect 122328 10296 122392 10300
rect 122328 10240 122378 10296
rect 122378 10240 122392 10296
rect 122328 10236 122392 10240
rect 123064 10236 123128 10300
rect 123800 10236 123864 10300
rect 124536 10236 124600 10300
rect 126008 10236 126072 10300
rect 126744 10236 126808 10300
rect 127480 10236 127544 10300
rect 128216 10296 128280 10300
rect 128216 10240 128266 10296
rect 128266 10240 128280 10296
rect 128216 10236 128280 10240
rect 128952 10236 129016 10300
rect 129688 10296 129752 10300
rect 129688 10240 129702 10296
rect 129702 10240 129752 10296
rect 129688 10236 129752 10240
rect 130424 10236 130488 10300
rect 131160 10236 131224 10300
rect 131896 10236 131960 10300
rect 132632 10236 132696 10300
rect 133368 10296 133432 10300
rect 133368 10240 133418 10296
rect 133418 10240 133432 10296
rect 133368 10236 133432 10240
rect 134104 10296 134168 10300
rect 134104 10240 134154 10296
rect 134154 10240 134168 10296
rect 134104 10236 134168 10240
rect 134840 10236 134904 10300
rect 138060 10236 138124 10300
rect 142476 10236 142540 10300
rect 148364 10236 148428 10300
rect 171456 10236 171520 10300
rect 173664 10236 173728 10300
rect 174400 10296 174464 10300
rect 174400 10240 174450 10296
rect 174450 10240 174464 10296
rect 174400 10236 174464 10240
rect 175136 10296 175200 10300
rect 175136 10240 175186 10296
rect 175186 10240 175200 10296
rect 175136 10236 175200 10240
rect 175872 10296 175936 10300
rect 175872 10240 175922 10296
rect 175922 10240 175936 10296
rect 175872 10236 175936 10240
rect 176608 10236 176672 10300
rect 177344 10236 177408 10300
rect 178080 10236 178144 10300
rect 178816 10236 178880 10300
rect 180288 10236 180352 10300
rect 181760 10236 181824 10300
rect 182496 10296 182560 10300
rect 182496 10240 182546 10296
rect 182546 10240 182560 10296
rect 182496 10236 182560 10240
rect 183232 10296 183296 10300
rect 183232 10240 183282 10296
rect 183282 10240 183296 10296
rect 183232 10236 183296 10240
rect 183968 10236 184032 10300
rect 184704 10296 184768 10300
rect 184704 10240 184754 10296
rect 184754 10240 184768 10296
rect 184704 10236 184768 10240
rect 185440 10296 185504 10300
rect 185440 10240 185490 10296
rect 185490 10240 185504 10296
rect 185440 10236 185504 10240
rect 186176 10296 186240 10300
rect 186176 10240 186226 10296
rect 186226 10240 186240 10296
rect 186176 10236 186240 10240
rect 186912 10296 186976 10300
rect 186912 10240 186962 10296
rect 186962 10240 186976 10296
rect 186912 10236 186976 10240
rect 187648 10296 187712 10300
rect 187648 10240 187698 10296
rect 187698 10240 187712 10296
rect 187648 10236 187712 10240
rect 188384 10236 188448 10300
rect 189120 10236 189184 10300
rect 189856 10296 189920 10300
rect 189856 10240 189906 10296
rect 189906 10240 189920 10296
rect 189856 10236 189920 10240
rect 191328 10296 191392 10300
rect 191328 10240 191378 10296
rect 191378 10240 191392 10296
rect 191328 10236 191392 10240
rect 192064 10236 192128 10300
rect 193536 10236 193600 10300
rect 194272 10296 194336 10300
rect 194272 10240 194322 10296
rect 194322 10240 194336 10296
rect 194272 10236 194336 10240
rect 195008 10236 195072 10300
rect 195744 10296 195808 10300
rect 195744 10240 195794 10296
rect 195794 10240 195808 10296
rect 195744 10236 195808 10240
rect 196480 10296 196544 10300
rect 196480 10240 196530 10296
rect 196530 10240 196544 10296
rect 196480 10236 196544 10240
rect 197216 10296 197280 10300
rect 197216 10240 197266 10296
rect 197266 10240 197280 10296
rect 197216 10236 197280 10240
rect 197952 10296 198016 10300
rect 197952 10240 198002 10296
rect 198002 10240 198016 10296
rect 197952 10236 198016 10240
rect 198688 10236 198752 10300
rect 199424 10236 199488 10300
rect 200160 10236 200224 10300
rect 200896 10296 200960 10300
rect 200896 10240 200946 10296
rect 200946 10240 200960 10296
rect 200896 10236 200960 10240
rect 201632 10236 201696 10300
rect 203104 10236 203168 10300
rect 205588 10236 205652 10300
rect 220308 10296 220372 10300
rect 220308 10240 220358 10296
rect 220358 10240 220372 10296
rect 220308 10236 220372 10240
rect 239720 10236 239784 10300
rect 240456 10236 240520 10300
rect 241192 10296 241256 10300
rect 241192 10240 241242 10296
rect 241242 10240 241256 10296
rect 241192 10236 241256 10240
rect 241928 10236 241992 10300
rect 242664 10236 242728 10300
rect 243400 10296 243464 10300
rect 243400 10240 243450 10296
rect 243450 10240 243464 10296
rect 243400 10236 243464 10240
rect 244136 10296 244200 10300
rect 244136 10240 244186 10296
rect 244186 10240 244200 10296
rect 244136 10236 244200 10240
rect 244872 10236 244936 10300
rect 246344 10296 246408 10300
rect 246344 10240 246394 10296
rect 246394 10240 246408 10296
rect 246344 10236 246408 10240
rect 247080 10296 247144 10300
rect 247080 10240 247130 10296
rect 247130 10240 247144 10296
rect 247080 10236 247144 10240
rect 247816 10236 247880 10300
rect 248552 10236 248616 10300
rect 249288 10296 249352 10300
rect 249288 10240 249338 10296
rect 249338 10240 249352 10296
rect 249288 10236 249352 10240
rect 250024 10236 250088 10300
rect 250760 10236 250824 10300
rect 251496 10296 251560 10300
rect 251496 10240 251546 10296
rect 251546 10240 251560 10296
rect 251496 10236 251560 10240
rect 252232 10296 252296 10300
rect 252232 10240 252282 10296
rect 252282 10240 252296 10296
rect 252232 10236 252296 10240
rect 253704 10296 253768 10300
rect 253704 10240 253754 10296
rect 253754 10240 253768 10296
rect 253704 10236 253768 10240
rect 254440 10236 254504 10300
rect 255176 10236 255240 10300
rect 255912 10236 255976 10300
rect 256648 10296 256712 10300
rect 256648 10240 256698 10296
rect 256698 10240 256712 10296
rect 256648 10236 256712 10240
rect 257384 10236 257448 10300
rect 258120 10236 258184 10300
rect 258856 10236 258920 10300
rect 259592 10236 259656 10300
rect 260328 10236 260392 10300
rect 261800 10296 261864 10300
rect 261800 10240 261850 10296
rect 261850 10240 261864 10296
rect 261800 10236 261864 10240
rect 262536 10296 262600 10300
rect 262536 10240 262550 10296
rect 262550 10240 262600 10296
rect 262536 10236 262600 10240
rect 263272 10296 263336 10300
rect 263272 10240 263322 10296
rect 263322 10240 263336 10296
rect 263272 10236 263336 10240
rect 264008 10236 264072 10300
rect 266216 10296 266280 10300
rect 266216 10240 266230 10296
rect 266230 10240 266280 10296
rect 266216 10236 266280 10240
rect 1532 10100 1596 10164
rect 2268 10100 2332 10164
rect 3740 10100 3804 10164
rect 4476 10100 4540 10164
rect 5212 10100 5276 10164
rect 5948 10100 6012 10164
rect 6684 10100 6748 10164
rect 7420 10100 7484 10164
rect 8892 10100 8956 10164
rect 9628 10160 9692 10164
rect 9628 10104 9642 10160
rect 9642 10104 9692 10160
rect 9628 10100 9692 10104
rect 10364 10100 10428 10164
rect 11100 10100 11164 10164
rect 11836 10100 11900 10164
rect 12572 10100 12636 10164
rect 14044 10100 14108 10164
rect 14780 10100 14844 10164
rect 15516 10100 15580 10164
rect 16252 10100 16316 10164
rect 16988 10100 17052 10164
rect 17724 10100 17788 10164
rect 18460 10100 18524 10164
rect 71268 10100 71332 10164
rect 79364 10100 79428 10164
rect 83044 10160 83108 10164
rect 83044 10104 83094 10160
rect 83094 10104 83108 10160
rect 83044 10100 83108 10104
rect 83780 10100 83844 10164
rect 84516 10100 84580 10164
rect 85252 10100 85316 10164
rect 138796 10100 138860 10164
rect 140268 10100 140332 10164
rect 141004 10100 141068 10164
rect 141740 10100 141804 10164
rect 143212 10100 143276 10164
rect 143948 10100 144012 10164
rect 145420 10100 145484 10164
rect 146156 10100 146220 10164
rect 146892 10100 146956 10164
rect 149100 10100 149164 10164
rect 150572 10100 150636 10164
rect 151308 10100 151372 10164
rect 152044 10100 152108 10164
rect 152780 10160 152844 10164
rect 152780 10104 152830 10160
rect 152830 10104 152844 10160
rect 152780 10100 152844 10104
rect 153516 10100 153580 10164
rect 206324 10100 206388 10164
rect 207060 10100 207124 10164
rect 208532 10100 208596 10164
rect 209268 10160 209332 10164
rect 209268 10104 209318 10160
rect 209318 10104 209332 10160
rect 209268 10100 209332 10104
rect 210740 10100 210804 10164
rect 212212 10100 212276 10164
rect 213684 10100 213748 10164
rect 214420 10160 214484 10164
rect 214420 10104 214470 10160
rect 214470 10104 214484 10160
rect 214420 10100 214484 10104
rect 215892 10100 215956 10164
rect 217364 10100 217428 10164
rect 218836 10100 218900 10164
rect 219572 10100 219636 10164
rect 222516 10100 222580 10164
rect 223252 10100 223316 10164
rect 91140 9964 91204 10028
rect 3004 9828 3068 9892
rect 8156 9888 8220 9892
rect 8156 9832 8206 9888
rect 8206 9832 8220 9888
rect 8156 9828 8220 9832
rect 13308 9828 13372 9892
rect 19932 9828 19996 9892
rect 69796 9828 69860 9892
rect 77156 9888 77220 9892
rect 77156 9832 77206 9888
rect 77206 9832 77220 9888
rect 77156 9828 77220 9832
rect 78628 9888 78692 9892
rect 78628 9832 78678 9888
rect 78678 9832 78692 9888
rect 78628 9828 78692 9832
rect 80836 9828 80900 9892
rect 85988 9828 86052 9892
rect 139532 9828 139596 9892
rect 144684 9828 144748 9892
rect 149836 9828 149900 9892
rect 154988 9828 155052 9892
rect 211476 9828 211540 9892
rect 216628 9828 216692 9892
rect 221780 9828 221844 9892
rect 68548 9820 68612 9824
rect 68548 9764 68552 9820
rect 68552 9764 68608 9820
rect 68608 9764 68612 9820
rect 68548 9760 68612 9764
rect 68628 9820 68692 9824
rect 68628 9764 68632 9820
rect 68632 9764 68688 9820
rect 68688 9764 68692 9820
rect 68628 9760 68692 9764
rect 68708 9820 68772 9824
rect 68708 9764 68712 9820
rect 68712 9764 68768 9820
rect 68768 9764 68772 9820
rect 68708 9760 68772 9764
rect 68788 9820 68852 9824
rect 68788 9764 68792 9820
rect 68792 9764 68848 9820
rect 68848 9764 68852 9820
rect 68788 9760 68852 9764
rect 136145 9820 136209 9824
rect 136145 9764 136149 9820
rect 136149 9764 136205 9820
rect 136205 9764 136209 9820
rect 136145 9760 136209 9764
rect 136225 9820 136289 9824
rect 136225 9764 136229 9820
rect 136229 9764 136285 9820
rect 136285 9764 136289 9820
rect 136225 9760 136289 9764
rect 136305 9820 136369 9824
rect 136305 9764 136309 9820
rect 136309 9764 136365 9820
rect 136365 9764 136369 9820
rect 136305 9760 136369 9764
rect 136385 9820 136449 9824
rect 136385 9764 136389 9820
rect 136389 9764 136445 9820
rect 136445 9764 136449 9820
rect 136385 9760 136449 9764
rect 203742 9820 203806 9824
rect 203742 9764 203746 9820
rect 203746 9764 203802 9820
rect 203802 9764 203806 9820
rect 203742 9760 203806 9764
rect 203822 9820 203886 9824
rect 203822 9764 203826 9820
rect 203826 9764 203882 9820
rect 203882 9764 203886 9820
rect 203822 9760 203886 9764
rect 203902 9820 203966 9824
rect 203902 9764 203906 9820
rect 203906 9764 203962 9820
rect 203962 9764 203966 9820
rect 203902 9760 203966 9764
rect 203982 9820 204046 9824
rect 203982 9764 203986 9820
rect 203986 9764 204042 9820
rect 204042 9764 204046 9820
rect 203982 9760 204046 9764
rect 271339 9820 271403 9824
rect 271339 9764 271343 9820
rect 271343 9764 271399 9820
rect 271399 9764 271403 9820
rect 271339 9760 271403 9764
rect 271419 9820 271483 9824
rect 271419 9764 271423 9820
rect 271423 9764 271479 9820
rect 271479 9764 271483 9820
rect 271419 9760 271483 9764
rect 271499 9820 271563 9824
rect 271499 9764 271503 9820
rect 271503 9764 271559 9820
rect 271559 9764 271563 9820
rect 271499 9760 271563 9764
rect 271579 9820 271643 9824
rect 271579 9764 271583 9820
rect 271583 9764 271639 9820
rect 271639 9764 271643 9820
rect 271579 9760 271643 9764
rect 25820 9752 25884 9756
rect 25820 9696 25870 9752
rect 25870 9696 25884 9752
rect 25820 9692 25884 9696
rect 26556 9692 26620 9756
rect 29500 9692 29564 9756
rect 30236 9752 30300 9756
rect 30236 9696 30286 9752
rect 30286 9696 30300 9752
rect 30236 9692 30300 9696
rect 92612 9692 92676 9756
rect 93348 9692 93412 9756
rect 95556 9692 95620 9756
rect 96292 9752 96356 9756
rect 96292 9696 96342 9752
rect 96342 9696 96356 9752
rect 96292 9692 96356 9696
rect 98500 9692 98564 9756
rect 99972 9692 100036 9756
rect 167500 9692 167564 9756
rect 168972 9692 169036 9756
rect 69060 9616 69124 9620
rect 69060 9560 69110 9616
rect 69110 9560 69124 9616
rect 69060 9556 69124 9560
rect 70532 9556 70596 9620
rect 72740 9556 72804 9620
rect 74212 9616 74276 9620
rect 74212 9560 74262 9616
rect 74262 9560 74276 9616
rect 74212 9556 74276 9560
rect 75684 9556 75748 9620
rect 76420 9616 76484 9620
rect 76420 9560 76470 9616
rect 76470 9560 76484 9616
rect 76420 9556 76484 9560
rect 77892 9556 77956 9620
rect 80100 9556 80164 9620
rect 137324 9556 137388 9620
rect 215156 9556 215220 9620
rect 156460 9420 156524 9484
rect 223988 9480 224052 9484
rect 223988 9424 224038 9480
rect 224038 9424 224052 9480
rect 223988 9420 224052 9424
rect 227668 9420 227732 9484
rect 228404 9420 228468 9484
rect 229876 9480 229940 9484
rect 229876 9424 229890 9480
rect 229890 9424 229940 9480
rect 229876 9420 229940 9424
rect 232084 9420 232148 9484
rect 233556 9420 233620 9484
rect 235764 9420 235828 9484
rect 267596 9480 267660 9484
rect 267596 9424 267610 9480
rect 267610 9424 267660 9480
rect 267596 9420 267660 9424
rect 34750 9276 34814 9280
rect 34750 9220 34754 9276
rect 34754 9220 34810 9276
rect 34810 9220 34814 9276
rect 34750 9216 34814 9220
rect 34830 9276 34894 9280
rect 34830 9220 34834 9276
rect 34834 9220 34890 9276
rect 34890 9220 34894 9276
rect 34830 9216 34894 9220
rect 34910 9276 34974 9280
rect 34910 9220 34914 9276
rect 34914 9220 34970 9276
rect 34970 9220 34974 9276
rect 34910 9216 34974 9220
rect 34990 9276 35054 9280
rect 34990 9220 34994 9276
rect 34994 9220 35050 9276
rect 35050 9220 35054 9276
rect 34990 9216 35054 9220
rect 102347 9276 102411 9280
rect 102347 9220 102351 9276
rect 102351 9220 102407 9276
rect 102407 9220 102411 9276
rect 102347 9216 102411 9220
rect 102427 9276 102491 9280
rect 102427 9220 102431 9276
rect 102431 9220 102487 9276
rect 102487 9220 102491 9276
rect 102427 9216 102491 9220
rect 102507 9276 102571 9280
rect 102507 9220 102511 9276
rect 102511 9220 102567 9276
rect 102567 9220 102571 9276
rect 102507 9216 102571 9220
rect 102587 9276 102651 9280
rect 102587 9220 102591 9276
rect 102591 9220 102647 9276
rect 102647 9220 102651 9276
rect 102587 9216 102651 9220
rect 169944 9276 170008 9280
rect 169944 9220 169948 9276
rect 169948 9220 170004 9276
rect 170004 9220 170008 9276
rect 169944 9216 170008 9220
rect 170024 9276 170088 9280
rect 170024 9220 170028 9276
rect 170028 9220 170084 9276
rect 170084 9220 170088 9276
rect 170024 9216 170088 9220
rect 170104 9276 170168 9280
rect 170104 9220 170108 9276
rect 170108 9220 170164 9276
rect 170164 9220 170168 9276
rect 170104 9216 170168 9220
rect 170184 9276 170248 9280
rect 170184 9220 170188 9276
rect 170188 9220 170244 9276
rect 170244 9220 170248 9276
rect 170184 9216 170248 9220
rect 237541 9276 237605 9280
rect 237541 9220 237545 9276
rect 237545 9220 237601 9276
rect 237601 9220 237605 9276
rect 237541 9216 237605 9220
rect 237621 9276 237685 9280
rect 237621 9220 237625 9276
rect 237625 9220 237681 9276
rect 237681 9220 237685 9276
rect 237621 9216 237685 9220
rect 237701 9276 237765 9280
rect 237701 9220 237705 9276
rect 237705 9220 237761 9276
rect 237761 9220 237765 9276
rect 237701 9216 237765 9220
rect 237781 9276 237845 9280
rect 237781 9220 237785 9276
rect 237785 9220 237841 9276
rect 237841 9220 237845 9276
rect 237781 9216 237845 9220
rect 796 9148 860 9212
rect 24348 9148 24412 9212
rect 32444 9148 32508 9212
rect 88196 9208 88260 9212
rect 88196 9152 88246 9208
rect 88246 9152 88260 9208
rect 88196 9148 88260 9152
rect 91876 9148 91940 9212
rect 100708 9148 100772 9212
rect 168236 9148 168300 9212
rect 236500 9148 236564 9212
rect 73476 9072 73540 9076
rect 73476 9016 73490 9072
rect 73490 9016 73540 9072
rect 73476 9012 73540 9016
rect 74948 9012 75012 9076
rect 213868 9012 213932 9076
rect 22140 8936 22204 8940
rect 22140 8880 22154 8936
rect 22154 8880 22204 8936
rect 22140 8876 22204 8880
rect 96292 8876 96356 8940
rect 68548 8732 68612 8736
rect 68548 8676 68552 8732
rect 68552 8676 68608 8732
rect 68608 8676 68612 8732
rect 68548 8672 68612 8676
rect 68628 8732 68692 8736
rect 68628 8676 68632 8732
rect 68632 8676 68688 8732
rect 68688 8676 68692 8732
rect 68628 8672 68692 8676
rect 68708 8732 68772 8736
rect 68708 8676 68712 8732
rect 68712 8676 68768 8732
rect 68768 8676 68772 8732
rect 68708 8672 68772 8676
rect 68788 8732 68852 8736
rect 68788 8676 68792 8732
rect 68792 8676 68848 8732
rect 68848 8676 68852 8732
rect 68788 8672 68852 8676
rect 136145 8732 136209 8736
rect 136145 8676 136149 8732
rect 136149 8676 136205 8732
rect 136205 8676 136209 8732
rect 136145 8672 136209 8676
rect 136225 8732 136289 8736
rect 136225 8676 136229 8732
rect 136229 8676 136285 8732
rect 136285 8676 136289 8732
rect 136225 8672 136289 8676
rect 136305 8732 136369 8736
rect 136305 8676 136309 8732
rect 136309 8676 136365 8732
rect 136365 8676 136369 8732
rect 136305 8672 136369 8676
rect 136385 8732 136449 8736
rect 136385 8676 136389 8732
rect 136389 8676 136445 8732
rect 136445 8676 136449 8732
rect 136385 8672 136449 8676
rect 203742 8732 203806 8736
rect 203742 8676 203746 8732
rect 203746 8676 203802 8732
rect 203802 8676 203806 8732
rect 203742 8672 203806 8676
rect 203822 8732 203886 8736
rect 203822 8676 203826 8732
rect 203826 8676 203882 8732
rect 203882 8676 203886 8732
rect 203822 8672 203886 8676
rect 203902 8732 203966 8736
rect 203902 8676 203906 8732
rect 203906 8676 203962 8732
rect 203962 8676 203966 8732
rect 203902 8672 203966 8676
rect 203982 8732 204046 8736
rect 203982 8676 203986 8732
rect 203986 8676 204042 8732
rect 204042 8676 204046 8732
rect 203982 8672 204046 8676
rect 21404 8664 21468 8668
rect 21404 8608 21418 8664
rect 21418 8608 21468 8664
rect 21404 8604 21468 8608
rect 27292 8604 27356 8668
rect 28028 8604 28092 8668
rect 28764 8604 28828 8668
rect 30972 8664 31036 8668
rect 30972 8608 31022 8664
rect 31022 8608 31036 8664
rect 30972 8604 31036 8608
rect 87460 8664 87524 8668
rect 87460 8608 87510 8664
rect 87510 8608 87524 8664
rect 87460 8604 87524 8608
rect 90404 8604 90468 8668
rect 94084 8604 94148 8668
rect 94820 8604 94884 8668
rect 97028 8604 97092 8668
rect 97764 8604 97828 8668
rect 99236 8604 99300 8668
rect 155724 8604 155788 8668
rect 227484 8876 227548 8940
rect 226012 8740 226076 8804
rect 271339 8732 271403 8736
rect 271339 8676 271343 8732
rect 271343 8676 271399 8732
rect 271399 8676 271403 8732
rect 271339 8672 271403 8676
rect 271419 8732 271483 8736
rect 271419 8676 271423 8732
rect 271423 8676 271479 8732
rect 271479 8676 271483 8732
rect 271419 8672 271483 8676
rect 271499 8732 271563 8736
rect 271499 8676 271503 8732
rect 271503 8676 271559 8732
rect 271559 8676 271563 8732
rect 271499 8672 271563 8676
rect 271579 8732 271643 8736
rect 271579 8676 271583 8732
rect 271583 8676 271639 8732
rect 271639 8676 271643 8732
rect 271579 8672 271643 8676
rect 224724 8664 224788 8668
rect 224724 8608 224738 8664
rect 224738 8608 224788 8664
rect 20668 8332 20732 8396
rect 22876 8392 22940 8396
rect 22876 8336 22926 8392
rect 22926 8336 22940 8392
rect 22876 8332 22940 8336
rect 23612 8392 23676 8396
rect 23612 8336 23662 8392
rect 23662 8336 23676 8392
rect 23612 8332 23676 8336
rect 25084 8332 25148 8396
rect 157196 8392 157260 8396
rect 157196 8336 157246 8392
rect 157246 8336 157260 8392
rect 157196 8332 157260 8336
rect 158668 8332 158732 8396
rect 160140 8332 160204 8396
rect 161612 8332 161676 8396
rect 163084 8332 163148 8396
rect 164556 8332 164620 8396
rect 166028 8332 166092 8396
rect 166764 8332 166828 8396
rect 34750 8188 34814 8192
rect 34750 8132 34754 8188
rect 34754 8132 34810 8188
rect 34810 8132 34814 8188
rect 34750 8128 34814 8132
rect 34830 8188 34894 8192
rect 34830 8132 34834 8188
rect 34834 8132 34890 8188
rect 34890 8132 34894 8188
rect 34830 8128 34894 8132
rect 34910 8188 34974 8192
rect 34910 8132 34914 8188
rect 34914 8132 34970 8188
rect 34970 8132 34974 8188
rect 34910 8128 34974 8132
rect 34990 8188 35054 8192
rect 34990 8132 34994 8188
rect 34994 8132 35050 8188
rect 35050 8132 35054 8188
rect 34990 8128 35054 8132
rect 102347 8188 102411 8192
rect 102347 8132 102351 8188
rect 102351 8132 102407 8188
rect 102407 8132 102411 8188
rect 102347 8128 102411 8132
rect 102427 8188 102491 8192
rect 102427 8132 102431 8188
rect 102431 8132 102487 8188
rect 102487 8132 102491 8188
rect 102427 8128 102491 8132
rect 102507 8188 102571 8192
rect 102507 8132 102511 8188
rect 102511 8132 102567 8188
rect 102567 8132 102571 8188
rect 102507 8128 102571 8132
rect 102587 8188 102651 8192
rect 102587 8132 102591 8188
rect 102591 8132 102647 8188
rect 102647 8132 102651 8188
rect 102587 8128 102651 8132
rect 169944 8188 170008 8192
rect 169944 8132 169948 8188
rect 169948 8132 170004 8188
rect 170004 8132 170008 8188
rect 169944 8128 170008 8132
rect 170024 8188 170088 8192
rect 170024 8132 170028 8188
rect 170028 8132 170084 8188
rect 170084 8132 170088 8188
rect 170024 8128 170088 8132
rect 170104 8188 170168 8192
rect 170104 8132 170108 8188
rect 170108 8132 170164 8188
rect 170164 8132 170168 8188
rect 170104 8128 170168 8132
rect 170184 8188 170248 8192
rect 170184 8132 170188 8188
rect 170188 8132 170244 8188
rect 170244 8132 170248 8188
rect 170184 8128 170248 8132
rect 224724 8604 224788 8608
rect 225460 8664 225524 8668
rect 225460 8608 225510 8664
rect 225510 8608 225524 8664
rect 225460 8604 225524 8608
rect 226196 8664 226260 8668
rect 226196 8608 226246 8664
rect 226246 8608 226260 8664
rect 226196 8604 226260 8608
rect 226932 8664 226996 8668
rect 226932 8608 226982 8664
rect 226982 8608 226996 8664
rect 226932 8604 226996 8608
rect 229140 8664 229204 8668
rect 229140 8608 229190 8664
rect 229190 8608 229204 8664
rect 229140 8604 229204 8608
rect 230612 8604 230676 8668
rect 231348 8604 231412 8668
rect 232820 8604 232884 8668
rect 234292 8604 234356 8668
rect 237236 8604 237300 8668
rect 227300 8468 227364 8532
rect 224356 8392 224420 8396
rect 224356 8336 224370 8392
rect 224370 8336 224420 8392
rect 224356 8332 224420 8336
rect 235028 8332 235092 8396
rect 237541 8188 237605 8192
rect 237541 8132 237545 8188
rect 237545 8132 237601 8188
rect 237601 8132 237605 8188
rect 237541 8128 237605 8132
rect 237621 8188 237685 8192
rect 237621 8132 237625 8188
rect 237625 8132 237681 8188
rect 237681 8132 237685 8188
rect 237621 8128 237685 8132
rect 237701 8188 237765 8192
rect 237701 8132 237705 8188
rect 237705 8132 237761 8188
rect 237761 8132 237765 8188
rect 237701 8128 237765 8132
rect 237781 8188 237845 8192
rect 237781 8132 237785 8188
rect 237785 8132 237841 8188
rect 237841 8132 237845 8188
rect 237781 8128 237845 8132
rect 88932 8060 88996 8124
rect 96844 8060 96908 8124
rect 157932 8060 157996 8124
rect 159404 8120 159468 8124
rect 159404 8064 159454 8120
rect 159454 8064 159468 8120
rect 159404 8060 159468 8064
rect 160876 8060 160940 8124
rect 163820 8060 163884 8124
rect 165292 8120 165356 8124
rect 165292 8064 165342 8120
rect 165342 8064 165356 8120
rect 165292 8060 165356 8064
rect 162348 7848 162412 7852
rect 162348 7792 162398 7848
rect 162398 7792 162412 7848
rect 162348 7788 162412 7792
rect 264836 8120 264900 8124
rect 264836 8064 264886 8120
rect 264886 8064 264900 8120
rect 264836 8060 264900 8064
rect 68548 7644 68612 7648
rect 68548 7588 68552 7644
rect 68552 7588 68608 7644
rect 68608 7588 68612 7644
rect 68548 7584 68612 7588
rect 68628 7644 68692 7648
rect 68628 7588 68632 7644
rect 68632 7588 68688 7644
rect 68688 7588 68692 7644
rect 68628 7584 68692 7588
rect 68708 7644 68772 7648
rect 68708 7588 68712 7644
rect 68712 7588 68768 7644
rect 68768 7588 68772 7644
rect 68708 7584 68772 7588
rect 68788 7644 68852 7648
rect 68788 7588 68792 7644
rect 68792 7588 68848 7644
rect 68848 7588 68852 7644
rect 68788 7584 68852 7588
rect 136145 7644 136209 7648
rect 136145 7588 136149 7644
rect 136149 7588 136205 7644
rect 136205 7588 136209 7644
rect 136145 7584 136209 7588
rect 136225 7644 136289 7648
rect 136225 7588 136229 7644
rect 136229 7588 136285 7644
rect 136285 7588 136289 7644
rect 136225 7584 136289 7588
rect 136305 7644 136369 7648
rect 136305 7588 136309 7644
rect 136309 7588 136365 7644
rect 136365 7588 136369 7644
rect 136305 7584 136369 7588
rect 136385 7644 136449 7648
rect 136385 7588 136389 7644
rect 136389 7588 136445 7644
rect 136445 7588 136449 7644
rect 136385 7584 136449 7588
rect 203742 7644 203806 7648
rect 203742 7588 203746 7644
rect 203746 7588 203802 7644
rect 203802 7588 203806 7644
rect 203742 7584 203806 7588
rect 203822 7644 203886 7648
rect 203822 7588 203826 7644
rect 203826 7588 203882 7644
rect 203882 7588 203886 7644
rect 203822 7584 203886 7588
rect 203902 7644 203966 7648
rect 203902 7588 203906 7644
rect 203906 7588 203962 7644
rect 203962 7588 203966 7644
rect 203902 7584 203966 7588
rect 203982 7644 204046 7648
rect 203982 7588 203986 7644
rect 203986 7588 204042 7644
rect 204042 7588 204046 7644
rect 203982 7584 204046 7588
rect 267780 7652 267844 7716
rect 219940 7516 220004 7580
rect 271339 7644 271403 7648
rect 271339 7588 271343 7644
rect 271343 7588 271399 7644
rect 271399 7588 271403 7644
rect 271339 7584 271403 7588
rect 271419 7644 271483 7648
rect 271419 7588 271423 7644
rect 271423 7588 271479 7644
rect 271479 7588 271483 7644
rect 271419 7584 271483 7588
rect 271499 7644 271563 7648
rect 271499 7588 271503 7644
rect 271503 7588 271559 7644
rect 271559 7588 271563 7644
rect 271499 7584 271563 7588
rect 271579 7644 271643 7648
rect 271579 7588 271583 7644
rect 271583 7588 271639 7644
rect 271639 7588 271643 7644
rect 271579 7584 271643 7588
rect 34750 7100 34814 7104
rect 34750 7044 34754 7100
rect 34754 7044 34810 7100
rect 34810 7044 34814 7100
rect 34750 7040 34814 7044
rect 34830 7100 34894 7104
rect 34830 7044 34834 7100
rect 34834 7044 34890 7100
rect 34890 7044 34894 7100
rect 34830 7040 34894 7044
rect 34910 7100 34974 7104
rect 34910 7044 34914 7100
rect 34914 7044 34970 7100
rect 34970 7044 34974 7100
rect 34910 7040 34974 7044
rect 34990 7100 35054 7104
rect 34990 7044 34994 7100
rect 34994 7044 35050 7100
rect 35050 7044 35054 7100
rect 34990 7040 35054 7044
rect 102347 7100 102411 7104
rect 102347 7044 102351 7100
rect 102351 7044 102407 7100
rect 102407 7044 102411 7100
rect 102347 7040 102411 7044
rect 102427 7100 102491 7104
rect 102427 7044 102431 7100
rect 102431 7044 102487 7100
rect 102487 7044 102491 7100
rect 102427 7040 102491 7044
rect 102507 7100 102571 7104
rect 102507 7044 102511 7100
rect 102511 7044 102567 7100
rect 102567 7044 102571 7100
rect 102507 7040 102571 7044
rect 102587 7100 102651 7104
rect 102587 7044 102591 7100
rect 102591 7044 102647 7100
rect 102647 7044 102651 7100
rect 102587 7040 102651 7044
rect 169944 7100 170008 7104
rect 169944 7044 169948 7100
rect 169948 7044 170004 7100
rect 170004 7044 170008 7100
rect 169944 7040 170008 7044
rect 170024 7100 170088 7104
rect 170024 7044 170028 7100
rect 170028 7044 170084 7100
rect 170084 7044 170088 7100
rect 170024 7040 170088 7044
rect 170104 7100 170168 7104
rect 170104 7044 170108 7100
rect 170108 7044 170164 7100
rect 170164 7044 170168 7100
rect 170104 7040 170168 7044
rect 170184 7100 170248 7104
rect 170184 7044 170188 7100
rect 170188 7044 170244 7100
rect 170244 7044 170248 7100
rect 170184 7040 170248 7044
rect 237541 7100 237605 7104
rect 237541 7044 237545 7100
rect 237545 7044 237601 7100
rect 237601 7044 237605 7100
rect 237541 7040 237605 7044
rect 237621 7100 237685 7104
rect 237621 7044 237625 7100
rect 237625 7044 237681 7100
rect 237681 7044 237685 7100
rect 237621 7040 237685 7044
rect 237701 7100 237765 7104
rect 237701 7044 237705 7100
rect 237705 7044 237761 7100
rect 237761 7044 237765 7100
rect 237701 7040 237765 7044
rect 237781 7100 237845 7104
rect 237781 7044 237785 7100
rect 237785 7044 237841 7100
rect 237841 7044 237845 7100
rect 237781 7040 237845 7044
rect 19196 6896 19260 6900
rect 19196 6840 19246 6896
rect 19246 6840 19260 6896
rect 19196 6836 19260 6840
rect 94268 6896 94332 6900
rect 94268 6840 94282 6896
rect 94282 6840 94332 6896
rect 94268 6836 94332 6840
rect 107148 6836 107212 6900
rect 220860 6700 220924 6764
rect 227484 6700 227548 6764
rect 266860 6836 266924 6900
rect 249012 6700 249076 6764
rect 151676 6564 151740 6628
rect 68548 6556 68612 6560
rect 68548 6500 68552 6556
rect 68552 6500 68608 6556
rect 68608 6500 68612 6556
rect 68548 6496 68612 6500
rect 68628 6556 68692 6560
rect 68628 6500 68632 6556
rect 68632 6500 68688 6556
rect 68688 6500 68692 6556
rect 68628 6496 68692 6500
rect 68708 6556 68772 6560
rect 68708 6500 68712 6556
rect 68712 6500 68768 6556
rect 68768 6500 68772 6556
rect 68708 6496 68772 6500
rect 68788 6556 68852 6560
rect 68788 6500 68792 6556
rect 68792 6500 68848 6556
rect 68848 6500 68852 6556
rect 68788 6496 68852 6500
rect 136145 6556 136209 6560
rect 136145 6500 136149 6556
rect 136149 6500 136205 6556
rect 136205 6500 136209 6556
rect 136145 6496 136209 6500
rect 136225 6556 136289 6560
rect 136225 6500 136229 6556
rect 136229 6500 136285 6556
rect 136285 6500 136289 6556
rect 136225 6496 136289 6500
rect 136305 6556 136369 6560
rect 136305 6500 136309 6556
rect 136309 6500 136365 6556
rect 136365 6500 136369 6556
rect 136305 6496 136369 6500
rect 136385 6556 136449 6560
rect 136385 6500 136389 6556
rect 136389 6500 136445 6556
rect 136445 6500 136449 6556
rect 136385 6496 136449 6500
rect 203742 6556 203806 6560
rect 203742 6500 203746 6556
rect 203746 6500 203802 6556
rect 203802 6500 203806 6556
rect 203742 6496 203806 6500
rect 203822 6556 203886 6560
rect 203822 6500 203826 6556
rect 203826 6500 203882 6556
rect 203882 6500 203886 6556
rect 203822 6496 203886 6500
rect 203902 6556 203966 6560
rect 203902 6500 203906 6556
rect 203906 6500 203962 6556
rect 203962 6500 203966 6556
rect 203902 6496 203966 6500
rect 203982 6556 204046 6560
rect 203982 6500 203986 6556
rect 203986 6500 204042 6556
rect 204042 6500 204046 6556
rect 203982 6496 204046 6500
rect 271339 6556 271403 6560
rect 271339 6500 271343 6556
rect 271343 6500 271399 6556
rect 271399 6500 271403 6556
rect 271339 6496 271403 6500
rect 271419 6556 271483 6560
rect 271419 6500 271423 6556
rect 271423 6500 271479 6556
rect 271479 6500 271483 6556
rect 271419 6496 271483 6500
rect 271499 6556 271563 6560
rect 271499 6500 271503 6556
rect 271503 6500 271559 6556
rect 271559 6500 271563 6556
rect 271499 6496 271563 6500
rect 271579 6556 271643 6560
rect 271579 6500 271583 6556
rect 271583 6500 271639 6556
rect 271639 6500 271643 6556
rect 271579 6496 271643 6500
rect 93900 6292 93964 6356
rect 268516 6156 268580 6220
rect 269988 6156 270052 6220
rect 271092 6292 271156 6356
rect 34750 6012 34814 6016
rect 34750 5956 34754 6012
rect 34754 5956 34810 6012
rect 34810 5956 34814 6012
rect 34750 5952 34814 5956
rect 34830 6012 34894 6016
rect 34830 5956 34834 6012
rect 34834 5956 34890 6012
rect 34890 5956 34894 6012
rect 34830 5952 34894 5956
rect 34910 6012 34974 6016
rect 34910 5956 34914 6012
rect 34914 5956 34970 6012
rect 34970 5956 34974 6012
rect 34910 5952 34974 5956
rect 34990 6012 35054 6016
rect 34990 5956 34994 6012
rect 34994 5956 35050 6012
rect 35050 5956 35054 6012
rect 34990 5952 35054 5956
rect 102347 6012 102411 6016
rect 102347 5956 102351 6012
rect 102351 5956 102407 6012
rect 102407 5956 102411 6012
rect 102347 5952 102411 5956
rect 102427 6012 102491 6016
rect 102427 5956 102431 6012
rect 102431 5956 102487 6012
rect 102487 5956 102491 6012
rect 102427 5952 102491 5956
rect 102507 6012 102571 6016
rect 102507 5956 102511 6012
rect 102511 5956 102567 6012
rect 102567 5956 102571 6012
rect 102507 5952 102571 5956
rect 102587 6012 102651 6016
rect 102587 5956 102591 6012
rect 102591 5956 102647 6012
rect 102647 5956 102651 6012
rect 102587 5952 102651 5956
rect 169944 6012 170008 6016
rect 169944 5956 169948 6012
rect 169948 5956 170004 6012
rect 170004 5956 170008 6012
rect 169944 5952 170008 5956
rect 170024 6012 170088 6016
rect 170024 5956 170028 6012
rect 170028 5956 170084 6012
rect 170084 5956 170088 6012
rect 170024 5952 170088 5956
rect 170104 6012 170168 6016
rect 170104 5956 170108 6012
rect 170108 5956 170164 6012
rect 170164 5956 170168 6012
rect 170104 5952 170168 5956
rect 170184 6012 170248 6016
rect 170184 5956 170188 6012
rect 170188 5956 170244 6012
rect 170244 5956 170248 6012
rect 170184 5952 170248 5956
rect 237541 6012 237605 6016
rect 237541 5956 237545 6012
rect 237545 5956 237601 6012
rect 237601 5956 237605 6012
rect 237541 5952 237605 5956
rect 237621 6012 237685 6016
rect 237621 5956 237625 6012
rect 237625 5956 237681 6012
rect 237681 5956 237685 6012
rect 237621 5952 237685 5956
rect 237701 6012 237765 6016
rect 237701 5956 237705 6012
rect 237705 5956 237761 6012
rect 237761 5956 237765 6012
rect 237701 5952 237765 5956
rect 237781 6012 237845 6016
rect 237781 5956 237785 6012
rect 237785 5956 237841 6012
rect 237841 5956 237845 6012
rect 237781 5952 237845 5956
rect 213868 5748 213932 5812
rect 95188 5476 95252 5540
rect 68548 5468 68612 5472
rect 68548 5412 68552 5468
rect 68552 5412 68608 5468
rect 68608 5412 68612 5468
rect 68548 5408 68612 5412
rect 68628 5468 68692 5472
rect 68628 5412 68632 5468
rect 68632 5412 68688 5468
rect 68688 5412 68692 5468
rect 68628 5408 68692 5412
rect 68708 5468 68772 5472
rect 68708 5412 68712 5468
rect 68712 5412 68768 5468
rect 68768 5412 68772 5468
rect 68708 5408 68772 5412
rect 68788 5468 68852 5472
rect 68788 5412 68792 5468
rect 68792 5412 68848 5468
rect 68848 5412 68852 5468
rect 68788 5408 68852 5412
rect 151860 5612 151924 5676
rect 266308 5808 266372 5812
rect 266308 5752 266358 5808
rect 266358 5752 266372 5808
rect 266308 5748 266372 5752
rect 269252 5612 269316 5676
rect 270540 5672 270604 5676
rect 270540 5616 270554 5672
rect 270554 5616 270604 5672
rect 270540 5612 270604 5616
rect 220860 5476 220924 5540
rect 136145 5468 136209 5472
rect 136145 5412 136149 5468
rect 136149 5412 136205 5468
rect 136205 5412 136209 5468
rect 136145 5408 136209 5412
rect 136225 5468 136289 5472
rect 136225 5412 136229 5468
rect 136229 5412 136285 5468
rect 136285 5412 136289 5468
rect 136225 5408 136289 5412
rect 136305 5468 136369 5472
rect 136305 5412 136309 5468
rect 136309 5412 136365 5468
rect 136365 5412 136369 5468
rect 136305 5408 136369 5412
rect 136385 5468 136449 5472
rect 136385 5412 136389 5468
rect 136389 5412 136445 5468
rect 136445 5412 136449 5468
rect 136385 5408 136449 5412
rect 203742 5468 203806 5472
rect 203742 5412 203746 5468
rect 203746 5412 203802 5468
rect 203802 5412 203806 5468
rect 203742 5408 203806 5412
rect 203822 5468 203886 5472
rect 203822 5412 203826 5468
rect 203826 5412 203882 5468
rect 203882 5412 203886 5468
rect 203822 5408 203886 5412
rect 203902 5468 203966 5472
rect 203902 5412 203906 5468
rect 203906 5412 203962 5468
rect 203962 5412 203966 5468
rect 203902 5408 203966 5412
rect 203982 5468 204046 5472
rect 203982 5412 203986 5468
rect 203986 5412 204042 5468
rect 204042 5412 204046 5468
rect 203982 5408 204046 5412
rect 271339 5468 271403 5472
rect 271339 5412 271343 5468
rect 271343 5412 271399 5468
rect 271399 5412 271403 5468
rect 271339 5408 271403 5412
rect 271419 5468 271483 5472
rect 271419 5412 271423 5468
rect 271423 5412 271479 5468
rect 271479 5412 271483 5468
rect 271419 5408 271483 5412
rect 271499 5468 271563 5472
rect 271499 5412 271503 5468
rect 271503 5412 271559 5468
rect 271559 5412 271563 5468
rect 271499 5408 271563 5412
rect 271579 5468 271643 5472
rect 271579 5412 271583 5468
rect 271583 5412 271639 5468
rect 271639 5412 271643 5468
rect 271579 5408 271643 5412
rect 113036 5340 113100 5404
rect 249012 5340 249076 5404
rect 219940 5204 220004 5268
rect 34750 4924 34814 4928
rect 34750 4868 34754 4924
rect 34754 4868 34810 4924
rect 34810 4868 34814 4924
rect 34750 4864 34814 4868
rect 34830 4924 34894 4928
rect 34830 4868 34834 4924
rect 34834 4868 34890 4924
rect 34890 4868 34894 4924
rect 34830 4864 34894 4868
rect 34910 4924 34974 4928
rect 34910 4868 34914 4924
rect 34914 4868 34970 4924
rect 34970 4868 34974 4924
rect 34910 4864 34974 4868
rect 34990 4924 35054 4928
rect 34990 4868 34994 4924
rect 34994 4868 35050 4924
rect 35050 4868 35054 4924
rect 34990 4864 35054 4868
rect 102347 4924 102411 4928
rect 102347 4868 102351 4924
rect 102351 4868 102407 4924
rect 102407 4868 102411 4924
rect 102347 4864 102411 4868
rect 102427 4924 102491 4928
rect 102427 4868 102431 4924
rect 102431 4868 102487 4924
rect 102487 4868 102491 4924
rect 102427 4864 102491 4868
rect 102507 4924 102571 4928
rect 102507 4868 102511 4924
rect 102511 4868 102567 4924
rect 102567 4868 102571 4924
rect 102507 4864 102571 4868
rect 102587 4924 102651 4928
rect 102587 4868 102591 4924
rect 102591 4868 102647 4924
rect 102647 4868 102651 4924
rect 102587 4864 102651 4868
rect 169944 4924 170008 4928
rect 169944 4868 169948 4924
rect 169948 4868 170004 4924
rect 170004 4868 170008 4924
rect 169944 4864 170008 4868
rect 170024 4924 170088 4928
rect 170024 4868 170028 4924
rect 170028 4868 170084 4924
rect 170084 4868 170088 4924
rect 170024 4864 170088 4868
rect 170104 4924 170168 4928
rect 170104 4868 170108 4924
rect 170108 4868 170164 4924
rect 170164 4868 170168 4924
rect 170104 4864 170168 4868
rect 170184 4924 170248 4928
rect 170184 4868 170188 4924
rect 170188 4868 170244 4924
rect 170244 4868 170248 4924
rect 170184 4864 170248 4868
rect 237541 4924 237605 4928
rect 237541 4868 237545 4924
rect 237545 4868 237601 4924
rect 237601 4868 237605 4924
rect 237541 4864 237605 4868
rect 237621 4924 237685 4928
rect 237621 4868 237625 4924
rect 237625 4868 237681 4924
rect 237681 4868 237685 4924
rect 237621 4864 237685 4868
rect 237701 4924 237765 4928
rect 237701 4868 237705 4924
rect 237705 4868 237761 4924
rect 237761 4868 237765 4924
rect 237701 4864 237765 4868
rect 237781 4924 237845 4928
rect 237781 4868 237785 4924
rect 237785 4868 237841 4924
rect 237841 4868 237845 4924
rect 237781 4864 237845 4868
rect 106044 4796 106108 4860
rect 110276 4796 110340 4860
rect 225092 4796 225156 4860
rect 226196 4524 226260 4588
rect 68548 4380 68612 4384
rect 68548 4324 68552 4380
rect 68552 4324 68608 4380
rect 68608 4324 68612 4380
rect 68548 4320 68612 4324
rect 68628 4380 68692 4384
rect 68628 4324 68632 4380
rect 68632 4324 68688 4380
rect 68688 4324 68692 4380
rect 68628 4320 68692 4324
rect 68708 4380 68772 4384
rect 68708 4324 68712 4380
rect 68712 4324 68768 4380
rect 68768 4324 68772 4380
rect 68708 4320 68772 4324
rect 68788 4380 68852 4384
rect 68788 4324 68792 4380
rect 68792 4324 68848 4380
rect 68848 4324 68852 4380
rect 68788 4320 68852 4324
rect 96476 4116 96540 4180
rect 136145 4380 136209 4384
rect 136145 4324 136149 4380
rect 136149 4324 136205 4380
rect 136205 4324 136209 4380
rect 136145 4320 136209 4324
rect 136225 4380 136289 4384
rect 136225 4324 136229 4380
rect 136229 4324 136285 4380
rect 136285 4324 136289 4380
rect 136225 4320 136289 4324
rect 136305 4380 136369 4384
rect 136305 4324 136309 4380
rect 136309 4324 136365 4380
rect 136365 4324 136369 4380
rect 136305 4320 136369 4324
rect 136385 4380 136449 4384
rect 136385 4324 136389 4380
rect 136389 4324 136445 4380
rect 136445 4324 136449 4380
rect 136385 4320 136449 4324
rect 203742 4380 203806 4384
rect 203742 4324 203746 4380
rect 203746 4324 203802 4380
rect 203802 4324 203806 4380
rect 203742 4320 203806 4324
rect 203822 4380 203886 4384
rect 203822 4324 203826 4380
rect 203826 4324 203882 4380
rect 203882 4324 203886 4380
rect 203822 4320 203886 4324
rect 203902 4380 203966 4384
rect 203902 4324 203906 4380
rect 203906 4324 203962 4380
rect 203962 4324 203966 4380
rect 203902 4320 203966 4324
rect 203982 4380 204046 4384
rect 203982 4324 203986 4380
rect 203986 4324 204042 4380
rect 204042 4324 204046 4380
rect 203982 4320 204046 4324
rect 271339 4380 271403 4384
rect 271339 4324 271343 4380
rect 271343 4324 271399 4380
rect 271399 4324 271403 4380
rect 271339 4320 271403 4324
rect 271419 4380 271483 4384
rect 271419 4324 271423 4380
rect 271423 4324 271479 4380
rect 271479 4324 271483 4380
rect 271419 4320 271483 4324
rect 271499 4380 271563 4384
rect 271499 4324 271503 4380
rect 271503 4324 271559 4380
rect 271559 4324 271563 4380
rect 271499 4320 271563 4324
rect 271579 4380 271643 4384
rect 271579 4324 271583 4380
rect 271583 4324 271639 4380
rect 271639 4324 271643 4380
rect 271579 4320 271643 4324
rect 103284 3980 103348 4044
rect 104572 4040 104636 4044
rect 104572 3984 104586 4040
rect 104586 3984 104636 4040
rect 104572 3980 104636 3984
rect 105492 3980 105556 4044
rect 106964 3980 107028 4044
rect 107700 3980 107764 4044
rect 108252 3980 108316 4044
rect 109172 4040 109236 4044
rect 109172 3984 109222 4040
rect 109222 3984 109236 4040
rect 109172 3980 109236 3984
rect 109908 3980 109972 4044
rect 110644 4040 110708 4044
rect 110644 3984 110694 4040
rect 110694 3984 110708 4040
rect 110644 3980 110708 3984
rect 111196 4040 111260 4044
rect 111196 3984 111246 4040
rect 111246 3984 111260 4040
rect 111196 3980 111260 3984
rect 112116 3980 112180 4044
rect 112852 3980 112916 4044
rect 113220 3980 113284 4044
rect 153148 3980 153212 4044
rect 215156 4040 215220 4044
rect 215156 3984 215206 4040
rect 215206 3984 215220 4040
rect 215156 3980 215220 3984
rect 223988 3980 224052 4044
rect 34750 3836 34814 3840
rect 34750 3780 34754 3836
rect 34754 3780 34810 3836
rect 34810 3780 34814 3836
rect 34750 3776 34814 3780
rect 34830 3836 34894 3840
rect 34830 3780 34834 3836
rect 34834 3780 34890 3836
rect 34890 3780 34894 3836
rect 34830 3776 34894 3780
rect 34910 3836 34974 3840
rect 34910 3780 34914 3836
rect 34914 3780 34970 3836
rect 34970 3780 34974 3836
rect 34910 3776 34974 3780
rect 34990 3836 35054 3840
rect 34990 3780 34994 3836
rect 34994 3780 35050 3836
rect 35050 3780 35054 3836
rect 34990 3776 35054 3780
rect 102347 3836 102411 3840
rect 102347 3780 102351 3836
rect 102351 3780 102407 3836
rect 102407 3780 102411 3836
rect 102347 3776 102411 3780
rect 102427 3836 102491 3840
rect 102427 3780 102431 3836
rect 102431 3780 102487 3836
rect 102487 3780 102491 3836
rect 102427 3776 102491 3780
rect 102507 3836 102571 3840
rect 102507 3780 102511 3836
rect 102511 3780 102567 3836
rect 102567 3780 102571 3836
rect 102507 3776 102571 3780
rect 102587 3836 102651 3840
rect 102587 3780 102591 3836
rect 102591 3780 102647 3836
rect 102647 3780 102651 3836
rect 102587 3776 102651 3780
rect 97764 3708 97828 3772
rect 104020 3844 104084 3908
rect 226012 3844 226076 3908
rect 169944 3836 170008 3840
rect 169944 3780 169948 3836
rect 169948 3780 170004 3836
rect 170004 3780 170008 3836
rect 169944 3776 170008 3780
rect 170024 3836 170088 3840
rect 170024 3780 170028 3836
rect 170028 3780 170084 3836
rect 170084 3780 170088 3836
rect 170024 3776 170088 3780
rect 170104 3836 170168 3840
rect 170104 3780 170108 3836
rect 170108 3780 170164 3836
rect 170164 3780 170168 3836
rect 170104 3776 170168 3780
rect 170184 3836 170248 3840
rect 170184 3780 170188 3836
rect 170188 3780 170244 3836
rect 170244 3780 170248 3836
rect 170184 3776 170248 3780
rect 237541 3836 237605 3840
rect 237541 3780 237545 3836
rect 237545 3780 237601 3836
rect 237601 3780 237605 3836
rect 237541 3776 237605 3780
rect 237621 3836 237685 3840
rect 237621 3780 237625 3836
rect 237625 3780 237681 3836
rect 237681 3780 237685 3836
rect 237621 3776 237685 3780
rect 237701 3836 237765 3840
rect 237701 3780 237705 3836
rect 237705 3780 237761 3836
rect 237761 3780 237765 3836
rect 237701 3776 237765 3780
rect 237781 3836 237845 3840
rect 237781 3780 237785 3836
rect 237785 3780 237841 3836
rect 237841 3780 237845 3836
rect 237781 3776 237845 3780
rect 107148 3708 107212 3772
rect 218836 3768 218900 3772
rect 218836 3712 218886 3768
rect 218886 3712 218900 3768
rect 218836 3708 218900 3712
rect 223252 3708 223316 3772
rect 227300 3708 227364 3772
rect 223988 3572 224052 3636
rect 154252 3360 154316 3364
rect 154252 3304 154302 3360
rect 154302 3304 154316 3360
rect 154252 3300 154316 3304
rect 68548 3292 68612 3296
rect 68548 3236 68552 3292
rect 68552 3236 68608 3292
rect 68608 3236 68612 3292
rect 68548 3232 68612 3236
rect 68628 3292 68692 3296
rect 68628 3236 68632 3292
rect 68632 3236 68688 3292
rect 68688 3236 68692 3292
rect 68628 3232 68692 3236
rect 68708 3292 68772 3296
rect 68708 3236 68712 3292
rect 68712 3236 68768 3292
rect 68768 3236 68772 3292
rect 68708 3232 68772 3236
rect 68788 3292 68852 3296
rect 68788 3236 68792 3292
rect 68792 3236 68848 3292
rect 68848 3236 68852 3292
rect 68788 3232 68852 3236
rect 136145 3292 136209 3296
rect 136145 3236 136149 3292
rect 136149 3236 136205 3292
rect 136205 3236 136209 3292
rect 136145 3232 136209 3236
rect 136225 3292 136289 3296
rect 136225 3236 136229 3292
rect 136229 3236 136285 3292
rect 136285 3236 136289 3292
rect 136225 3232 136289 3236
rect 136305 3292 136369 3296
rect 136305 3236 136309 3292
rect 136309 3236 136365 3292
rect 136365 3236 136369 3292
rect 136305 3232 136369 3236
rect 136385 3292 136449 3296
rect 136385 3236 136389 3292
rect 136389 3236 136445 3292
rect 136445 3236 136449 3292
rect 136385 3232 136449 3236
rect 203742 3292 203806 3296
rect 203742 3236 203746 3292
rect 203746 3236 203802 3292
rect 203802 3236 203806 3292
rect 203742 3232 203806 3236
rect 203822 3292 203886 3296
rect 203822 3236 203826 3292
rect 203826 3236 203882 3292
rect 203882 3236 203886 3292
rect 203822 3232 203886 3236
rect 203902 3292 203966 3296
rect 203902 3236 203906 3292
rect 203906 3236 203962 3292
rect 203962 3236 203966 3292
rect 203902 3232 203966 3236
rect 203982 3292 204046 3296
rect 203982 3236 203986 3292
rect 203986 3236 204042 3292
rect 204042 3236 204046 3292
rect 203982 3232 204046 3236
rect 93900 3164 93964 3228
rect 96292 3164 96356 3228
rect 96844 3164 96908 3228
rect 100708 3224 100772 3228
rect 100708 3168 100758 3224
rect 100758 3168 100772 3224
rect 100708 3164 100772 3168
rect 110276 3164 110340 3228
rect 144684 3224 144748 3228
rect 144684 3168 144734 3224
rect 144734 3168 144748 3224
rect 144684 3164 144748 3168
rect 94084 3028 94148 3092
rect 211476 3088 211540 3092
rect 211476 3032 211526 3088
rect 211526 3032 211540 3088
rect 211476 3028 211540 3032
rect 217364 3164 217428 3228
rect 221044 3164 221108 3228
rect 271339 3292 271403 3296
rect 271339 3236 271343 3292
rect 271343 3236 271399 3292
rect 271399 3236 271403 3292
rect 271339 3232 271403 3236
rect 271419 3292 271483 3296
rect 271419 3236 271423 3292
rect 271423 3236 271479 3292
rect 271479 3236 271483 3292
rect 271419 3232 271483 3236
rect 271499 3292 271563 3296
rect 271499 3236 271503 3292
rect 271503 3236 271559 3292
rect 271559 3236 271563 3292
rect 271499 3232 271563 3236
rect 271579 3292 271643 3296
rect 271579 3236 271583 3292
rect 271583 3236 271639 3292
rect 271639 3236 271643 3292
rect 271579 3232 271643 3236
rect 258948 3224 259012 3228
rect 258948 3168 258998 3224
rect 258998 3168 259012 3224
rect 258948 3164 259012 3168
rect 796 2816 860 2820
rect 796 2760 846 2816
rect 846 2760 860 2816
rect 796 2756 860 2760
rect 19196 2816 19260 2820
rect 19196 2760 19246 2816
rect 19246 2760 19260 2816
rect 19196 2756 19260 2760
rect 22876 2816 22940 2820
rect 22876 2760 22890 2816
rect 22890 2760 22940 2816
rect 22876 2756 22940 2760
rect 25084 2816 25148 2820
rect 25084 2760 25098 2816
rect 25098 2760 25148 2816
rect 25084 2756 25148 2760
rect 27292 2756 27356 2820
rect 54892 2756 54956 2820
rect 95556 2756 95620 2820
rect 97028 2816 97092 2820
rect 97028 2760 97042 2816
rect 97042 2760 97092 2816
rect 97028 2756 97092 2760
rect 116532 2756 116596 2820
rect 123892 2756 123956 2820
rect 133460 2756 133524 2820
rect 145420 2816 145484 2820
rect 145420 2760 145470 2816
rect 145470 2760 145484 2816
rect 145420 2756 145484 2760
rect 149100 2892 149164 2956
rect 153516 2892 153580 2956
rect 154988 2952 155052 2956
rect 154988 2896 155038 2952
rect 155038 2896 155052 2952
rect 154988 2892 155052 2896
rect 156460 2816 156524 2820
rect 156460 2760 156474 2816
rect 156474 2760 156524 2816
rect 156460 2756 156524 2760
rect 189948 2756 190012 2820
rect 191420 2756 191484 2820
rect 198044 2756 198108 2820
rect 199516 2756 199580 2820
rect 200988 2756 201052 2820
rect 210740 2756 210804 2820
rect 216628 2892 216692 2956
rect 224356 2756 224420 2820
rect 226196 2892 226260 2956
rect 250852 3028 250916 3092
rect 246436 2892 246500 2956
rect 256004 2892 256068 2956
rect 259684 2756 259748 2820
rect 260420 2816 260484 2820
rect 260420 2760 260470 2816
rect 260470 2760 260484 2816
rect 260420 2756 260484 2760
rect 261892 2756 261956 2820
rect 271092 2756 271156 2820
rect 34750 2748 34814 2752
rect 34750 2692 34754 2748
rect 34754 2692 34810 2748
rect 34810 2692 34814 2748
rect 34750 2688 34814 2692
rect 34830 2748 34894 2752
rect 34830 2692 34834 2748
rect 34834 2692 34890 2748
rect 34890 2692 34894 2748
rect 34830 2688 34894 2692
rect 34910 2748 34974 2752
rect 34910 2692 34914 2748
rect 34914 2692 34970 2748
rect 34970 2692 34974 2748
rect 34910 2688 34974 2692
rect 34990 2748 35054 2752
rect 34990 2692 34994 2748
rect 34994 2692 35050 2748
rect 35050 2692 35054 2748
rect 34990 2688 35054 2692
rect 102347 2748 102411 2752
rect 102347 2692 102351 2748
rect 102351 2692 102407 2748
rect 102407 2692 102411 2748
rect 102347 2688 102411 2692
rect 102427 2748 102491 2752
rect 102427 2692 102431 2748
rect 102431 2692 102487 2748
rect 102487 2692 102491 2748
rect 102427 2688 102491 2692
rect 102507 2748 102571 2752
rect 102507 2692 102511 2748
rect 102511 2692 102567 2748
rect 102567 2692 102571 2748
rect 102507 2688 102571 2692
rect 102587 2748 102651 2752
rect 102587 2692 102591 2748
rect 102591 2692 102647 2748
rect 102647 2692 102651 2748
rect 102587 2688 102651 2692
rect 169944 2748 170008 2752
rect 169944 2692 169948 2748
rect 169948 2692 170004 2748
rect 170004 2692 170008 2748
rect 169944 2688 170008 2692
rect 170024 2748 170088 2752
rect 170024 2692 170028 2748
rect 170028 2692 170084 2748
rect 170084 2692 170088 2748
rect 170024 2688 170088 2692
rect 170104 2748 170168 2752
rect 170104 2692 170108 2748
rect 170108 2692 170164 2748
rect 170164 2692 170168 2748
rect 170104 2688 170168 2692
rect 170184 2748 170248 2752
rect 170184 2692 170188 2748
rect 170188 2692 170244 2748
rect 170244 2692 170248 2748
rect 170184 2688 170248 2692
rect 237541 2748 237605 2752
rect 237541 2692 237545 2748
rect 237545 2692 237601 2748
rect 237601 2692 237605 2748
rect 237541 2688 237605 2692
rect 237621 2748 237685 2752
rect 237621 2692 237625 2748
rect 237625 2692 237681 2748
rect 237681 2692 237685 2748
rect 237621 2688 237685 2692
rect 237701 2748 237765 2752
rect 237701 2692 237705 2748
rect 237705 2692 237761 2748
rect 237761 2692 237765 2748
rect 237701 2688 237765 2692
rect 237781 2748 237845 2752
rect 237781 2692 237785 2748
rect 237785 2692 237841 2748
rect 237841 2692 237845 2748
rect 237781 2688 237845 2692
rect 96660 2348 96724 2412
rect 151676 2408 151740 2412
rect 151676 2352 151726 2408
rect 151726 2352 151740 2408
rect 68548 2204 68612 2208
rect 68548 2148 68552 2204
rect 68552 2148 68608 2204
rect 68608 2148 68612 2204
rect 68548 2144 68612 2148
rect 68628 2204 68692 2208
rect 68628 2148 68632 2204
rect 68632 2148 68688 2204
rect 68688 2148 68692 2204
rect 68628 2144 68692 2148
rect 68708 2204 68772 2208
rect 68708 2148 68712 2204
rect 68712 2148 68768 2204
rect 68768 2148 68772 2204
rect 68708 2144 68772 2148
rect 68788 2204 68852 2208
rect 68788 2148 68792 2204
rect 68792 2148 68848 2204
rect 68848 2148 68852 2204
rect 68788 2144 68852 2148
rect 94268 2136 94332 2140
rect 94268 2080 94282 2136
rect 94282 2080 94332 2136
rect 94268 2076 94332 2080
rect 96476 2136 96540 2140
rect 96476 2080 96490 2136
rect 96490 2080 96540 2136
rect 96476 2076 96540 2080
rect 114324 2212 114388 2276
rect 151676 2348 151740 2352
rect 136145 2204 136209 2208
rect 136145 2148 136149 2204
rect 136149 2148 136205 2204
rect 136205 2148 136209 2204
rect 136145 2144 136209 2148
rect 136225 2204 136289 2208
rect 136225 2148 136229 2204
rect 136229 2148 136285 2204
rect 136285 2148 136289 2204
rect 136225 2144 136289 2148
rect 136305 2204 136369 2208
rect 136305 2148 136309 2204
rect 136309 2148 136365 2204
rect 136365 2148 136369 2204
rect 136305 2144 136369 2148
rect 136385 2204 136449 2208
rect 136385 2148 136389 2204
rect 136389 2148 136445 2204
rect 136445 2148 136449 2204
rect 136385 2144 136449 2148
rect 203742 2204 203806 2208
rect 203742 2148 203746 2204
rect 203746 2148 203802 2204
rect 203802 2148 203806 2204
rect 203742 2144 203806 2148
rect 203822 2204 203886 2208
rect 203822 2148 203826 2204
rect 203826 2148 203882 2204
rect 203882 2148 203886 2204
rect 203822 2144 203886 2148
rect 203902 2204 203966 2208
rect 203902 2148 203906 2204
rect 203906 2148 203962 2204
rect 203962 2148 203966 2204
rect 203902 2144 203966 2148
rect 203982 2204 204046 2208
rect 203982 2148 203986 2204
rect 203986 2148 204042 2204
rect 204042 2148 204046 2204
rect 203982 2144 204046 2148
rect 22140 1668 22204 1732
rect 271339 2204 271403 2208
rect 271339 2148 271343 2204
rect 271343 2148 271399 2204
rect 271399 2148 271403 2204
rect 271339 2144 271403 2148
rect 271419 2204 271483 2208
rect 271419 2148 271423 2204
rect 271423 2148 271479 2204
rect 271479 2148 271483 2204
rect 271419 2144 271483 2148
rect 271499 2204 271563 2208
rect 271499 2148 271503 2204
rect 271503 2148 271559 2204
rect 271559 2148 271563 2204
rect 271499 2144 271563 2148
rect 271579 2204 271643 2208
rect 271579 2148 271583 2204
rect 271583 2148 271639 2204
rect 271639 2148 271643 2204
rect 271579 2144 271643 2148
rect 267596 2076 267660 2140
rect 140268 1864 140332 1868
rect 140268 1808 140282 1864
rect 140282 1808 140332 1864
rect 34750 1660 34814 1664
rect 34750 1604 34754 1660
rect 34754 1604 34810 1660
rect 34810 1604 34814 1660
rect 34750 1600 34814 1604
rect 34830 1660 34894 1664
rect 34830 1604 34834 1660
rect 34834 1604 34890 1660
rect 34890 1604 34894 1660
rect 34830 1600 34894 1604
rect 34910 1660 34974 1664
rect 34910 1604 34914 1660
rect 34914 1604 34970 1660
rect 34970 1604 34974 1660
rect 34910 1600 34974 1604
rect 34990 1660 35054 1664
rect 34990 1604 34994 1660
rect 34994 1604 35050 1660
rect 35050 1604 35054 1660
rect 34990 1600 35054 1604
rect 19932 1532 19996 1596
rect 32444 1532 32508 1596
rect 57836 1532 57900 1596
rect 59308 1592 59372 1596
rect 59308 1536 59358 1592
rect 59358 1536 59372 1592
rect 59308 1532 59372 1536
rect 102347 1660 102411 1664
rect 102347 1604 102351 1660
rect 102351 1604 102407 1660
rect 102407 1604 102411 1660
rect 102347 1600 102411 1604
rect 102427 1660 102491 1664
rect 102427 1604 102431 1660
rect 102431 1604 102487 1660
rect 102487 1604 102491 1660
rect 102427 1600 102491 1604
rect 102507 1660 102571 1664
rect 102507 1604 102511 1660
rect 102511 1604 102567 1660
rect 102567 1604 102571 1660
rect 102507 1600 102571 1604
rect 102587 1660 102651 1664
rect 102587 1604 102591 1660
rect 102591 1604 102647 1660
rect 102647 1604 102651 1660
rect 102587 1600 102651 1604
rect 91140 1592 91204 1596
rect 91140 1536 91190 1592
rect 91190 1536 91204 1592
rect 91140 1532 91204 1536
rect 96292 1592 96356 1596
rect 96292 1536 96306 1592
rect 96306 1536 96356 1592
rect 96292 1532 96356 1536
rect 98500 1532 98564 1596
rect 20668 1396 20732 1460
rect 4476 1320 4540 1324
rect 4476 1264 4526 1320
rect 4526 1264 4540 1320
rect 4476 1260 4540 1264
rect 6684 1320 6748 1324
rect 6684 1264 6734 1320
rect 6734 1264 6748 1320
rect 6684 1260 6748 1264
rect 14780 1320 14844 1324
rect 14780 1264 14830 1320
rect 14830 1264 14844 1320
rect 14780 1260 14844 1264
rect 23612 1320 23676 1324
rect 23612 1264 23626 1320
rect 23626 1264 23676 1320
rect 23612 1260 23676 1264
rect 24348 1260 24412 1324
rect 25820 1320 25884 1324
rect 25820 1264 25834 1320
rect 25834 1264 25884 1320
rect 25820 1260 25884 1264
rect 26556 1320 26620 1324
rect 26556 1264 26570 1320
rect 26570 1264 26620 1320
rect 26556 1260 26620 1264
rect 76420 1320 76484 1324
rect 76420 1264 76470 1320
rect 76470 1264 76484 1320
rect 76420 1260 76484 1264
rect 78628 1320 78692 1324
rect 78628 1264 78678 1320
rect 78678 1264 78692 1320
rect 78628 1260 78692 1264
rect 81572 1320 81636 1324
rect 81572 1264 81622 1320
rect 81622 1264 81636 1320
rect 81572 1260 81636 1264
rect 83780 1320 83844 1324
rect 83780 1264 83830 1320
rect 83830 1264 83844 1320
rect 83780 1260 83844 1264
rect 88196 1396 88260 1460
rect 140268 1804 140332 1808
rect 194364 1804 194428 1868
rect 195836 1804 195900 1868
rect 212212 1804 212276 1868
rect 169944 1660 170008 1664
rect 169944 1604 169948 1660
rect 169948 1604 170004 1660
rect 170004 1604 170008 1660
rect 169944 1600 170008 1604
rect 170024 1660 170088 1664
rect 170024 1604 170028 1660
rect 170028 1604 170084 1660
rect 170084 1604 170088 1660
rect 170024 1600 170088 1604
rect 170104 1660 170168 1664
rect 170104 1604 170108 1660
rect 170108 1604 170164 1660
rect 170164 1604 170168 1660
rect 170104 1600 170168 1604
rect 170184 1660 170248 1664
rect 170184 1604 170188 1660
rect 170188 1604 170244 1660
rect 170244 1604 170248 1660
rect 170184 1600 170248 1604
rect 237541 1660 237605 1664
rect 237541 1604 237545 1660
rect 237545 1604 237601 1660
rect 237601 1604 237605 1660
rect 237541 1600 237605 1604
rect 237621 1660 237685 1664
rect 237621 1604 237625 1660
rect 237625 1604 237681 1660
rect 237681 1604 237685 1660
rect 237621 1600 237685 1604
rect 237701 1660 237765 1664
rect 237701 1604 237705 1660
rect 237705 1604 237761 1660
rect 237761 1604 237765 1660
rect 237701 1600 237765 1604
rect 237781 1660 237845 1664
rect 237781 1604 237785 1660
rect 237785 1604 237841 1660
rect 237841 1604 237845 1660
rect 237781 1600 237845 1604
rect 237236 1532 237300 1596
rect 113588 1396 113652 1460
rect 114876 1456 114940 1460
rect 114876 1400 114890 1456
rect 114890 1400 114940 1456
rect 114876 1396 114940 1400
rect 115612 1456 115676 1460
rect 115612 1400 115626 1456
rect 115626 1400 115676 1456
rect 115612 1396 115676 1400
rect 117268 1456 117332 1460
rect 117268 1400 117318 1456
rect 117318 1400 117332 1456
rect 117268 1396 117332 1400
rect 126836 1396 126900 1460
rect 128308 1396 128372 1460
rect 134932 1396 134996 1460
rect 137324 1396 137388 1460
rect 141004 1396 141068 1460
rect 150572 1456 150636 1460
rect 150572 1400 150622 1456
rect 150622 1400 150636 1456
rect 150572 1396 150636 1400
rect 152044 1456 152108 1460
rect 152044 1400 152094 1456
rect 152094 1400 152108 1456
rect 152044 1396 152108 1400
rect 155724 1396 155788 1460
rect 157196 1456 157260 1460
rect 157196 1400 157246 1456
rect 157246 1400 157260 1456
rect 157196 1396 157260 1400
rect 168236 1396 168300 1460
rect 186268 1456 186332 1460
rect 186268 1400 186318 1456
rect 186318 1400 186332 1456
rect 186268 1396 186332 1400
rect 197308 1456 197372 1460
rect 197308 1400 197358 1456
rect 197358 1400 197372 1456
rect 197308 1396 197372 1400
rect 201724 1396 201788 1460
rect 210004 1396 210068 1460
rect 218100 1396 218164 1460
rect 219572 1396 219636 1460
rect 222516 1456 222580 1460
rect 222516 1400 222566 1456
rect 222566 1400 222580 1456
rect 222516 1396 222580 1400
rect 226196 1396 226260 1460
rect 249380 1532 249444 1596
rect 251588 1532 251652 1596
rect 256740 1532 256804 1596
rect 242756 1456 242820 1460
rect 242756 1400 242806 1456
rect 242806 1400 242820 1456
rect 242756 1396 242820 1400
rect 245700 1456 245764 1460
rect 245700 1400 245750 1456
rect 245750 1400 245764 1456
rect 245700 1396 245764 1400
rect 248644 1396 248708 1460
rect 252324 1396 252388 1460
rect 257476 1456 257540 1460
rect 257476 1400 257526 1456
rect 257526 1400 257540 1456
rect 88932 1260 88996 1324
rect 89852 1260 89916 1324
rect 90404 1260 90468 1324
rect 91876 1260 91940 1324
rect 93348 1260 93412 1324
rect 152780 1260 152844 1324
rect 157932 1260 157996 1324
rect 257476 1396 257540 1400
rect 29500 1124 29564 1188
rect 158668 1124 158732 1188
rect 160140 1124 160204 1188
rect 161612 1184 161676 1188
rect 161612 1128 161662 1184
rect 161662 1128 161676 1184
rect 161612 1124 161676 1128
rect 163820 1184 163884 1188
rect 163820 1128 163870 1184
rect 163870 1128 163884 1184
rect 163820 1124 163884 1128
rect 165292 1184 165356 1188
rect 165292 1128 165306 1184
rect 165306 1128 165356 1184
rect 165292 1124 165356 1128
rect 166028 1184 166092 1188
rect 166028 1128 166042 1184
rect 166042 1128 166092 1184
rect 166028 1124 166092 1128
rect 166764 1184 166828 1188
rect 166764 1128 166814 1184
rect 166814 1128 166828 1184
rect 166764 1124 166828 1128
rect 223988 1124 224052 1188
rect 225460 1124 225524 1188
rect 227668 1124 227732 1188
rect 229876 1124 229940 1188
rect 230612 1124 230676 1188
rect 232084 1124 232148 1188
rect 232820 1124 232884 1188
rect 235028 1124 235092 1188
rect 236500 1124 236564 1188
rect 68548 1116 68612 1120
rect 68548 1060 68552 1116
rect 68552 1060 68608 1116
rect 68608 1060 68612 1116
rect 68548 1056 68612 1060
rect 68628 1116 68692 1120
rect 68628 1060 68632 1116
rect 68632 1060 68688 1116
rect 68688 1060 68692 1116
rect 68628 1056 68692 1060
rect 68708 1116 68772 1120
rect 68708 1060 68712 1116
rect 68712 1060 68768 1116
rect 68768 1060 68772 1116
rect 68708 1056 68772 1060
rect 68788 1116 68852 1120
rect 68788 1060 68792 1116
rect 68792 1060 68848 1116
rect 68848 1060 68852 1116
rect 68788 1056 68852 1060
rect 136145 1116 136209 1120
rect 136145 1060 136149 1116
rect 136149 1060 136205 1116
rect 136205 1060 136209 1116
rect 136145 1056 136209 1060
rect 136225 1116 136289 1120
rect 136225 1060 136229 1116
rect 136229 1060 136285 1116
rect 136285 1060 136289 1116
rect 136225 1056 136289 1060
rect 136305 1116 136369 1120
rect 136305 1060 136309 1116
rect 136309 1060 136365 1116
rect 136365 1060 136369 1116
rect 136305 1056 136369 1060
rect 136385 1116 136449 1120
rect 136385 1060 136389 1116
rect 136389 1060 136445 1116
rect 136445 1060 136449 1116
rect 136385 1056 136449 1060
rect 203742 1116 203806 1120
rect 203742 1060 203746 1116
rect 203746 1060 203802 1116
rect 203802 1060 203806 1116
rect 203742 1056 203806 1060
rect 203822 1116 203886 1120
rect 203822 1060 203826 1116
rect 203826 1060 203882 1116
rect 203882 1060 203886 1116
rect 203822 1056 203886 1060
rect 203902 1116 203966 1120
rect 203902 1060 203906 1116
rect 203906 1060 203962 1116
rect 203962 1060 203966 1116
rect 203902 1056 203966 1060
rect 203982 1116 204046 1120
rect 203982 1060 203986 1116
rect 203986 1060 204042 1116
rect 204042 1060 204046 1116
rect 203982 1056 204046 1060
rect 271339 1116 271403 1120
rect 271339 1060 271343 1116
rect 271343 1060 271399 1116
rect 271399 1060 271403 1116
rect 271339 1056 271403 1060
rect 271419 1116 271483 1120
rect 271419 1060 271423 1116
rect 271423 1060 271479 1116
rect 271479 1060 271483 1116
rect 271419 1056 271483 1060
rect 271499 1116 271563 1120
rect 271499 1060 271503 1116
rect 271503 1060 271559 1116
rect 271559 1060 271563 1116
rect 271499 1056 271563 1060
rect 271579 1116 271643 1120
rect 271579 1060 271583 1116
rect 271583 1060 271639 1116
rect 271639 1060 271643 1116
rect 271579 1056 271643 1060
rect 1532 988 1596 1052
rect 3740 1048 3804 1052
rect 3740 992 3790 1048
rect 3790 992 3804 1048
rect 3740 988 3804 992
rect 5212 1048 5276 1052
rect 5212 992 5226 1048
rect 5226 992 5276 1048
rect 5212 988 5276 992
rect 7420 988 7484 1052
rect 9628 1048 9692 1052
rect 9628 992 9678 1048
rect 9678 992 9692 1048
rect 9628 988 9692 992
rect 11836 988 11900 1052
rect 12572 988 12636 1052
rect 14044 1048 14108 1052
rect 14044 992 14094 1048
rect 14094 992 14108 1048
rect 14044 988 14108 992
rect 15516 1048 15580 1052
rect 15516 992 15530 1048
rect 15530 992 15580 1048
rect 15516 988 15580 992
rect 17724 988 17788 1052
rect 71268 988 71332 1052
rect 72004 988 72068 1052
rect 73476 988 73540 1052
rect 75684 1048 75748 1052
rect 75684 992 75734 1048
rect 75734 992 75748 1048
rect 75684 988 75748 992
rect 77156 1048 77220 1052
rect 77156 992 77206 1048
rect 77206 992 77220 1048
rect 77156 988 77220 992
rect 79364 1048 79428 1052
rect 79364 992 79414 1048
rect 79414 992 79428 1048
rect 79364 988 79428 992
rect 80836 1048 80900 1052
rect 80836 992 80886 1048
rect 80886 992 80900 1048
rect 80836 988 80900 992
rect 82308 1048 82372 1052
rect 82308 992 82358 1048
rect 82358 992 82372 1048
rect 82308 988 82372 992
rect 84516 1048 84580 1052
rect 84516 992 84566 1048
rect 84566 992 84580 1048
rect 84516 988 84580 992
rect 85988 1048 86052 1052
rect 85988 992 86038 1048
rect 86038 992 86052 1048
rect 85988 988 86052 992
rect 69060 912 69124 916
rect 69060 856 69110 912
rect 69110 856 69124 912
rect 69060 852 69124 856
rect 69796 852 69860 916
rect 70532 852 70596 916
rect 72740 852 72804 916
rect 74212 912 74276 916
rect 74212 856 74262 912
rect 74262 856 74276 912
rect 74212 852 74276 856
rect 74948 852 75012 916
rect 77892 852 77956 916
rect 80100 852 80164 916
rect 83044 852 83108 916
rect 86724 912 86788 916
rect 86724 856 86774 912
rect 86774 856 86788 912
rect 86724 852 86788 856
rect 139532 988 139596 1052
rect 99236 852 99300 916
rect 3004 776 3068 780
rect 3004 720 3018 776
rect 3018 720 3068 776
rect 3004 716 3068 720
rect 5948 716 6012 780
rect 10364 776 10428 780
rect 10364 720 10378 776
rect 10378 720 10428 776
rect 10364 716 10428 720
rect 11100 716 11164 780
rect 16252 716 16316 780
rect 16988 776 17052 780
rect 16988 720 17038 776
rect 17038 720 17052 776
rect 16988 716 17052 720
rect 2268 580 2332 644
rect 13308 580 13372 644
rect 21404 640 21468 644
rect 21404 584 21454 640
rect 21454 584 21468 640
rect 21404 580 21468 584
rect 28028 580 28092 644
rect 30236 640 30300 644
rect 30236 584 30286 640
rect 30286 584 30300 640
rect 30236 580 30300 584
rect 30972 580 31036 644
rect 31708 580 31772 644
rect 34928 580 34992 644
rect 35664 640 35728 644
rect 35664 584 35678 640
rect 35678 584 35728 640
rect 35664 580 35728 584
rect 36400 580 36464 644
rect 37136 580 37200 644
rect 37872 580 37936 644
rect 38608 640 38672 644
rect 38608 584 38622 640
rect 38622 584 38672 640
rect 38608 580 38672 584
rect 40080 580 40144 644
rect 40816 640 40880 644
rect 40816 584 40830 640
rect 40830 584 40880 640
rect 40816 580 40880 584
rect 41552 580 41616 644
rect 42288 580 42352 644
rect 43024 580 43088 644
rect 43760 580 43824 644
rect 44496 580 44560 644
rect 45232 580 45296 644
rect 45968 640 46032 644
rect 45968 584 45982 640
rect 45982 584 46032 640
rect 45968 580 46032 584
rect 46704 580 46768 644
rect 47440 580 47504 644
rect 48176 640 48240 644
rect 48176 584 48226 640
rect 48226 584 48240 640
rect 48176 580 48240 584
rect 48912 580 48976 644
rect 49648 580 49712 644
rect 50384 580 50448 644
rect 51120 580 51184 644
rect 51856 580 51920 644
rect 53328 580 53392 644
rect 54064 580 54128 644
rect 8156 444 8220 508
rect 92612 580 92676 644
rect 94820 640 94884 644
rect 94820 584 94834 640
rect 94834 584 94884 640
rect 94820 580 94884 584
rect 99972 580 100036 644
rect 266308 988 266372 1052
rect 205588 852 205652 916
rect 206324 852 206388 916
rect 207060 852 207124 916
rect 208532 852 208596 916
rect 138796 776 138860 780
rect 138796 720 138846 776
rect 138846 720 138860 776
rect 138796 716 138860 720
rect 141740 776 141804 780
rect 141740 720 141790 776
rect 141790 720 141804 776
rect 141740 716 141804 720
rect 142476 716 142540 780
rect 146156 716 146220 780
rect 148364 776 148428 780
rect 148364 720 148414 776
rect 148414 720 148428 776
rect 148364 716 148428 720
rect 149836 716 149900 780
rect 151860 716 151924 780
rect 124536 580 124600 644
rect 125272 640 125336 644
rect 125272 584 125322 640
rect 125322 584 125336 640
rect 125272 580 125336 584
rect 126008 580 126072 644
rect 128952 580 129016 644
rect 130424 580 130488 644
rect 131160 580 131224 644
rect 134104 580 134168 644
rect 138060 580 138124 644
rect 143212 580 143276 644
rect 147628 580 147692 644
rect 151308 580 151372 644
rect 159404 580 159468 644
rect 162348 580 162412 644
rect 163084 580 163148 644
rect 164556 640 164620 644
rect 164556 584 164606 640
rect 164606 584 164620 640
rect 164556 580 164620 584
rect 168972 640 169036 644
rect 168972 584 169022 640
rect 169022 584 169036 640
rect 168972 580 169036 584
rect 171456 580 171520 644
rect 172192 640 172256 644
rect 172192 584 172242 640
rect 172242 584 172256 640
rect 172192 580 172256 584
rect 172928 640 172992 644
rect 172928 584 172978 640
rect 172978 584 172992 640
rect 172928 580 172992 584
rect 173664 580 173728 644
rect 174400 640 174464 644
rect 174400 584 174450 640
rect 174450 584 174464 640
rect 174400 580 174464 584
rect 175136 580 175200 644
rect 176608 640 176672 644
rect 176608 584 176658 640
rect 176658 584 176672 640
rect 176608 580 176672 584
rect 177344 580 177408 644
rect 178080 580 178144 644
rect 178816 580 178880 644
rect 179552 640 179616 644
rect 179552 584 179602 640
rect 179602 584 179616 640
rect 179552 580 179616 584
rect 180288 640 180352 644
rect 180288 584 180338 640
rect 180338 584 180352 640
rect 180288 580 180352 584
rect 215892 716 215956 780
rect 224724 776 224788 780
rect 224724 720 224774 776
rect 224774 720 224788 776
rect 224724 716 224788 720
rect 225092 716 225156 780
rect 55536 444 55600 508
rect 56272 444 56336 508
rect 57008 444 57072 508
rect 58480 444 58544 508
rect 59952 504 60016 508
rect 59952 448 60002 504
rect 60002 448 60016 504
rect 59952 444 60016 448
rect 60688 444 60752 508
rect 61424 504 61488 508
rect 61424 448 61474 504
rect 61474 448 61488 504
rect 61424 444 61488 448
rect 62160 444 62224 508
rect 62896 444 62960 508
rect 65840 504 65904 508
rect 65840 448 65890 504
rect 65890 448 65904 504
rect 65840 444 65904 448
rect 66576 444 66640 508
rect 87460 504 87524 508
rect 87460 448 87510 504
rect 87510 448 87524 504
rect 87460 444 87524 448
rect 8892 308 8956 372
rect 18460 308 18524 372
rect 28764 368 28828 372
rect 28764 312 28814 368
rect 28814 312 28828 368
rect 28764 308 28828 312
rect 39344 308 39408 372
rect 52592 308 52656 372
rect 63632 308 63696 372
rect 64368 308 64432 372
rect 65104 308 65168 372
rect 85252 308 85316 372
rect 117912 444 117976 508
rect 118648 504 118712 508
rect 118648 448 118698 504
rect 118698 448 118712 504
rect 118648 444 118712 448
rect 119384 504 119448 508
rect 119384 448 119398 504
rect 119398 448 119448 504
rect 119384 444 119448 448
rect 120120 444 120184 508
rect 120856 444 120920 508
rect 121592 444 121656 508
rect 122328 444 122392 508
rect 123064 444 123128 508
rect 127480 444 127544 508
rect 143948 504 144012 508
rect 143948 448 143998 504
rect 143998 448 144012 504
rect 143948 444 144012 448
rect 95188 308 95252 372
rect 129688 308 129752 372
rect 131896 308 131960 372
rect 132632 308 132696 372
rect 146892 368 146956 372
rect 146892 312 146942 368
rect 146942 312 146956 368
rect 146892 308 146956 312
rect 153148 172 153212 236
rect 160876 308 160940 372
rect 167500 308 167564 372
rect 175872 444 175936 508
rect 181760 504 181824 508
rect 181760 448 181810 504
rect 181810 448 181824 504
rect 181760 444 181824 448
rect 182496 444 182560 508
rect 183232 504 183296 508
rect 183232 448 183282 504
rect 183282 448 183296 504
rect 183232 444 183296 448
rect 183968 444 184032 508
rect 184704 504 184768 508
rect 184704 448 184754 504
rect 184754 448 184768 504
rect 184704 444 184768 448
rect 185440 504 185504 508
rect 185440 448 185490 504
rect 185490 448 185504 504
rect 185440 444 185504 448
rect 186912 504 186976 508
rect 186912 448 186962 504
rect 186962 448 186976 504
rect 186912 444 186976 448
rect 187648 444 187712 508
rect 188384 444 188448 508
rect 189120 444 189184 508
rect 190592 444 190656 508
rect 192800 504 192864 508
rect 192800 448 192850 504
rect 192850 448 192864 504
rect 192800 444 192864 448
rect 193536 504 193600 508
rect 193536 448 193586 504
rect 193586 448 193600 504
rect 193536 444 193600 448
rect 195008 444 195072 508
rect 196480 444 196544 508
rect 198688 444 198752 508
rect 200160 444 200224 508
rect 202368 504 202432 508
rect 202368 448 202418 504
rect 202418 448 202432 504
rect 202368 444 202432 448
rect 203104 444 203168 508
rect 209268 444 209332 508
rect 213684 444 213748 508
rect 181024 308 181088 372
rect 192064 308 192128 372
rect 207796 308 207860 372
rect 212948 368 213012 372
rect 212948 312 212998 368
rect 212998 312 213012 368
rect 212948 308 213012 312
rect 214420 368 214484 372
rect 214420 312 214470 368
rect 214470 312 214484 368
rect 214420 308 214484 312
rect 221780 580 221844 644
rect 226932 580 226996 644
rect 228404 580 228468 644
rect 229140 580 229204 644
rect 231348 580 231412 644
rect 233556 580 233620 644
rect 234292 580 234356 644
rect 235764 640 235828 644
rect 235764 584 235814 640
rect 235814 584 235828 640
rect 235764 580 235828 584
rect 239720 580 239784 644
rect 240456 580 240520 644
rect 241192 640 241256 644
rect 241192 584 241242 640
rect 241242 584 241256 640
rect 241192 580 241256 584
rect 241928 640 241992 644
rect 241928 584 241978 640
rect 241978 584 241992 640
rect 241928 580 241992 584
rect 243400 640 243464 644
rect 243400 584 243450 640
rect 243450 584 243464 640
rect 243400 580 243464 584
rect 244136 640 244200 644
rect 244136 584 244186 640
rect 244186 584 244200 640
rect 244136 580 244200 584
rect 244872 640 244936 644
rect 244872 584 244922 640
rect 244922 584 244936 640
rect 244872 580 244936 584
rect 247080 640 247144 644
rect 247080 584 247094 640
rect 247094 584 247144 640
rect 247080 580 247144 584
rect 247816 580 247880 644
rect 250024 640 250088 644
rect 250024 584 250074 640
rect 250074 584 250088 640
rect 250024 580 250088 584
rect 254440 580 254504 644
rect 255176 580 255240 644
rect 258120 640 258184 644
rect 258120 584 258134 640
rect 258134 584 258184 640
rect 258120 580 258184 584
rect 261064 640 261128 644
rect 261064 584 261114 640
rect 261114 584 261128 640
rect 261064 580 261128 584
rect 262536 580 262600 644
rect 263272 640 263336 644
rect 263272 584 263322 640
rect 263322 584 263336 640
rect 263272 580 263336 584
rect 264008 580 264072 644
rect 264744 580 264808 644
rect 265480 580 265544 644
rect 266216 580 266280 644
rect 266952 640 267016 644
rect 266952 584 266966 640
rect 266966 584 267016 640
rect 266952 580 267016 584
rect 267688 640 267752 644
rect 267688 584 267702 640
rect 267702 584 267752 640
rect 267688 580 267752 584
rect 268424 640 268488 644
rect 268424 584 268438 640
rect 268438 584 268488 640
rect 268424 580 268488 584
rect 269160 580 269224 644
rect 270632 580 270696 644
rect 252968 444 253032 508
rect 220308 308 220372 372
rect 253704 308 253768 372
rect 269896 308 269960 372
<< metal4 >>
rect 798 9213 858 10880
rect 1534 10165 1594 10880
rect 2270 10165 2330 10880
rect 1531 10164 1597 10165
rect 1531 10100 1532 10164
rect 1596 10100 1597 10164
rect 1531 10099 1597 10100
rect 2267 10164 2333 10165
rect 2267 10100 2268 10164
rect 2332 10100 2333 10164
rect 2267 10099 2333 10100
rect 3006 9893 3066 10880
rect 3742 10165 3802 10880
rect 4478 10165 4538 10880
rect 5214 10165 5274 10880
rect 5950 10165 6010 10880
rect 6686 10165 6746 10880
rect 7422 10165 7482 10880
rect 3739 10164 3805 10165
rect 3739 10100 3740 10164
rect 3804 10100 3805 10164
rect 3739 10099 3805 10100
rect 4475 10164 4541 10165
rect 4475 10100 4476 10164
rect 4540 10100 4541 10164
rect 4475 10099 4541 10100
rect 5211 10164 5277 10165
rect 5211 10100 5212 10164
rect 5276 10100 5277 10164
rect 5211 10099 5277 10100
rect 5947 10164 6013 10165
rect 5947 10100 5948 10164
rect 6012 10100 6013 10164
rect 5947 10099 6013 10100
rect 6683 10164 6749 10165
rect 6683 10100 6684 10164
rect 6748 10100 6749 10164
rect 6683 10099 6749 10100
rect 7419 10164 7485 10165
rect 7419 10100 7420 10164
rect 7484 10100 7485 10164
rect 7419 10099 7485 10100
rect 8158 9893 8218 10880
rect 8894 10165 8954 10880
rect 9630 10165 9690 10880
rect 10366 10165 10426 10880
rect 11102 10165 11162 10880
rect 11838 10165 11898 10880
rect 12574 10165 12634 10880
rect 8891 10164 8957 10165
rect 8891 10100 8892 10164
rect 8956 10100 8957 10164
rect 8891 10099 8957 10100
rect 9627 10164 9693 10165
rect 9627 10100 9628 10164
rect 9692 10100 9693 10164
rect 9627 10099 9693 10100
rect 10363 10164 10429 10165
rect 10363 10100 10364 10164
rect 10428 10100 10429 10164
rect 10363 10099 10429 10100
rect 11099 10164 11165 10165
rect 11099 10100 11100 10164
rect 11164 10100 11165 10164
rect 11099 10099 11165 10100
rect 11835 10164 11901 10165
rect 11835 10100 11836 10164
rect 11900 10100 11901 10164
rect 11835 10099 11901 10100
rect 12571 10164 12637 10165
rect 12571 10100 12572 10164
rect 12636 10100 12637 10164
rect 12571 10099 12637 10100
rect 13310 9893 13370 10880
rect 14046 10165 14106 10880
rect 14782 10165 14842 10880
rect 15518 10165 15578 10880
rect 16254 10165 16314 10880
rect 16990 10165 17050 10880
rect 17726 10165 17786 10880
rect 18462 10165 18522 10880
rect 14043 10164 14109 10165
rect 14043 10100 14044 10164
rect 14108 10100 14109 10164
rect 14043 10099 14109 10100
rect 14779 10164 14845 10165
rect 14779 10100 14780 10164
rect 14844 10100 14845 10164
rect 14779 10099 14845 10100
rect 15515 10164 15581 10165
rect 15515 10100 15516 10164
rect 15580 10100 15581 10164
rect 15515 10099 15581 10100
rect 16251 10164 16317 10165
rect 16251 10100 16252 10164
rect 16316 10100 16317 10164
rect 16251 10099 16317 10100
rect 16987 10164 17053 10165
rect 16987 10100 16988 10164
rect 17052 10100 17053 10164
rect 16987 10099 17053 10100
rect 17723 10164 17789 10165
rect 17723 10100 17724 10164
rect 17788 10100 17789 10164
rect 17723 10099 17789 10100
rect 18459 10164 18525 10165
rect 18459 10100 18460 10164
rect 18524 10100 18525 10164
rect 18459 10099 18525 10100
rect 3003 9892 3069 9893
rect 3003 9828 3004 9892
rect 3068 9828 3069 9892
rect 3003 9827 3069 9828
rect 8155 9892 8221 9893
rect 8155 9828 8156 9892
rect 8220 9828 8221 9892
rect 8155 9827 8221 9828
rect 13307 9892 13373 9893
rect 13307 9828 13308 9892
rect 13372 9828 13373 9892
rect 13307 9827 13373 9828
rect 795 9212 861 9213
rect 795 9148 796 9212
rect 860 9148 861 9212
rect 795 9147 861 9148
rect 19198 6901 19258 10880
rect 19934 9893 19994 10880
rect 19931 9892 19997 9893
rect 19931 9828 19932 9892
rect 19996 9828 19997 9892
rect 19931 9827 19997 9828
rect 20670 8397 20730 10880
rect 21406 8669 21466 10880
rect 22142 8941 22202 10880
rect 22139 8940 22205 8941
rect 22139 8876 22140 8940
rect 22204 8876 22205 8940
rect 22139 8875 22205 8876
rect 21403 8668 21469 8669
rect 21403 8604 21404 8668
rect 21468 8604 21469 8668
rect 21403 8603 21469 8604
rect 22878 8397 22938 10880
rect 23614 8397 23674 10880
rect 24350 9213 24410 10880
rect 24347 9212 24413 9213
rect 24347 9148 24348 9212
rect 24412 9148 24413 9212
rect 24347 9147 24413 9148
rect 25086 8397 25146 10880
rect 25822 9757 25882 10880
rect 26558 9757 26618 10880
rect 25819 9756 25885 9757
rect 25819 9692 25820 9756
rect 25884 9692 25885 9756
rect 25819 9691 25885 9692
rect 26555 9756 26621 9757
rect 26555 9692 26556 9756
rect 26620 9692 26621 9756
rect 26555 9691 26621 9692
rect 27294 8669 27354 10880
rect 28030 8669 28090 10880
rect 28766 8669 28826 10880
rect 29502 9757 29562 10880
rect 30238 9757 30298 10880
rect 29499 9756 29565 9757
rect 29499 9692 29500 9756
rect 29564 9692 29565 9756
rect 29499 9691 29565 9692
rect 30235 9756 30301 9757
rect 30235 9692 30236 9756
rect 30300 9692 30301 9756
rect 30235 9691 30301 9692
rect 30974 8669 31034 10880
rect 31710 10301 31770 10880
rect 31707 10300 31773 10301
rect 31707 10236 31708 10300
rect 31772 10236 31773 10300
rect 31707 10235 31773 10236
rect 32446 9213 32506 10880
rect 34930 10301 34990 10880
rect 35666 10301 35726 10880
rect 36402 10301 36462 10880
rect 37138 10301 37198 10880
rect 37874 10301 37934 10880
rect 38610 10301 38670 10880
rect 39346 10301 39406 10880
rect 40082 10301 40142 10880
rect 40818 10301 40878 10880
rect 41554 10301 41614 10880
rect 42290 10301 42350 10880
rect 43026 10301 43086 10880
rect 43762 10301 43822 10880
rect 44498 10301 44558 10880
rect 45234 10301 45294 10880
rect 45970 10301 46030 10880
rect 46706 10301 46766 10880
rect 47442 10301 47502 10880
rect 48178 10301 48238 10880
rect 48914 10301 48974 10880
rect 49650 10301 49710 10880
rect 50386 10301 50446 10880
rect 51122 10301 51182 10880
rect 51858 10301 51918 10880
rect 52594 10573 52654 10880
rect 52591 10572 52657 10573
rect 52591 10508 52592 10572
rect 52656 10508 52657 10572
rect 52591 10507 52657 10508
rect 53330 10301 53390 10880
rect 54066 10301 54126 10880
rect 54802 10301 54862 10880
rect 55538 10301 55598 10880
rect 56274 10301 56334 10880
rect 57010 10301 57070 10880
rect 57746 10301 57806 10880
rect 58482 10301 58542 10880
rect 59218 10301 59278 10880
rect 59954 10301 60014 10880
rect 60690 10301 60750 10880
rect 61426 10301 61486 10880
rect 62162 10301 62222 10880
rect 62898 10301 62958 10880
rect 63634 10301 63694 10880
rect 64370 10301 64430 10880
rect 65106 10301 65166 10880
rect 65842 10301 65902 10880
rect 66578 10301 66638 10880
rect 34927 10300 34993 10301
rect 34927 10236 34928 10300
rect 34992 10236 34993 10300
rect 34927 10235 34993 10236
rect 35663 10300 35729 10301
rect 35663 10236 35664 10300
rect 35728 10236 35729 10300
rect 35663 10235 35729 10236
rect 36399 10300 36465 10301
rect 36399 10236 36400 10300
rect 36464 10236 36465 10300
rect 36399 10235 36465 10236
rect 37135 10300 37201 10301
rect 37135 10236 37136 10300
rect 37200 10236 37201 10300
rect 37135 10235 37201 10236
rect 37871 10300 37937 10301
rect 37871 10236 37872 10300
rect 37936 10236 37937 10300
rect 37871 10235 37937 10236
rect 38607 10300 38673 10301
rect 38607 10236 38608 10300
rect 38672 10236 38673 10300
rect 38607 10235 38673 10236
rect 39343 10300 39409 10301
rect 39343 10236 39344 10300
rect 39408 10236 39409 10300
rect 39343 10235 39409 10236
rect 40079 10300 40145 10301
rect 40079 10236 40080 10300
rect 40144 10236 40145 10300
rect 40079 10235 40145 10236
rect 40815 10300 40881 10301
rect 40815 10236 40816 10300
rect 40880 10236 40881 10300
rect 40815 10235 40881 10236
rect 41551 10300 41617 10301
rect 41551 10236 41552 10300
rect 41616 10236 41617 10300
rect 41551 10235 41617 10236
rect 42287 10300 42353 10301
rect 42287 10236 42288 10300
rect 42352 10236 42353 10300
rect 42287 10235 42353 10236
rect 43023 10300 43089 10301
rect 43023 10236 43024 10300
rect 43088 10236 43089 10300
rect 43023 10235 43089 10236
rect 43759 10300 43825 10301
rect 43759 10236 43760 10300
rect 43824 10236 43825 10300
rect 43759 10235 43825 10236
rect 44495 10300 44561 10301
rect 44495 10236 44496 10300
rect 44560 10236 44561 10300
rect 44495 10235 44561 10236
rect 45231 10300 45297 10301
rect 45231 10236 45232 10300
rect 45296 10236 45297 10300
rect 45231 10235 45297 10236
rect 45967 10300 46033 10301
rect 45967 10236 45968 10300
rect 46032 10236 46033 10300
rect 45967 10235 46033 10236
rect 46703 10300 46769 10301
rect 46703 10236 46704 10300
rect 46768 10236 46769 10300
rect 46703 10235 46769 10236
rect 47439 10300 47505 10301
rect 47439 10236 47440 10300
rect 47504 10236 47505 10300
rect 47439 10235 47505 10236
rect 48175 10300 48241 10301
rect 48175 10236 48176 10300
rect 48240 10236 48241 10300
rect 48175 10235 48241 10236
rect 48911 10300 48977 10301
rect 48911 10236 48912 10300
rect 48976 10236 48977 10300
rect 48911 10235 48977 10236
rect 49647 10300 49713 10301
rect 49647 10236 49648 10300
rect 49712 10236 49713 10300
rect 49647 10235 49713 10236
rect 50383 10300 50449 10301
rect 50383 10236 50384 10300
rect 50448 10236 50449 10300
rect 50383 10235 50449 10236
rect 51119 10300 51185 10301
rect 51119 10236 51120 10300
rect 51184 10236 51185 10300
rect 51119 10235 51185 10236
rect 51855 10300 51921 10301
rect 51855 10236 51856 10300
rect 51920 10236 51921 10300
rect 51855 10235 51921 10236
rect 53327 10300 53393 10301
rect 53327 10236 53328 10300
rect 53392 10236 53393 10300
rect 53327 10235 53393 10236
rect 54063 10300 54129 10301
rect 54063 10236 54064 10300
rect 54128 10236 54129 10300
rect 54063 10235 54129 10236
rect 54799 10300 54865 10301
rect 54799 10236 54800 10300
rect 54864 10236 54865 10300
rect 54799 10235 54865 10236
rect 55535 10300 55601 10301
rect 55535 10236 55536 10300
rect 55600 10236 55601 10300
rect 55535 10235 55601 10236
rect 56271 10300 56337 10301
rect 56271 10236 56272 10300
rect 56336 10236 56337 10300
rect 56271 10235 56337 10236
rect 57007 10300 57073 10301
rect 57007 10236 57008 10300
rect 57072 10236 57073 10300
rect 57007 10235 57073 10236
rect 57743 10300 57809 10301
rect 57743 10236 57744 10300
rect 57808 10236 57809 10300
rect 57743 10235 57809 10236
rect 58479 10300 58545 10301
rect 58479 10236 58480 10300
rect 58544 10236 58545 10300
rect 58479 10235 58545 10236
rect 59215 10300 59281 10301
rect 59215 10236 59216 10300
rect 59280 10236 59281 10300
rect 59215 10235 59281 10236
rect 59951 10300 60017 10301
rect 59951 10236 59952 10300
rect 60016 10236 60017 10300
rect 59951 10235 60017 10236
rect 60687 10300 60753 10301
rect 60687 10236 60688 10300
rect 60752 10236 60753 10300
rect 60687 10235 60753 10236
rect 61423 10300 61489 10301
rect 61423 10236 61424 10300
rect 61488 10236 61489 10300
rect 61423 10235 61489 10236
rect 62159 10300 62225 10301
rect 62159 10236 62160 10300
rect 62224 10236 62225 10300
rect 62159 10235 62225 10236
rect 62895 10300 62961 10301
rect 62895 10236 62896 10300
rect 62960 10236 62961 10300
rect 62895 10235 62961 10236
rect 63631 10300 63697 10301
rect 63631 10236 63632 10300
rect 63696 10236 63697 10300
rect 63631 10235 63697 10236
rect 64367 10300 64433 10301
rect 64367 10236 64368 10300
rect 64432 10236 64433 10300
rect 64367 10235 64433 10236
rect 65103 10300 65169 10301
rect 65103 10236 65104 10300
rect 65168 10236 65169 10300
rect 65103 10235 65169 10236
rect 65839 10300 65905 10301
rect 65839 10236 65840 10300
rect 65904 10236 65905 10300
rect 65839 10235 65905 10236
rect 66575 10300 66641 10301
rect 66575 10236 66576 10300
rect 66640 10236 66641 10300
rect 66575 10235 66641 10236
rect 34742 9280 35062 9840
rect 34742 9216 34750 9280
rect 34814 9216 34830 9280
rect 34894 9216 34910 9280
rect 34974 9216 34990 9280
rect 35054 9216 35062 9280
rect 32443 9212 32509 9213
rect 32443 9148 32444 9212
rect 32508 9148 32509 9212
rect 32443 9147 32509 9148
rect 27291 8668 27357 8669
rect 27291 8604 27292 8668
rect 27356 8604 27357 8668
rect 27291 8603 27357 8604
rect 28027 8668 28093 8669
rect 28027 8604 28028 8668
rect 28092 8604 28093 8668
rect 28027 8603 28093 8604
rect 28763 8668 28829 8669
rect 28763 8604 28764 8668
rect 28828 8604 28829 8668
rect 28763 8603 28829 8604
rect 30971 8668 31037 8669
rect 30971 8604 30972 8668
rect 31036 8604 31037 8668
rect 30971 8603 31037 8604
rect 20667 8396 20733 8397
rect 20667 8332 20668 8396
rect 20732 8332 20733 8396
rect 20667 8331 20733 8332
rect 22875 8396 22941 8397
rect 22875 8332 22876 8396
rect 22940 8332 22941 8396
rect 22875 8331 22941 8332
rect 23611 8396 23677 8397
rect 23611 8332 23612 8396
rect 23676 8332 23677 8396
rect 23611 8331 23677 8332
rect 25083 8396 25149 8397
rect 25083 8332 25084 8396
rect 25148 8332 25149 8396
rect 25083 8331 25149 8332
rect 34742 8192 35062 9216
rect 34742 8128 34750 8192
rect 34814 8128 34830 8192
rect 34894 8128 34910 8192
rect 34974 8128 34990 8192
rect 35054 8128 35062 8192
rect 34742 7104 35062 8128
rect 34742 7040 34750 7104
rect 34814 7040 34830 7104
rect 34894 7040 34910 7104
rect 34974 7040 34990 7104
rect 35054 7040 35062 7104
rect 19195 6900 19261 6901
rect 19195 6836 19196 6900
rect 19260 6836 19261 6900
rect 19195 6835 19261 6836
rect 34742 6016 35062 7040
rect 34742 5952 34750 6016
rect 34814 5952 34830 6016
rect 34894 5952 34910 6016
rect 34974 5952 34990 6016
rect 35054 5952 35062 6016
rect 34742 4928 35062 5952
rect 34742 4864 34750 4928
rect 34814 4864 34830 4928
rect 34894 4864 34910 4928
rect 34974 4864 34990 4928
rect 35054 4864 35062 4928
rect 34742 3840 35062 4864
rect 34742 3776 34750 3840
rect 34814 3776 34830 3840
rect 34894 3776 34910 3840
rect 34974 3776 34990 3840
rect 35054 3776 35062 3840
rect 795 2820 861 2821
rect 795 2756 796 2820
rect 860 2756 861 2820
rect 795 2755 861 2756
rect 19195 2820 19261 2821
rect 19195 2756 19196 2820
rect 19260 2756 19261 2820
rect 19195 2755 19261 2756
rect 22875 2820 22941 2821
rect 22875 2756 22876 2820
rect 22940 2756 22941 2820
rect 22875 2755 22941 2756
rect 25083 2820 25149 2821
rect 25083 2756 25084 2820
rect 25148 2756 25149 2820
rect 25083 2755 25149 2756
rect 27291 2820 27357 2821
rect 27291 2756 27292 2820
rect 27356 2756 27357 2820
rect 27291 2755 27357 2756
rect 798 0 858 2755
rect 4475 1324 4541 1325
rect 4475 1260 4476 1324
rect 4540 1260 4541 1324
rect 4475 1259 4541 1260
rect 6683 1324 6749 1325
rect 6683 1260 6684 1324
rect 6748 1260 6749 1324
rect 6683 1259 6749 1260
rect 14779 1324 14845 1325
rect 14779 1260 14780 1324
rect 14844 1260 14845 1324
rect 14779 1259 14845 1260
rect 1531 1052 1597 1053
rect 1531 988 1532 1052
rect 1596 988 1597 1052
rect 1531 987 1597 988
rect 3739 1052 3805 1053
rect 3739 988 3740 1052
rect 3804 988 3805 1052
rect 3739 987 3805 988
rect 1534 0 1594 987
rect 3003 780 3069 781
rect 3003 716 3004 780
rect 3068 716 3069 780
rect 3003 715 3069 716
rect 2267 644 2333 645
rect 2267 580 2268 644
rect 2332 580 2333 644
rect 2267 579 2333 580
rect 2270 0 2330 579
rect 3006 0 3066 715
rect 3742 0 3802 987
rect 4478 0 4538 1259
rect 5211 1052 5277 1053
rect 5211 988 5212 1052
rect 5276 988 5277 1052
rect 5211 987 5277 988
rect 5214 0 5274 987
rect 5947 780 6013 781
rect 5947 716 5948 780
rect 6012 716 6013 780
rect 5947 715 6013 716
rect 5950 0 6010 715
rect 6686 0 6746 1259
rect 7419 1052 7485 1053
rect 7419 988 7420 1052
rect 7484 988 7485 1052
rect 7419 987 7485 988
rect 9627 1052 9693 1053
rect 9627 988 9628 1052
rect 9692 988 9693 1052
rect 9627 987 9693 988
rect 11835 1052 11901 1053
rect 11835 988 11836 1052
rect 11900 988 11901 1052
rect 11835 987 11901 988
rect 12571 1052 12637 1053
rect 12571 988 12572 1052
rect 12636 988 12637 1052
rect 12571 987 12637 988
rect 14043 1052 14109 1053
rect 14043 988 14044 1052
rect 14108 988 14109 1052
rect 14043 987 14109 988
rect 7422 0 7482 987
rect 8155 508 8221 509
rect 8155 444 8156 508
rect 8220 444 8221 508
rect 8155 443 8221 444
rect 8158 0 8218 443
rect 8891 372 8957 373
rect 8891 308 8892 372
rect 8956 308 8957 372
rect 8891 307 8957 308
rect 8894 0 8954 307
rect 9630 0 9690 987
rect 10363 780 10429 781
rect 10363 716 10364 780
rect 10428 716 10429 780
rect 10363 715 10429 716
rect 11099 780 11165 781
rect 11099 716 11100 780
rect 11164 716 11165 780
rect 11099 715 11165 716
rect 10366 0 10426 715
rect 11102 0 11162 715
rect 11838 0 11898 987
rect 12574 0 12634 987
rect 13307 644 13373 645
rect 13307 580 13308 644
rect 13372 580 13373 644
rect 13307 579 13373 580
rect 13310 0 13370 579
rect 14046 0 14106 987
rect 14782 0 14842 1259
rect 15515 1052 15581 1053
rect 15515 988 15516 1052
rect 15580 988 15581 1052
rect 15515 987 15581 988
rect 17723 1052 17789 1053
rect 17723 988 17724 1052
rect 17788 988 17789 1052
rect 17723 987 17789 988
rect 15518 0 15578 987
rect 16251 780 16317 781
rect 16251 716 16252 780
rect 16316 716 16317 780
rect 16251 715 16317 716
rect 16987 780 17053 781
rect 16987 716 16988 780
rect 17052 716 17053 780
rect 16987 715 17053 716
rect 16254 0 16314 715
rect 16990 0 17050 715
rect 17726 0 17786 987
rect 18459 372 18525 373
rect 18459 308 18460 372
rect 18524 308 18525 372
rect 18459 307 18525 308
rect 18462 0 18522 307
rect 19198 0 19258 2755
rect 22139 1732 22205 1733
rect 22139 1668 22140 1732
rect 22204 1668 22205 1732
rect 22139 1667 22205 1668
rect 19931 1596 19997 1597
rect 19931 1532 19932 1596
rect 19996 1532 19997 1596
rect 19931 1531 19997 1532
rect 19934 0 19994 1531
rect 20667 1460 20733 1461
rect 20667 1396 20668 1460
rect 20732 1396 20733 1460
rect 20667 1395 20733 1396
rect 20670 0 20730 1395
rect 21403 644 21469 645
rect 21403 580 21404 644
rect 21468 580 21469 644
rect 21403 579 21469 580
rect 21406 0 21466 579
rect 22142 0 22202 1667
rect 22878 0 22938 2755
rect 23611 1324 23677 1325
rect 23611 1260 23612 1324
rect 23676 1260 23677 1324
rect 23611 1259 23677 1260
rect 24347 1324 24413 1325
rect 24347 1260 24348 1324
rect 24412 1260 24413 1324
rect 24347 1259 24413 1260
rect 23614 0 23674 1259
rect 24350 0 24410 1259
rect 25086 0 25146 2755
rect 25819 1324 25885 1325
rect 25819 1260 25820 1324
rect 25884 1260 25885 1324
rect 25819 1259 25885 1260
rect 26555 1324 26621 1325
rect 26555 1260 26556 1324
rect 26620 1260 26621 1324
rect 26555 1259 26621 1260
rect 25822 0 25882 1259
rect 26558 0 26618 1259
rect 27294 0 27354 2755
rect 34742 2752 35062 3776
rect 68540 9824 68860 9840
rect 68540 9760 68548 9824
rect 68612 9760 68628 9824
rect 68692 9760 68708 9824
rect 68772 9760 68788 9824
rect 68852 9760 68860 9824
rect 68540 8736 68860 9760
rect 69062 9621 69122 10880
rect 69798 9893 69858 10880
rect 69795 9892 69861 9893
rect 69795 9828 69796 9892
rect 69860 9828 69861 9892
rect 69795 9827 69861 9828
rect 70534 9621 70594 10880
rect 71270 10165 71330 10880
rect 72006 10437 72066 10880
rect 72003 10436 72069 10437
rect 72003 10372 72004 10436
rect 72068 10372 72069 10436
rect 72003 10371 72069 10372
rect 71267 10164 71333 10165
rect 71267 10100 71268 10164
rect 71332 10100 71333 10164
rect 71267 10099 71333 10100
rect 72742 9621 72802 10880
rect 69059 9620 69125 9621
rect 69059 9556 69060 9620
rect 69124 9556 69125 9620
rect 69059 9555 69125 9556
rect 70531 9620 70597 9621
rect 70531 9556 70532 9620
rect 70596 9556 70597 9620
rect 70531 9555 70597 9556
rect 72739 9620 72805 9621
rect 72739 9556 72740 9620
rect 72804 9556 72805 9620
rect 72739 9555 72805 9556
rect 73478 9077 73538 10880
rect 74214 9621 74274 10880
rect 74211 9620 74277 9621
rect 74211 9556 74212 9620
rect 74276 9556 74277 9620
rect 74211 9555 74277 9556
rect 74950 9077 75010 10880
rect 75686 9621 75746 10880
rect 76422 9621 76482 10880
rect 77158 9893 77218 10880
rect 77155 9892 77221 9893
rect 77155 9828 77156 9892
rect 77220 9828 77221 9892
rect 77155 9827 77221 9828
rect 77894 9621 77954 10880
rect 78630 9893 78690 10880
rect 79366 10165 79426 10880
rect 79363 10164 79429 10165
rect 79363 10100 79364 10164
rect 79428 10100 79429 10164
rect 79363 10099 79429 10100
rect 78627 9892 78693 9893
rect 78627 9828 78628 9892
rect 78692 9828 78693 9892
rect 78627 9827 78693 9828
rect 80102 9621 80162 10880
rect 80838 9893 80898 10880
rect 81574 10573 81634 10880
rect 82310 10573 82370 10880
rect 81571 10572 81637 10573
rect 81571 10508 81572 10572
rect 81636 10508 81637 10572
rect 81571 10507 81637 10508
rect 82307 10572 82373 10573
rect 82307 10508 82308 10572
rect 82372 10508 82373 10572
rect 82307 10507 82373 10508
rect 83046 10165 83106 10880
rect 83782 10165 83842 10880
rect 84518 10165 84578 10880
rect 85254 10165 85314 10880
rect 83043 10164 83109 10165
rect 83043 10100 83044 10164
rect 83108 10100 83109 10164
rect 83043 10099 83109 10100
rect 83779 10164 83845 10165
rect 83779 10100 83780 10164
rect 83844 10100 83845 10164
rect 83779 10099 83845 10100
rect 84515 10164 84581 10165
rect 84515 10100 84516 10164
rect 84580 10100 84581 10164
rect 84515 10099 84581 10100
rect 85251 10164 85317 10165
rect 85251 10100 85252 10164
rect 85316 10100 85317 10164
rect 85251 10099 85317 10100
rect 85990 9893 86050 10880
rect 86726 10573 86786 10880
rect 86723 10572 86789 10573
rect 86723 10508 86724 10572
rect 86788 10508 86789 10572
rect 86723 10507 86789 10508
rect 80835 9892 80901 9893
rect 80835 9828 80836 9892
rect 80900 9828 80901 9892
rect 80835 9827 80901 9828
rect 85987 9892 86053 9893
rect 85987 9828 85988 9892
rect 86052 9828 86053 9892
rect 85987 9827 86053 9828
rect 75683 9620 75749 9621
rect 75683 9556 75684 9620
rect 75748 9556 75749 9620
rect 75683 9555 75749 9556
rect 76419 9620 76485 9621
rect 76419 9556 76420 9620
rect 76484 9556 76485 9620
rect 76419 9555 76485 9556
rect 77891 9620 77957 9621
rect 77891 9556 77892 9620
rect 77956 9556 77957 9620
rect 77891 9555 77957 9556
rect 80099 9620 80165 9621
rect 80099 9556 80100 9620
rect 80164 9556 80165 9620
rect 80099 9555 80165 9556
rect 73475 9076 73541 9077
rect 73475 9012 73476 9076
rect 73540 9012 73541 9076
rect 73475 9011 73541 9012
rect 74947 9076 75013 9077
rect 74947 9012 74948 9076
rect 75012 9012 75013 9076
rect 74947 9011 75013 9012
rect 68540 8672 68548 8736
rect 68612 8672 68628 8736
rect 68692 8672 68708 8736
rect 68772 8672 68788 8736
rect 68852 8672 68860 8736
rect 68540 7648 68860 8672
rect 87462 8669 87522 10880
rect 88198 9213 88258 10880
rect 88195 9212 88261 9213
rect 88195 9148 88196 9212
rect 88260 9148 88261 9212
rect 88195 9147 88261 9148
rect 87459 8668 87525 8669
rect 87459 8604 87460 8668
rect 87524 8604 87525 8668
rect 87459 8603 87525 8604
rect 88934 8125 88994 10880
rect 89670 10301 89730 10880
rect 89667 10300 89733 10301
rect 89667 10236 89668 10300
rect 89732 10236 89733 10300
rect 89667 10235 89733 10236
rect 90406 8669 90466 10880
rect 91142 10029 91202 10880
rect 91139 10028 91205 10029
rect 91139 9964 91140 10028
rect 91204 9964 91205 10028
rect 91139 9963 91205 9964
rect 91878 9213 91938 10880
rect 92614 9757 92674 10880
rect 93350 9757 93410 10880
rect 92611 9756 92677 9757
rect 92611 9692 92612 9756
rect 92676 9692 92677 9756
rect 92611 9691 92677 9692
rect 93347 9756 93413 9757
rect 93347 9692 93348 9756
rect 93412 9692 93413 9756
rect 93347 9691 93413 9692
rect 91875 9212 91941 9213
rect 91875 9148 91876 9212
rect 91940 9148 91941 9212
rect 91875 9147 91941 9148
rect 94086 8669 94146 10880
rect 94822 8669 94882 10880
rect 95558 9757 95618 10880
rect 96294 9757 96354 10880
rect 96659 10436 96725 10437
rect 96659 10372 96660 10436
rect 96724 10372 96725 10436
rect 96659 10371 96725 10372
rect 95555 9756 95621 9757
rect 95555 9692 95556 9756
rect 95620 9692 95621 9756
rect 95555 9691 95621 9692
rect 96291 9756 96357 9757
rect 96291 9692 96292 9756
rect 96356 9692 96357 9756
rect 96291 9691 96357 9692
rect 96291 8940 96357 8941
rect 96291 8876 96292 8940
rect 96356 8876 96357 8940
rect 96291 8875 96357 8876
rect 90403 8668 90469 8669
rect 90403 8604 90404 8668
rect 90468 8604 90469 8668
rect 90403 8603 90469 8604
rect 94083 8668 94149 8669
rect 94083 8604 94084 8668
rect 94148 8604 94149 8668
rect 94083 8603 94149 8604
rect 94819 8668 94885 8669
rect 94819 8604 94820 8668
rect 94884 8604 94885 8668
rect 94819 8603 94885 8604
rect 88931 8124 88997 8125
rect 88931 8060 88932 8124
rect 88996 8060 88997 8124
rect 88931 8059 88997 8060
rect 68540 7584 68548 7648
rect 68612 7584 68628 7648
rect 68692 7584 68708 7648
rect 68772 7584 68788 7648
rect 68852 7584 68860 7648
rect 68540 6560 68860 7584
rect 94267 6900 94333 6901
rect 94267 6836 94268 6900
rect 94332 6836 94333 6900
rect 94267 6835 94333 6836
rect 68540 6496 68548 6560
rect 68612 6496 68628 6560
rect 68692 6496 68708 6560
rect 68772 6496 68788 6560
rect 68852 6496 68860 6560
rect 68540 5472 68860 6496
rect 93899 6356 93965 6357
rect 93899 6292 93900 6356
rect 93964 6292 93965 6356
rect 93899 6291 93965 6292
rect 68540 5408 68548 5472
rect 68612 5408 68628 5472
rect 68692 5408 68708 5472
rect 68772 5408 68788 5472
rect 68852 5408 68860 5472
rect 68540 4384 68860 5408
rect 68540 4320 68548 4384
rect 68612 4320 68628 4384
rect 68692 4320 68708 4384
rect 68772 4320 68788 4384
rect 68852 4320 68860 4384
rect 68540 3296 68860 4320
rect 68540 3232 68548 3296
rect 68612 3232 68628 3296
rect 68692 3232 68708 3296
rect 68772 3232 68788 3296
rect 68852 3232 68860 3296
rect 54891 2820 54957 2821
rect 54891 2756 54892 2820
rect 54956 2756 54957 2820
rect 54891 2755 54957 2756
rect 34742 2688 34750 2752
rect 34814 2688 34830 2752
rect 34894 2688 34910 2752
rect 34974 2688 34990 2752
rect 35054 2688 35062 2752
rect 34742 1664 35062 2688
rect 34742 1600 34750 1664
rect 34814 1600 34830 1664
rect 34894 1600 34910 1664
rect 34974 1600 34990 1664
rect 35054 1600 35062 1664
rect 32443 1596 32509 1597
rect 32443 1532 32444 1596
rect 32508 1532 32509 1596
rect 32443 1531 32509 1532
rect 29499 1188 29565 1189
rect 29499 1124 29500 1188
rect 29564 1124 29565 1188
rect 29499 1123 29565 1124
rect 28027 644 28093 645
rect 28027 580 28028 644
rect 28092 580 28093 644
rect 28027 579 28093 580
rect 28030 0 28090 579
rect 28763 372 28829 373
rect 28763 308 28764 372
rect 28828 308 28829 372
rect 28763 307 28829 308
rect 28766 0 28826 307
rect 29502 0 29562 1123
rect 30235 644 30301 645
rect 30235 580 30236 644
rect 30300 580 30301 644
rect 30235 579 30301 580
rect 30971 644 31037 645
rect 30971 580 30972 644
rect 31036 580 31037 644
rect 30971 579 31037 580
rect 31707 644 31773 645
rect 31707 580 31708 644
rect 31772 580 31773 644
rect 31707 579 31773 580
rect 30238 0 30298 579
rect 30974 0 31034 579
rect 31710 0 31770 579
rect 32446 0 32506 1531
rect 34742 1040 35062 1600
rect 34927 644 34993 645
rect 34927 580 34928 644
rect 34992 580 34993 644
rect 34927 579 34993 580
rect 35663 644 35729 645
rect 35663 580 35664 644
rect 35728 580 35729 644
rect 35663 579 35729 580
rect 36399 644 36465 645
rect 36399 580 36400 644
rect 36464 580 36465 644
rect 36399 579 36465 580
rect 37135 644 37201 645
rect 37135 580 37136 644
rect 37200 580 37201 644
rect 37135 579 37201 580
rect 37871 644 37937 645
rect 37871 580 37872 644
rect 37936 580 37937 644
rect 37871 579 37937 580
rect 38607 644 38673 645
rect 38607 580 38608 644
rect 38672 580 38673 644
rect 38607 579 38673 580
rect 40079 644 40145 645
rect 40079 580 40080 644
rect 40144 580 40145 644
rect 40079 579 40145 580
rect 40815 644 40881 645
rect 40815 580 40816 644
rect 40880 580 40881 644
rect 40815 579 40881 580
rect 41551 644 41617 645
rect 41551 580 41552 644
rect 41616 580 41617 644
rect 41551 579 41617 580
rect 42287 644 42353 645
rect 42287 580 42288 644
rect 42352 580 42353 644
rect 42287 579 42353 580
rect 43023 644 43089 645
rect 43023 580 43024 644
rect 43088 580 43089 644
rect 43023 579 43089 580
rect 43759 644 43825 645
rect 43759 580 43760 644
rect 43824 580 43825 644
rect 43759 579 43825 580
rect 44495 644 44561 645
rect 44495 580 44496 644
rect 44560 580 44561 644
rect 44495 579 44561 580
rect 45231 644 45297 645
rect 45231 580 45232 644
rect 45296 580 45297 644
rect 45231 579 45297 580
rect 45967 644 46033 645
rect 45967 580 45968 644
rect 46032 580 46033 644
rect 45967 579 46033 580
rect 46703 644 46769 645
rect 46703 580 46704 644
rect 46768 580 46769 644
rect 46703 579 46769 580
rect 47439 644 47505 645
rect 47439 580 47440 644
rect 47504 580 47505 644
rect 47439 579 47505 580
rect 48175 644 48241 645
rect 48175 580 48176 644
rect 48240 580 48241 644
rect 48175 579 48241 580
rect 48911 644 48977 645
rect 48911 580 48912 644
rect 48976 580 48977 644
rect 48911 579 48977 580
rect 49647 644 49713 645
rect 49647 580 49648 644
rect 49712 580 49713 644
rect 49647 579 49713 580
rect 50383 644 50449 645
rect 50383 580 50384 644
rect 50448 580 50449 644
rect 50383 579 50449 580
rect 51119 644 51185 645
rect 51119 580 51120 644
rect 51184 580 51185 644
rect 51119 579 51185 580
rect 51855 644 51921 645
rect 51855 580 51856 644
rect 51920 580 51921 644
rect 51855 579 51921 580
rect 53327 644 53393 645
rect 53327 580 53328 644
rect 53392 580 53393 644
rect 53327 579 53393 580
rect 54063 644 54129 645
rect 54063 580 54064 644
rect 54128 580 54129 644
rect 54063 579 54129 580
rect 34930 0 34990 579
rect 35666 0 35726 579
rect 36402 0 36462 579
rect 37138 0 37198 579
rect 37874 0 37934 579
rect 38610 0 38670 579
rect 39343 372 39409 373
rect 39343 308 39344 372
rect 39408 308 39409 372
rect 39343 307 39409 308
rect 39346 0 39406 307
rect 40082 0 40142 579
rect 40818 0 40878 579
rect 41554 0 41614 579
rect 42290 0 42350 579
rect 43026 0 43086 579
rect 43762 0 43822 579
rect 44498 0 44558 579
rect 45234 0 45294 579
rect 45970 0 46030 579
rect 46706 0 46766 579
rect 47442 0 47502 579
rect 48178 0 48238 579
rect 48914 0 48974 579
rect 49650 0 49710 579
rect 50386 0 50446 579
rect 51122 0 51182 579
rect 51858 0 51918 579
rect 52591 372 52657 373
rect 52591 308 52592 372
rect 52656 308 52657 372
rect 52591 307 52657 308
rect 52594 0 52654 307
rect 53330 0 53390 579
rect 54066 0 54126 579
rect 54894 370 54954 2755
rect 68540 2208 68860 3232
rect 93902 3229 93962 6291
rect 93899 3228 93965 3229
rect 93899 3164 93900 3228
rect 93964 3164 93965 3228
rect 93899 3163 93965 3164
rect 94083 3092 94149 3093
rect 94083 3028 94084 3092
rect 94148 3028 94149 3092
rect 94083 3027 94149 3028
rect 68540 2144 68548 2208
rect 68612 2144 68628 2208
rect 68692 2144 68708 2208
rect 68772 2144 68788 2208
rect 68852 2144 68860 2208
rect 57835 1596 57901 1597
rect 57835 1532 57836 1596
rect 57900 1532 57901 1596
rect 57835 1531 57901 1532
rect 59307 1596 59373 1597
rect 59307 1532 59308 1596
rect 59372 1532 59373 1596
rect 59307 1531 59373 1532
rect 55535 508 55601 509
rect 55535 444 55536 508
rect 55600 444 55601 508
rect 55535 443 55601 444
rect 56271 508 56337 509
rect 56271 444 56272 508
rect 56336 444 56337 508
rect 56271 443 56337 444
rect 57007 508 57073 509
rect 57007 444 57008 508
rect 57072 444 57073 508
rect 57007 443 57073 444
rect 54802 310 54954 370
rect 54802 0 54862 310
rect 55538 0 55598 443
rect 56274 0 56334 443
rect 57010 0 57070 443
rect 57838 370 57898 1531
rect 58479 508 58545 509
rect 58479 444 58480 508
rect 58544 444 58545 508
rect 58479 443 58545 444
rect 57746 310 57898 370
rect 57746 0 57806 310
rect 58482 0 58542 443
rect 59310 370 59370 1531
rect 68540 1120 68860 2144
rect 91139 1596 91205 1597
rect 91139 1532 91140 1596
rect 91204 1532 91205 1596
rect 91139 1531 91205 1532
rect 88195 1460 88261 1461
rect 88195 1396 88196 1460
rect 88260 1396 88261 1460
rect 88195 1395 88261 1396
rect 76419 1324 76485 1325
rect 76419 1260 76420 1324
rect 76484 1260 76485 1324
rect 76419 1259 76485 1260
rect 78627 1324 78693 1325
rect 78627 1260 78628 1324
rect 78692 1260 78693 1324
rect 78627 1259 78693 1260
rect 81571 1324 81637 1325
rect 81571 1260 81572 1324
rect 81636 1260 81637 1324
rect 81571 1259 81637 1260
rect 83779 1324 83845 1325
rect 83779 1260 83780 1324
rect 83844 1260 83845 1324
rect 83779 1259 83845 1260
rect 68540 1056 68548 1120
rect 68612 1056 68628 1120
rect 68692 1056 68708 1120
rect 68772 1056 68788 1120
rect 68852 1056 68860 1120
rect 68540 1040 68860 1056
rect 71267 1052 71333 1053
rect 71267 988 71268 1052
rect 71332 988 71333 1052
rect 71267 987 71333 988
rect 72003 1052 72069 1053
rect 72003 988 72004 1052
rect 72068 988 72069 1052
rect 72003 987 72069 988
rect 73475 1052 73541 1053
rect 73475 988 73476 1052
rect 73540 988 73541 1052
rect 73475 987 73541 988
rect 75683 1052 75749 1053
rect 75683 988 75684 1052
rect 75748 988 75749 1052
rect 75683 987 75749 988
rect 69059 916 69125 917
rect 69059 852 69060 916
rect 69124 852 69125 916
rect 69059 851 69125 852
rect 69795 916 69861 917
rect 69795 852 69796 916
rect 69860 852 69861 916
rect 69795 851 69861 852
rect 70531 916 70597 917
rect 70531 852 70532 916
rect 70596 852 70597 916
rect 70531 851 70597 852
rect 59951 508 60017 509
rect 59951 444 59952 508
rect 60016 444 60017 508
rect 59951 443 60017 444
rect 60687 508 60753 509
rect 60687 444 60688 508
rect 60752 444 60753 508
rect 60687 443 60753 444
rect 61423 508 61489 509
rect 61423 444 61424 508
rect 61488 444 61489 508
rect 61423 443 61489 444
rect 62159 508 62225 509
rect 62159 444 62160 508
rect 62224 444 62225 508
rect 62159 443 62225 444
rect 62895 508 62961 509
rect 62895 444 62896 508
rect 62960 444 62961 508
rect 62895 443 62961 444
rect 65839 508 65905 509
rect 65839 444 65840 508
rect 65904 444 65905 508
rect 65839 443 65905 444
rect 66575 508 66641 509
rect 66575 444 66576 508
rect 66640 444 66641 508
rect 66575 443 66641 444
rect 59218 310 59370 370
rect 59218 0 59278 310
rect 59954 0 60014 443
rect 60690 0 60750 443
rect 61426 0 61486 443
rect 62162 0 62222 443
rect 62898 0 62958 443
rect 63631 372 63697 373
rect 63631 308 63632 372
rect 63696 308 63697 372
rect 63631 307 63697 308
rect 64367 372 64433 373
rect 64367 308 64368 372
rect 64432 308 64433 372
rect 64367 307 64433 308
rect 65103 372 65169 373
rect 65103 308 65104 372
rect 65168 308 65169 372
rect 65103 307 65169 308
rect 63634 0 63694 307
rect 64370 0 64430 307
rect 65106 0 65166 307
rect 65842 0 65902 443
rect 66578 0 66638 443
rect 69062 0 69122 851
rect 69798 0 69858 851
rect 70534 0 70594 851
rect 71270 0 71330 987
rect 72006 0 72066 987
rect 72739 916 72805 917
rect 72739 852 72740 916
rect 72804 852 72805 916
rect 72739 851 72805 852
rect 72742 0 72802 851
rect 73478 0 73538 987
rect 74211 916 74277 917
rect 74211 852 74212 916
rect 74276 852 74277 916
rect 74211 851 74277 852
rect 74947 916 75013 917
rect 74947 852 74948 916
rect 75012 852 75013 916
rect 74947 851 75013 852
rect 74214 0 74274 851
rect 74950 0 75010 851
rect 75686 0 75746 987
rect 76422 0 76482 1259
rect 77155 1052 77221 1053
rect 77155 988 77156 1052
rect 77220 988 77221 1052
rect 77155 987 77221 988
rect 77158 0 77218 987
rect 77891 916 77957 917
rect 77891 852 77892 916
rect 77956 852 77957 916
rect 77891 851 77957 852
rect 77894 0 77954 851
rect 78630 0 78690 1259
rect 79363 1052 79429 1053
rect 79363 988 79364 1052
rect 79428 988 79429 1052
rect 79363 987 79429 988
rect 80835 1052 80901 1053
rect 80835 988 80836 1052
rect 80900 988 80901 1052
rect 80835 987 80901 988
rect 79366 0 79426 987
rect 80099 916 80165 917
rect 80099 852 80100 916
rect 80164 852 80165 916
rect 80099 851 80165 852
rect 80102 0 80162 851
rect 80838 0 80898 987
rect 81574 0 81634 1259
rect 82307 1052 82373 1053
rect 82307 988 82308 1052
rect 82372 988 82373 1052
rect 82307 987 82373 988
rect 82310 0 82370 987
rect 83043 916 83109 917
rect 83043 852 83044 916
rect 83108 852 83109 916
rect 83043 851 83109 852
rect 83046 0 83106 851
rect 83782 0 83842 1259
rect 84515 1052 84581 1053
rect 84515 988 84516 1052
rect 84580 988 84581 1052
rect 84515 987 84581 988
rect 85987 1052 86053 1053
rect 85987 988 85988 1052
rect 86052 988 86053 1052
rect 85987 987 86053 988
rect 84518 0 84578 987
rect 85251 372 85317 373
rect 85251 308 85252 372
rect 85316 308 85317 372
rect 85251 307 85317 308
rect 85254 0 85314 307
rect 85990 0 86050 987
rect 86723 916 86789 917
rect 86723 852 86724 916
rect 86788 852 86789 916
rect 86723 851 86789 852
rect 86726 0 86786 851
rect 87459 508 87525 509
rect 87459 444 87460 508
rect 87524 444 87525 508
rect 87459 443 87525 444
rect 87462 0 87522 443
rect 88198 0 88258 1395
rect 88931 1324 88997 1325
rect 88931 1260 88932 1324
rect 88996 1260 88997 1324
rect 88931 1259 88997 1260
rect 89851 1324 89917 1325
rect 89851 1260 89852 1324
rect 89916 1260 89917 1324
rect 89851 1259 89917 1260
rect 90403 1324 90469 1325
rect 90403 1260 90404 1324
rect 90468 1260 90469 1324
rect 90403 1259 90469 1260
rect 88934 0 88994 1259
rect 89854 370 89914 1259
rect 89670 310 89914 370
rect 89670 0 89730 310
rect 90406 0 90466 1259
rect 91142 0 91202 1531
rect 91875 1324 91941 1325
rect 91875 1260 91876 1324
rect 91940 1260 91941 1324
rect 91875 1259 91941 1260
rect 93347 1324 93413 1325
rect 93347 1260 93348 1324
rect 93412 1260 93413 1324
rect 93347 1259 93413 1260
rect 91878 0 91938 1259
rect 92611 644 92677 645
rect 92611 580 92612 644
rect 92676 580 92677 644
rect 92611 579 92677 580
rect 92614 0 92674 579
rect 93350 0 93410 1259
rect 94086 0 94146 3027
rect 94270 2141 94330 6835
rect 95187 5540 95253 5541
rect 95187 5476 95188 5540
rect 95252 5476 95253 5540
rect 95187 5475 95253 5476
rect 94267 2140 94333 2141
rect 94267 2076 94268 2140
rect 94332 2076 94333 2140
rect 94267 2075 94333 2076
rect 94819 644 94885 645
rect 94819 580 94820 644
rect 94884 580 94885 644
rect 94819 579 94885 580
rect 94822 0 94882 579
rect 95190 373 95250 5475
rect 96294 3229 96354 8875
rect 96475 4180 96541 4181
rect 96475 4116 96476 4180
rect 96540 4116 96541 4180
rect 96475 4115 96541 4116
rect 96291 3228 96357 3229
rect 96291 3164 96292 3228
rect 96356 3164 96357 3228
rect 96291 3163 96357 3164
rect 95555 2820 95621 2821
rect 95555 2756 95556 2820
rect 95620 2756 95621 2820
rect 95555 2755 95621 2756
rect 95187 372 95253 373
rect 95187 308 95188 372
rect 95252 308 95253 372
rect 95187 307 95253 308
rect 95558 0 95618 2755
rect 96478 2141 96538 4115
rect 96662 2413 96722 10371
rect 97030 8669 97090 10880
rect 97766 8669 97826 10880
rect 98502 9757 98562 10880
rect 98499 9756 98565 9757
rect 98499 9692 98500 9756
rect 98564 9692 98565 9756
rect 98499 9691 98565 9692
rect 99238 8669 99298 10880
rect 99974 9757 100034 10880
rect 99971 9756 100037 9757
rect 99971 9692 99972 9756
rect 100036 9692 100037 9756
rect 99971 9691 100037 9692
rect 100710 9213 100770 10880
rect 103194 10301 103254 10880
rect 103930 10301 103990 10880
rect 104666 10301 104726 10880
rect 105402 10301 105462 10880
rect 106138 10301 106198 10880
rect 106874 10301 106934 10880
rect 107610 10301 107670 10880
rect 108346 10301 108406 10880
rect 109082 10301 109142 10880
rect 109818 10301 109878 10880
rect 110554 10301 110614 10880
rect 111290 10301 111350 10880
rect 112026 10301 112086 10880
rect 112762 10301 112822 10880
rect 113498 10301 113558 10880
rect 114234 10301 114294 10880
rect 114970 10301 115030 10880
rect 115706 10301 115766 10880
rect 116442 10301 116502 10880
rect 117178 10301 117238 10880
rect 117914 10301 117974 10880
rect 118650 10301 118710 10880
rect 119386 10301 119446 10880
rect 120122 10301 120182 10880
rect 120858 10301 120918 10880
rect 121594 10301 121654 10880
rect 122330 10301 122390 10880
rect 123066 10301 123126 10880
rect 123802 10301 123862 10880
rect 124538 10301 124598 10880
rect 125274 10437 125334 10880
rect 125271 10436 125337 10437
rect 125271 10372 125272 10436
rect 125336 10372 125337 10436
rect 125271 10371 125337 10372
rect 126010 10301 126070 10880
rect 126746 10301 126806 10880
rect 127482 10301 127542 10880
rect 128218 10301 128278 10880
rect 128954 10301 129014 10880
rect 129690 10301 129750 10880
rect 130426 10301 130486 10880
rect 131162 10301 131222 10880
rect 131898 10301 131958 10880
rect 132634 10301 132694 10880
rect 133370 10301 133430 10880
rect 134106 10301 134166 10880
rect 134842 10301 134902 10880
rect 103191 10300 103257 10301
rect 103191 10236 103192 10300
rect 103256 10236 103257 10300
rect 103191 10235 103257 10236
rect 103927 10300 103993 10301
rect 103927 10236 103928 10300
rect 103992 10236 103993 10300
rect 103927 10235 103993 10236
rect 104663 10300 104729 10301
rect 104663 10236 104664 10300
rect 104728 10236 104729 10300
rect 104663 10235 104729 10236
rect 105399 10300 105465 10301
rect 105399 10236 105400 10300
rect 105464 10236 105465 10300
rect 105399 10235 105465 10236
rect 106135 10300 106201 10301
rect 106135 10236 106136 10300
rect 106200 10236 106201 10300
rect 106135 10235 106201 10236
rect 106871 10300 106937 10301
rect 106871 10236 106872 10300
rect 106936 10236 106937 10300
rect 106871 10235 106937 10236
rect 107607 10300 107673 10301
rect 107607 10236 107608 10300
rect 107672 10236 107673 10300
rect 107607 10235 107673 10236
rect 108343 10300 108409 10301
rect 108343 10236 108344 10300
rect 108408 10236 108409 10300
rect 108343 10235 108409 10236
rect 109079 10300 109145 10301
rect 109079 10236 109080 10300
rect 109144 10236 109145 10300
rect 109079 10235 109145 10236
rect 109815 10300 109881 10301
rect 109815 10236 109816 10300
rect 109880 10236 109881 10300
rect 109815 10235 109881 10236
rect 110551 10300 110617 10301
rect 110551 10236 110552 10300
rect 110616 10236 110617 10300
rect 110551 10235 110617 10236
rect 111287 10300 111353 10301
rect 111287 10236 111288 10300
rect 111352 10236 111353 10300
rect 111287 10235 111353 10236
rect 112023 10300 112089 10301
rect 112023 10236 112024 10300
rect 112088 10236 112089 10300
rect 112023 10235 112089 10236
rect 112759 10300 112825 10301
rect 112759 10236 112760 10300
rect 112824 10236 112825 10300
rect 112759 10235 112825 10236
rect 113495 10300 113561 10301
rect 113495 10236 113496 10300
rect 113560 10236 113561 10300
rect 113495 10235 113561 10236
rect 114231 10300 114297 10301
rect 114231 10236 114232 10300
rect 114296 10236 114297 10300
rect 114231 10235 114297 10236
rect 114967 10300 115033 10301
rect 114967 10236 114968 10300
rect 115032 10236 115033 10300
rect 114967 10235 115033 10236
rect 115703 10300 115769 10301
rect 115703 10236 115704 10300
rect 115768 10236 115769 10300
rect 115703 10235 115769 10236
rect 116439 10300 116505 10301
rect 116439 10236 116440 10300
rect 116504 10236 116505 10300
rect 116439 10235 116505 10236
rect 117175 10300 117241 10301
rect 117175 10236 117176 10300
rect 117240 10236 117241 10300
rect 117175 10235 117241 10236
rect 117911 10300 117977 10301
rect 117911 10236 117912 10300
rect 117976 10236 117977 10300
rect 117911 10235 117977 10236
rect 118647 10300 118713 10301
rect 118647 10236 118648 10300
rect 118712 10236 118713 10300
rect 118647 10235 118713 10236
rect 119383 10300 119449 10301
rect 119383 10236 119384 10300
rect 119448 10236 119449 10300
rect 119383 10235 119449 10236
rect 120119 10300 120185 10301
rect 120119 10236 120120 10300
rect 120184 10236 120185 10300
rect 120119 10235 120185 10236
rect 120855 10300 120921 10301
rect 120855 10236 120856 10300
rect 120920 10236 120921 10300
rect 120855 10235 120921 10236
rect 121591 10300 121657 10301
rect 121591 10236 121592 10300
rect 121656 10236 121657 10300
rect 121591 10235 121657 10236
rect 122327 10300 122393 10301
rect 122327 10236 122328 10300
rect 122392 10236 122393 10300
rect 122327 10235 122393 10236
rect 123063 10300 123129 10301
rect 123063 10236 123064 10300
rect 123128 10236 123129 10300
rect 123063 10235 123129 10236
rect 123799 10300 123865 10301
rect 123799 10236 123800 10300
rect 123864 10236 123865 10300
rect 123799 10235 123865 10236
rect 124535 10300 124601 10301
rect 124535 10236 124536 10300
rect 124600 10236 124601 10300
rect 124535 10235 124601 10236
rect 126007 10300 126073 10301
rect 126007 10236 126008 10300
rect 126072 10236 126073 10300
rect 126007 10235 126073 10236
rect 126743 10300 126809 10301
rect 126743 10236 126744 10300
rect 126808 10236 126809 10300
rect 126743 10235 126809 10236
rect 127479 10300 127545 10301
rect 127479 10236 127480 10300
rect 127544 10236 127545 10300
rect 127479 10235 127545 10236
rect 128215 10300 128281 10301
rect 128215 10236 128216 10300
rect 128280 10236 128281 10300
rect 128215 10235 128281 10236
rect 128951 10300 129017 10301
rect 128951 10236 128952 10300
rect 129016 10236 129017 10300
rect 128951 10235 129017 10236
rect 129687 10300 129753 10301
rect 129687 10236 129688 10300
rect 129752 10236 129753 10300
rect 129687 10235 129753 10236
rect 130423 10300 130489 10301
rect 130423 10236 130424 10300
rect 130488 10236 130489 10300
rect 130423 10235 130489 10236
rect 131159 10300 131225 10301
rect 131159 10236 131160 10300
rect 131224 10236 131225 10300
rect 131159 10235 131225 10236
rect 131895 10300 131961 10301
rect 131895 10236 131896 10300
rect 131960 10236 131961 10300
rect 131895 10235 131961 10236
rect 132631 10300 132697 10301
rect 132631 10236 132632 10300
rect 132696 10236 132697 10300
rect 132631 10235 132697 10236
rect 133367 10300 133433 10301
rect 133367 10236 133368 10300
rect 133432 10236 133433 10300
rect 133367 10235 133433 10236
rect 134103 10300 134169 10301
rect 134103 10236 134104 10300
rect 134168 10236 134169 10300
rect 134103 10235 134169 10236
rect 134839 10300 134905 10301
rect 134839 10236 134840 10300
rect 134904 10236 134905 10300
rect 134839 10235 134905 10236
rect 102339 9280 102659 9840
rect 102339 9216 102347 9280
rect 102411 9216 102427 9280
rect 102491 9216 102507 9280
rect 102571 9216 102587 9280
rect 102651 9216 102659 9280
rect 100707 9212 100773 9213
rect 100707 9148 100708 9212
rect 100772 9148 100773 9212
rect 100707 9147 100773 9148
rect 97027 8668 97093 8669
rect 97027 8604 97028 8668
rect 97092 8604 97093 8668
rect 97027 8603 97093 8604
rect 97763 8668 97829 8669
rect 97763 8604 97764 8668
rect 97828 8604 97829 8668
rect 97763 8603 97829 8604
rect 99235 8668 99301 8669
rect 99235 8604 99236 8668
rect 99300 8604 99301 8668
rect 99235 8603 99301 8604
rect 102339 8192 102659 9216
rect 102339 8128 102347 8192
rect 102411 8128 102427 8192
rect 102491 8128 102507 8192
rect 102571 8128 102587 8192
rect 102651 8128 102659 8192
rect 96843 8124 96909 8125
rect 96843 8060 96844 8124
rect 96908 8060 96909 8124
rect 96843 8059 96909 8060
rect 96846 3229 96906 8059
rect 102339 7104 102659 8128
rect 102339 7040 102347 7104
rect 102411 7040 102427 7104
rect 102491 7040 102507 7104
rect 102571 7040 102587 7104
rect 102651 7040 102659 7104
rect 102339 6016 102659 7040
rect 136137 9824 136457 9840
rect 136137 9760 136145 9824
rect 136209 9760 136225 9824
rect 136289 9760 136305 9824
rect 136369 9760 136385 9824
rect 136449 9760 136457 9824
rect 136137 8736 136457 9760
rect 137326 9621 137386 10880
rect 138062 10301 138122 10880
rect 138059 10300 138125 10301
rect 138059 10236 138060 10300
rect 138124 10236 138125 10300
rect 138059 10235 138125 10236
rect 138798 10165 138858 10880
rect 138795 10164 138861 10165
rect 138795 10100 138796 10164
rect 138860 10100 138861 10164
rect 138795 10099 138861 10100
rect 139534 9893 139594 10880
rect 140270 10165 140330 10880
rect 141006 10165 141066 10880
rect 141742 10165 141802 10880
rect 142478 10301 142538 10880
rect 142475 10300 142541 10301
rect 142475 10236 142476 10300
rect 142540 10236 142541 10300
rect 142475 10235 142541 10236
rect 143214 10165 143274 10880
rect 143950 10165 144010 10880
rect 140267 10164 140333 10165
rect 140267 10100 140268 10164
rect 140332 10100 140333 10164
rect 140267 10099 140333 10100
rect 141003 10164 141069 10165
rect 141003 10100 141004 10164
rect 141068 10100 141069 10164
rect 141003 10099 141069 10100
rect 141739 10164 141805 10165
rect 141739 10100 141740 10164
rect 141804 10100 141805 10164
rect 141739 10099 141805 10100
rect 143211 10164 143277 10165
rect 143211 10100 143212 10164
rect 143276 10100 143277 10164
rect 143211 10099 143277 10100
rect 143947 10164 144013 10165
rect 143947 10100 143948 10164
rect 144012 10100 144013 10164
rect 143947 10099 144013 10100
rect 144686 9893 144746 10880
rect 145422 10165 145482 10880
rect 146158 10165 146218 10880
rect 146894 10165 146954 10880
rect 147630 10573 147690 10880
rect 147627 10572 147693 10573
rect 147627 10508 147628 10572
rect 147692 10508 147693 10572
rect 147627 10507 147693 10508
rect 148366 10301 148426 10880
rect 148363 10300 148429 10301
rect 148363 10236 148364 10300
rect 148428 10236 148429 10300
rect 148363 10235 148429 10236
rect 149102 10165 149162 10880
rect 145419 10164 145485 10165
rect 145419 10100 145420 10164
rect 145484 10100 145485 10164
rect 145419 10099 145485 10100
rect 146155 10164 146221 10165
rect 146155 10100 146156 10164
rect 146220 10100 146221 10164
rect 146155 10099 146221 10100
rect 146891 10164 146957 10165
rect 146891 10100 146892 10164
rect 146956 10100 146957 10164
rect 146891 10099 146957 10100
rect 149099 10164 149165 10165
rect 149099 10100 149100 10164
rect 149164 10100 149165 10164
rect 149099 10099 149165 10100
rect 149838 9893 149898 10880
rect 150574 10165 150634 10880
rect 151310 10165 151370 10880
rect 152046 10165 152106 10880
rect 152782 10165 152842 10880
rect 153518 10165 153578 10880
rect 154254 10437 154314 10880
rect 154251 10436 154317 10437
rect 154251 10372 154252 10436
rect 154316 10372 154317 10436
rect 154251 10371 154317 10372
rect 150571 10164 150637 10165
rect 150571 10100 150572 10164
rect 150636 10100 150637 10164
rect 150571 10099 150637 10100
rect 151307 10164 151373 10165
rect 151307 10100 151308 10164
rect 151372 10100 151373 10164
rect 151307 10099 151373 10100
rect 152043 10164 152109 10165
rect 152043 10100 152044 10164
rect 152108 10100 152109 10164
rect 152043 10099 152109 10100
rect 152779 10164 152845 10165
rect 152779 10100 152780 10164
rect 152844 10100 152845 10164
rect 152779 10099 152845 10100
rect 153515 10164 153581 10165
rect 153515 10100 153516 10164
rect 153580 10100 153581 10164
rect 153515 10099 153581 10100
rect 154990 9893 155050 10880
rect 139531 9892 139597 9893
rect 139531 9828 139532 9892
rect 139596 9828 139597 9892
rect 139531 9827 139597 9828
rect 144683 9892 144749 9893
rect 144683 9828 144684 9892
rect 144748 9828 144749 9892
rect 144683 9827 144749 9828
rect 149835 9892 149901 9893
rect 149835 9828 149836 9892
rect 149900 9828 149901 9892
rect 149835 9827 149901 9828
rect 154987 9892 155053 9893
rect 154987 9828 154988 9892
rect 155052 9828 155053 9892
rect 154987 9827 155053 9828
rect 137323 9620 137389 9621
rect 137323 9556 137324 9620
rect 137388 9556 137389 9620
rect 137323 9555 137389 9556
rect 136137 8672 136145 8736
rect 136209 8672 136225 8736
rect 136289 8672 136305 8736
rect 136369 8672 136385 8736
rect 136449 8672 136457 8736
rect 136137 7648 136457 8672
rect 155726 8669 155786 10880
rect 156462 9485 156522 10880
rect 156459 9484 156525 9485
rect 156459 9420 156460 9484
rect 156524 9420 156525 9484
rect 156459 9419 156525 9420
rect 155723 8668 155789 8669
rect 155723 8604 155724 8668
rect 155788 8604 155789 8668
rect 155723 8603 155789 8604
rect 157198 8397 157258 10880
rect 157195 8396 157261 8397
rect 157195 8332 157196 8396
rect 157260 8332 157261 8396
rect 157195 8331 157261 8332
rect 157934 8125 157994 10880
rect 158670 8397 158730 10880
rect 158667 8396 158733 8397
rect 158667 8332 158668 8396
rect 158732 8332 158733 8396
rect 158667 8331 158733 8332
rect 159406 8125 159466 10880
rect 160142 8397 160202 10880
rect 160139 8396 160205 8397
rect 160139 8332 160140 8396
rect 160204 8332 160205 8396
rect 160139 8331 160205 8332
rect 160878 8125 160938 10880
rect 161614 8397 161674 10880
rect 161611 8396 161677 8397
rect 161611 8332 161612 8396
rect 161676 8332 161677 8396
rect 161611 8331 161677 8332
rect 157931 8124 157997 8125
rect 157931 8060 157932 8124
rect 157996 8060 157997 8124
rect 157931 8059 157997 8060
rect 159403 8124 159469 8125
rect 159403 8060 159404 8124
rect 159468 8060 159469 8124
rect 159403 8059 159469 8060
rect 160875 8124 160941 8125
rect 160875 8060 160876 8124
rect 160940 8060 160941 8124
rect 160875 8059 160941 8060
rect 162350 7853 162410 10880
rect 163086 8397 163146 10880
rect 163083 8396 163149 8397
rect 163083 8332 163084 8396
rect 163148 8332 163149 8396
rect 163083 8331 163149 8332
rect 163822 8125 163882 10880
rect 164558 8397 164618 10880
rect 164555 8396 164621 8397
rect 164555 8332 164556 8396
rect 164620 8332 164621 8396
rect 164555 8331 164621 8332
rect 165294 8125 165354 10880
rect 166030 8397 166090 10880
rect 166766 8397 166826 10880
rect 167502 9757 167562 10880
rect 167499 9756 167565 9757
rect 167499 9692 167500 9756
rect 167564 9692 167565 9756
rect 167499 9691 167565 9692
rect 168238 9213 168298 10880
rect 168974 9757 169034 10880
rect 171458 10301 171518 10880
rect 172194 10573 172254 10880
rect 172191 10572 172257 10573
rect 172191 10508 172192 10572
rect 172256 10508 172257 10572
rect 172191 10507 172257 10508
rect 172930 10437 172990 10880
rect 172927 10436 172993 10437
rect 172927 10372 172928 10436
rect 172992 10372 172993 10436
rect 172927 10371 172993 10372
rect 173666 10301 173726 10880
rect 174402 10301 174462 10880
rect 175138 10301 175198 10880
rect 175874 10301 175934 10880
rect 176610 10301 176670 10880
rect 177346 10301 177406 10880
rect 178082 10301 178142 10880
rect 178818 10301 178878 10880
rect 179554 10573 179614 10880
rect 179551 10572 179617 10573
rect 179551 10508 179552 10572
rect 179616 10508 179617 10572
rect 179551 10507 179617 10508
rect 180290 10301 180350 10880
rect 181026 10437 181086 10880
rect 181023 10436 181089 10437
rect 181023 10372 181024 10436
rect 181088 10372 181089 10436
rect 181023 10371 181089 10372
rect 181762 10301 181822 10880
rect 182498 10301 182558 10880
rect 183234 10301 183294 10880
rect 183970 10301 184030 10880
rect 184706 10301 184766 10880
rect 185442 10301 185502 10880
rect 186178 10301 186238 10880
rect 186914 10301 186974 10880
rect 187650 10301 187710 10880
rect 188386 10301 188446 10880
rect 189122 10301 189182 10880
rect 189858 10301 189918 10880
rect 190594 10437 190654 10880
rect 190591 10436 190657 10437
rect 190591 10372 190592 10436
rect 190656 10372 190657 10436
rect 190591 10371 190657 10372
rect 191330 10301 191390 10880
rect 192066 10301 192126 10880
rect 192802 10437 192862 10880
rect 192799 10436 192865 10437
rect 192799 10372 192800 10436
rect 192864 10372 192865 10436
rect 192799 10371 192865 10372
rect 193538 10301 193598 10880
rect 194274 10301 194334 10880
rect 195010 10301 195070 10880
rect 195746 10301 195806 10880
rect 196482 10301 196542 10880
rect 197218 10301 197278 10880
rect 197954 10301 198014 10880
rect 198690 10301 198750 10880
rect 199426 10301 199486 10880
rect 200162 10301 200222 10880
rect 200898 10301 200958 10880
rect 201634 10301 201694 10880
rect 202370 10437 202430 10880
rect 202367 10436 202433 10437
rect 202367 10372 202368 10436
rect 202432 10372 202433 10436
rect 202367 10371 202433 10372
rect 203106 10301 203166 10880
rect 205590 10301 205650 10880
rect 171455 10300 171521 10301
rect 171455 10236 171456 10300
rect 171520 10236 171521 10300
rect 171455 10235 171521 10236
rect 173663 10300 173729 10301
rect 173663 10236 173664 10300
rect 173728 10236 173729 10300
rect 173663 10235 173729 10236
rect 174399 10300 174465 10301
rect 174399 10236 174400 10300
rect 174464 10236 174465 10300
rect 174399 10235 174465 10236
rect 175135 10300 175201 10301
rect 175135 10236 175136 10300
rect 175200 10236 175201 10300
rect 175135 10235 175201 10236
rect 175871 10300 175937 10301
rect 175871 10236 175872 10300
rect 175936 10236 175937 10300
rect 175871 10235 175937 10236
rect 176607 10300 176673 10301
rect 176607 10236 176608 10300
rect 176672 10236 176673 10300
rect 176607 10235 176673 10236
rect 177343 10300 177409 10301
rect 177343 10236 177344 10300
rect 177408 10236 177409 10300
rect 177343 10235 177409 10236
rect 178079 10300 178145 10301
rect 178079 10236 178080 10300
rect 178144 10236 178145 10300
rect 178079 10235 178145 10236
rect 178815 10300 178881 10301
rect 178815 10236 178816 10300
rect 178880 10236 178881 10300
rect 178815 10235 178881 10236
rect 180287 10300 180353 10301
rect 180287 10236 180288 10300
rect 180352 10236 180353 10300
rect 180287 10235 180353 10236
rect 181759 10300 181825 10301
rect 181759 10236 181760 10300
rect 181824 10236 181825 10300
rect 181759 10235 181825 10236
rect 182495 10300 182561 10301
rect 182495 10236 182496 10300
rect 182560 10236 182561 10300
rect 182495 10235 182561 10236
rect 183231 10300 183297 10301
rect 183231 10236 183232 10300
rect 183296 10236 183297 10300
rect 183231 10235 183297 10236
rect 183967 10300 184033 10301
rect 183967 10236 183968 10300
rect 184032 10236 184033 10300
rect 183967 10235 184033 10236
rect 184703 10300 184769 10301
rect 184703 10236 184704 10300
rect 184768 10236 184769 10300
rect 184703 10235 184769 10236
rect 185439 10300 185505 10301
rect 185439 10236 185440 10300
rect 185504 10236 185505 10300
rect 185439 10235 185505 10236
rect 186175 10300 186241 10301
rect 186175 10236 186176 10300
rect 186240 10236 186241 10300
rect 186175 10235 186241 10236
rect 186911 10300 186977 10301
rect 186911 10236 186912 10300
rect 186976 10236 186977 10300
rect 186911 10235 186977 10236
rect 187647 10300 187713 10301
rect 187647 10236 187648 10300
rect 187712 10236 187713 10300
rect 187647 10235 187713 10236
rect 188383 10300 188449 10301
rect 188383 10236 188384 10300
rect 188448 10236 188449 10300
rect 188383 10235 188449 10236
rect 189119 10300 189185 10301
rect 189119 10236 189120 10300
rect 189184 10236 189185 10300
rect 189119 10235 189185 10236
rect 189855 10300 189921 10301
rect 189855 10236 189856 10300
rect 189920 10236 189921 10300
rect 189855 10235 189921 10236
rect 191327 10300 191393 10301
rect 191327 10236 191328 10300
rect 191392 10236 191393 10300
rect 191327 10235 191393 10236
rect 192063 10300 192129 10301
rect 192063 10236 192064 10300
rect 192128 10236 192129 10300
rect 192063 10235 192129 10236
rect 193535 10300 193601 10301
rect 193535 10236 193536 10300
rect 193600 10236 193601 10300
rect 193535 10235 193601 10236
rect 194271 10300 194337 10301
rect 194271 10236 194272 10300
rect 194336 10236 194337 10300
rect 194271 10235 194337 10236
rect 195007 10300 195073 10301
rect 195007 10236 195008 10300
rect 195072 10236 195073 10300
rect 195007 10235 195073 10236
rect 195743 10300 195809 10301
rect 195743 10236 195744 10300
rect 195808 10236 195809 10300
rect 195743 10235 195809 10236
rect 196479 10300 196545 10301
rect 196479 10236 196480 10300
rect 196544 10236 196545 10300
rect 196479 10235 196545 10236
rect 197215 10300 197281 10301
rect 197215 10236 197216 10300
rect 197280 10236 197281 10300
rect 197215 10235 197281 10236
rect 197951 10300 198017 10301
rect 197951 10236 197952 10300
rect 198016 10236 198017 10300
rect 197951 10235 198017 10236
rect 198687 10300 198753 10301
rect 198687 10236 198688 10300
rect 198752 10236 198753 10300
rect 198687 10235 198753 10236
rect 199423 10300 199489 10301
rect 199423 10236 199424 10300
rect 199488 10236 199489 10300
rect 199423 10235 199489 10236
rect 200159 10300 200225 10301
rect 200159 10236 200160 10300
rect 200224 10236 200225 10300
rect 200159 10235 200225 10236
rect 200895 10300 200961 10301
rect 200895 10236 200896 10300
rect 200960 10236 200961 10300
rect 200895 10235 200961 10236
rect 201631 10300 201697 10301
rect 201631 10236 201632 10300
rect 201696 10236 201697 10300
rect 201631 10235 201697 10236
rect 203103 10300 203169 10301
rect 203103 10236 203104 10300
rect 203168 10236 203169 10300
rect 203103 10235 203169 10236
rect 205587 10300 205653 10301
rect 205587 10236 205588 10300
rect 205652 10236 205653 10300
rect 205587 10235 205653 10236
rect 206326 10165 206386 10880
rect 207062 10165 207122 10880
rect 207798 10573 207858 10880
rect 207795 10572 207861 10573
rect 207795 10508 207796 10572
rect 207860 10508 207861 10572
rect 207795 10507 207861 10508
rect 208534 10165 208594 10880
rect 209270 10165 209330 10880
rect 210006 10437 210066 10880
rect 210003 10436 210069 10437
rect 210003 10372 210004 10436
rect 210068 10372 210069 10436
rect 210003 10371 210069 10372
rect 210742 10165 210802 10880
rect 206323 10164 206389 10165
rect 206323 10100 206324 10164
rect 206388 10100 206389 10164
rect 206323 10099 206389 10100
rect 207059 10164 207125 10165
rect 207059 10100 207060 10164
rect 207124 10100 207125 10164
rect 207059 10099 207125 10100
rect 208531 10164 208597 10165
rect 208531 10100 208532 10164
rect 208596 10100 208597 10164
rect 208531 10099 208597 10100
rect 209267 10164 209333 10165
rect 209267 10100 209268 10164
rect 209332 10100 209333 10164
rect 209267 10099 209333 10100
rect 210739 10164 210805 10165
rect 210739 10100 210740 10164
rect 210804 10100 210805 10164
rect 210739 10099 210805 10100
rect 211478 9893 211538 10880
rect 212214 10165 212274 10880
rect 212950 10573 213010 10880
rect 212947 10572 213013 10573
rect 212947 10508 212948 10572
rect 213012 10508 213013 10572
rect 212947 10507 213013 10508
rect 213686 10165 213746 10880
rect 214422 10165 214482 10880
rect 212211 10164 212277 10165
rect 212211 10100 212212 10164
rect 212276 10100 212277 10164
rect 212211 10099 212277 10100
rect 213683 10164 213749 10165
rect 213683 10100 213684 10164
rect 213748 10100 213749 10164
rect 213683 10099 213749 10100
rect 214419 10164 214485 10165
rect 214419 10100 214420 10164
rect 214484 10100 214485 10164
rect 214419 10099 214485 10100
rect 211475 9892 211541 9893
rect 168971 9756 169037 9757
rect 168971 9692 168972 9756
rect 169036 9692 169037 9756
rect 168971 9691 169037 9692
rect 169936 9280 170256 9840
rect 169936 9216 169944 9280
rect 170008 9216 170024 9280
rect 170088 9216 170104 9280
rect 170168 9216 170184 9280
rect 170248 9216 170256 9280
rect 168235 9212 168301 9213
rect 168235 9148 168236 9212
rect 168300 9148 168301 9212
rect 168235 9147 168301 9148
rect 166027 8396 166093 8397
rect 166027 8332 166028 8396
rect 166092 8332 166093 8396
rect 166027 8331 166093 8332
rect 166763 8396 166829 8397
rect 166763 8332 166764 8396
rect 166828 8332 166829 8396
rect 166763 8331 166829 8332
rect 169936 8192 170256 9216
rect 169936 8128 169944 8192
rect 170008 8128 170024 8192
rect 170088 8128 170104 8192
rect 170168 8128 170184 8192
rect 170248 8128 170256 8192
rect 163819 8124 163885 8125
rect 163819 8060 163820 8124
rect 163884 8060 163885 8124
rect 163819 8059 163885 8060
rect 165291 8124 165357 8125
rect 165291 8060 165292 8124
rect 165356 8060 165357 8124
rect 165291 8059 165357 8060
rect 162347 7852 162413 7853
rect 162347 7788 162348 7852
rect 162412 7788 162413 7852
rect 162347 7787 162413 7788
rect 136137 7584 136145 7648
rect 136209 7584 136225 7648
rect 136289 7584 136305 7648
rect 136369 7584 136385 7648
rect 136449 7584 136457 7648
rect 107147 6900 107213 6901
rect 107147 6836 107148 6900
rect 107212 6836 107213 6900
rect 107147 6835 107213 6836
rect 102339 5952 102347 6016
rect 102411 5952 102427 6016
rect 102491 5952 102507 6016
rect 102571 5952 102587 6016
rect 102651 5952 102659 6016
rect 102339 4928 102659 5952
rect 102339 4864 102347 4928
rect 102411 4864 102427 4928
rect 102491 4864 102507 4928
rect 102571 4864 102587 4928
rect 102651 4864 102659 4928
rect 102339 3840 102659 4864
rect 106043 4860 106109 4861
rect 106043 4796 106044 4860
rect 106108 4796 106109 4860
rect 106043 4795 106109 4796
rect 103283 4044 103349 4045
rect 103283 3980 103284 4044
rect 103348 3980 103349 4044
rect 103283 3979 103349 3980
rect 104571 4044 104637 4045
rect 104571 3980 104572 4044
rect 104636 3980 104637 4044
rect 104571 3979 104637 3980
rect 105491 4044 105557 4045
rect 105491 3980 105492 4044
rect 105556 3980 105557 4044
rect 105491 3979 105557 3980
rect 102339 3776 102347 3840
rect 102411 3776 102427 3840
rect 102491 3776 102507 3840
rect 102571 3776 102587 3840
rect 102651 3776 102659 3840
rect 97763 3772 97829 3773
rect 97763 3708 97764 3772
rect 97828 3708 97829 3772
rect 97763 3707 97829 3708
rect 96843 3228 96909 3229
rect 96843 3164 96844 3228
rect 96908 3164 96909 3228
rect 96843 3163 96909 3164
rect 97027 2820 97093 2821
rect 97027 2756 97028 2820
rect 97092 2756 97093 2820
rect 97027 2755 97093 2756
rect 96659 2412 96725 2413
rect 96659 2348 96660 2412
rect 96724 2348 96725 2412
rect 96659 2347 96725 2348
rect 96475 2140 96541 2141
rect 96475 2076 96476 2140
rect 96540 2076 96541 2140
rect 96475 2075 96541 2076
rect 96291 1596 96357 1597
rect 96291 1532 96292 1596
rect 96356 1532 96357 1596
rect 96291 1531 96357 1532
rect 96294 0 96354 1531
rect 97030 0 97090 2755
rect 97766 0 97826 3707
rect 100707 3228 100773 3229
rect 100707 3164 100708 3228
rect 100772 3164 100773 3228
rect 100707 3163 100773 3164
rect 98499 1596 98565 1597
rect 98499 1532 98500 1596
rect 98564 1532 98565 1596
rect 98499 1531 98565 1532
rect 98502 0 98562 1531
rect 99235 916 99301 917
rect 99235 852 99236 916
rect 99300 852 99301 916
rect 99235 851 99301 852
rect 99238 0 99298 851
rect 99971 644 100037 645
rect 99971 580 99972 644
rect 100036 580 100037 644
rect 99971 579 100037 580
rect 99974 0 100034 579
rect 100710 0 100770 3163
rect 102339 2752 102659 3776
rect 102339 2688 102347 2752
rect 102411 2688 102427 2752
rect 102491 2688 102507 2752
rect 102571 2688 102587 2752
rect 102651 2688 102659 2752
rect 102339 1664 102659 2688
rect 102339 1600 102347 1664
rect 102411 1600 102427 1664
rect 102491 1600 102507 1664
rect 102571 1600 102587 1664
rect 102651 1600 102659 1664
rect 102339 1040 102659 1600
rect 103286 370 103346 3979
rect 104019 3908 104085 3909
rect 104019 3844 104020 3908
rect 104084 3844 104085 3908
rect 104019 3843 104085 3844
rect 104022 370 104082 3843
rect 103194 310 103346 370
rect 103930 310 104082 370
rect 104574 370 104634 3979
rect 105494 370 105554 3979
rect 104574 310 104726 370
rect 103194 0 103254 310
rect 103930 0 103990 310
rect 104666 0 104726 310
rect 105402 310 105554 370
rect 106046 370 106106 4795
rect 106963 4044 107029 4045
rect 106963 3980 106964 4044
rect 107028 3980 107029 4044
rect 106963 3979 107029 3980
rect 106966 370 107026 3979
rect 107150 3773 107210 6835
rect 136137 6560 136457 7584
rect 169936 7104 170256 8128
rect 169936 7040 169944 7104
rect 170008 7040 170024 7104
rect 170088 7040 170104 7104
rect 170168 7040 170184 7104
rect 170248 7040 170256 7104
rect 151675 6628 151741 6629
rect 151675 6564 151676 6628
rect 151740 6564 151741 6628
rect 151675 6563 151741 6564
rect 136137 6496 136145 6560
rect 136209 6496 136225 6560
rect 136289 6496 136305 6560
rect 136369 6496 136385 6560
rect 136449 6496 136457 6560
rect 136137 5472 136457 6496
rect 136137 5408 136145 5472
rect 136209 5408 136225 5472
rect 136289 5408 136305 5472
rect 136369 5408 136385 5472
rect 136449 5408 136457 5472
rect 113035 5404 113101 5405
rect 113035 5340 113036 5404
rect 113100 5340 113101 5404
rect 113035 5339 113101 5340
rect 110275 4860 110341 4861
rect 110275 4796 110276 4860
rect 110340 4796 110341 4860
rect 110275 4795 110341 4796
rect 107699 4044 107765 4045
rect 107699 3980 107700 4044
rect 107764 3980 107765 4044
rect 107699 3979 107765 3980
rect 108251 4044 108317 4045
rect 108251 3980 108252 4044
rect 108316 3980 108317 4044
rect 108251 3979 108317 3980
rect 109171 4044 109237 4045
rect 109171 3980 109172 4044
rect 109236 3980 109237 4044
rect 109171 3979 109237 3980
rect 109907 4044 109973 4045
rect 109907 3980 109908 4044
rect 109972 3980 109973 4044
rect 109907 3979 109973 3980
rect 107147 3772 107213 3773
rect 107147 3708 107148 3772
rect 107212 3708 107213 3772
rect 107147 3707 107213 3708
rect 107702 370 107762 3979
rect 106046 310 106198 370
rect 105402 0 105462 310
rect 106138 0 106198 310
rect 106874 310 107026 370
rect 107610 310 107762 370
rect 108254 370 108314 3979
rect 109174 370 109234 3979
rect 109910 370 109970 3979
rect 110278 3229 110338 4795
rect 113038 4450 113098 5339
rect 113038 4390 113282 4450
rect 113222 4045 113282 4390
rect 136137 4384 136457 5408
rect 136137 4320 136145 4384
rect 136209 4320 136225 4384
rect 136289 4320 136305 4384
rect 136369 4320 136385 4384
rect 136449 4320 136457 4384
rect 110643 4044 110709 4045
rect 110643 3980 110644 4044
rect 110708 3980 110709 4044
rect 110643 3979 110709 3980
rect 111195 4044 111261 4045
rect 111195 3980 111196 4044
rect 111260 3980 111261 4044
rect 111195 3979 111261 3980
rect 112115 4044 112181 4045
rect 112115 3980 112116 4044
rect 112180 3980 112181 4044
rect 112115 3979 112181 3980
rect 112851 4044 112917 4045
rect 112851 3980 112852 4044
rect 112916 3980 112917 4044
rect 112851 3979 112917 3980
rect 113219 4044 113285 4045
rect 113219 3980 113220 4044
rect 113284 3980 113285 4044
rect 113219 3979 113285 3980
rect 110275 3228 110341 3229
rect 110275 3164 110276 3228
rect 110340 3164 110341 3228
rect 110275 3163 110341 3164
rect 110646 370 110706 3979
rect 108254 310 108406 370
rect 106874 0 106934 310
rect 107610 0 107670 310
rect 108346 0 108406 310
rect 109082 310 109234 370
rect 109818 310 109970 370
rect 110554 310 110706 370
rect 111198 370 111258 3979
rect 112118 370 112178 3979
rect 112854 370 112914 3979
rect 136137 3296 136457 4320
rect 136137 3232 136145 3296
rect 136209 3232 136225 3296
rect 136289 3232 136305 3296
rect 136369 3232 136385 3296
rect 136449 3232 136457 3296
rect 116531 2820 116597 2821
rect 116531 2756 116532 2820
rect 116596 2756 116597 2820
rect 116531 2755 116597 2756
rect 123891 2820 123957 2821
rect 123891 2756 123892 2820
rect 123956 2756 123957 2820
rect 123891 2755 123957 2756
rect 133459 2820 133525 2821
rect 133459 2756 133460 2820
rect 133524 2756 133525 2820
rect 133459 2755 133525 2756
rect 114323 2276 114389 2277
rect 114323 2212 114324 2276
rect 114388 2212 114389 2276
rect 114323 2211 114389 2212
rect 113587 1460 113653 1461
rect 113587 1396 113588 1460
rect 113652 1396 113653 1460
rect 113587 1395 113653 1396
rect 113590 370 113650 1395
rect 114326 370 114386 2211
rect 114875 1460 114941 1461
rect 114875 1396 114876 1460
rect 114940 1396 114941 1460
rect 114875 1395 114941 1396
rect 115611 1460 115677 1461
rect 115611 1396 115612 1460
rect 115676 1396 115677 1460
rect 115611 1395 115677 1396
rect 111198 310 111350 370
rect 109082 0 109142 310
rect 109818 0 109878 310
rect 110554 0 110614 310
rect 111290 0 111350 310
rect 112026 310 112178 370
rect 112762 310 112914 370
rect 113498 310 113650 370
rect 114234 310 114386 370
rect 114878 370 114938 1395
rect 115614 370 115674 1395
rect 116534 370 116594 2755
rect 117267 1460 117333 1461
rect 117267 1396 117268 1460
rect 117332 1396 117333 1460
rect 117267 1395 117333 1396
rect 117270 370 117330 1395
rect 117911 508 117977 509
rect 117911 444 117912 508
rect 117976 444 117977 508
rect 117911 443 117977 444
rect 118647 508 118713 509
rect 118647 444 118648 508
rect 118712 444 118713 508
rect 118647 443 118713 444
rect 119383 508 119449 509
rect 119383 444 119384 508
rect 119448 444 119449 508
rect 119383 443 119449 444
rect 120119 508 120185 509
rect 120119 444 120120 508
rect 120184 444 120185 508
rect 120119 443 120185 444
rect 120855 508 120921 509
rect 120855 444 120856 508
rect 120920 444 120921 508
rect 120855 443 120921 444
rect 121591 508 121657 509
rect 121591 444 121592 508
rect 121656 444 121657 508
rect 121591 443 121657 444
rect 122327 508 122393 509
rect 122327 444 122328 508
rect 122392 444 122393 508
rect 122327 443 122393 444
rect 123063 508 123129 509
rect 123063 444 123064 508
rect 123128 444 123129 508
rect 123063 443 123129 444
rect 114878 310 115030 370
rect 115614 310 115766 370
rect 112026 0 112086 310
rect 112762 0 112822 310
rect 113498 0 113558 310
rect 114234 0 114294 310
rect 114970 0 115030 310
rect 115706 0 115766 310
rect 116442 310 116594 370
rect 117178 310 117330 370
rect 116442 0 116502 310
rect 117178 0 117238 310
rect 117914 0 117974 443
rect 118650 0 118710 443
rect 119386 0 119446 443
rect 120122 0 120182 443
rect 120858 0 120918 443
rect 121594 0 121654 443
rect 122330 0 122390 443
rect 123066 0 123126 443
rect 123894 370 123954 2755
rect 126835 1460 126901 1461
rect 126835 1396 126836 1460
rect 126900 1396 126901 1460
rect 126835 1395 126901 1396
rect 128307 1460 128373 1461
rect 128307 1396 128308 1460
rect 128372 1396 128373 1460
rect 128307 1395 128373 1396
rect 124535 644 124601 645
rect 124535 580 124536 644
rect 124600 580 124601 644
rect 124535 579 124601 580
rect 125271 644 125337 645
rect 125271 580 125272 644
rect 125336 580 125337 644
rect 125271 579 125337 580
rect 126007 644 126073 645
rect 126007 580 126008 644
rect 126072 580 126073 644
rect 126007 579 126073 580
rect 123802 310 123954 370
rect 123802 0 123862 310
rect 124538 0 124598 579
rect 125274 0 125334 579
rect 126010 0 126070 579
rect 126838 370 126898 1395
rect 127479 508 127545 509
rect 127479 444 127480 508
rect 127544 444 127545 508
rect 127479 443 127545 444
rect 126746 310 126898 370
rect 126746 0 126806 310
rect 127482 0 127542 443
rect 128310 370 128370 1395
rect 128951 644 129017 645
rect 128951 580 128952 644
rect 129016 580 129017 644
rect 128951 579 129017 580
rect 130423 644 130489 645
rect 130423 580 130424 644
rect 130488 580 130489 644
rect 130423 579 130489 580
rect 131159 644 131225 645
rect 131159 580 131160 644
rect 131224 580 131225 644
rect 131159 579 131225 580
rect 128218 310 128370 370
rect 128218 0 128278 310
rect 128954 0 129014 579
rect 129687 372 129753 373
rect 129687 308 129688 372
rect 129752 308 129753 372
rect 129687 307 129753 308
rect 129690 0 129750 307
rect 130426 0 130486 579
rect 131162 0 131222 579
rect 131895 372 131961 373
rect 131895 308 131896 372
rect 131960 308 131961 372
rect 131895 307 131961 308
rect 132631 372 132697 373
rect 132631 308 132632 372
rect 132696 308 132697 372
rect 133462 370 133522 2755
rect 136137 2208 136457 3232
rect 144683 3228 144749 3229
rect 144683 3164 144684 3228
rect 144748 3164 144749 3228
rect 144683 3163 144749 3164
rect 136137 2144 136145 2208
rect 136209 2144 136225 2208
rect 136289 2144 136305 2208
rect 136369 2144 136385 2208
rect 136449 2144 136457 2208
rect 134931 1460 134997 1461
rect 134931 1396 134932 1460
rect 134996 1396 134997 1460
rect 134931 1395 134997 1396
rect 134103 644 134169 645
rect 134103 580 134104 644
rect 134168 580 134169 644
rect 134103 579 134169 580
rect 132631 307 132697 308
rect 133370 310 133522 370
rect 131898 0 131958 307
rect 132634 0 132694 307
rect 133370 0 133430 310
rect 134106 0 134166 579
rect 134934 370 134994 1395
rect 136137 1120 136457 2144
rect 140267 1868 140333 1869
rect 140267 1804 140268 1868
rect 140332 1804 140333 1868
rect 140267 1803 140333 1804
rect 137323 1460 137389 1461
rect 137323 1396 137324 1460
rect 137388 1396 137389 1460
rect 137323 1395 137389 1396
rect 136137 1056 136145 1120
rect 136209 1056 136225 1120
rect 136289 1056 136305 1120
rect 136369 1056 136385 1120
rect 136449 1056 136457 1120
rect 136137 1040 136457 1056
rect 134842 310 134994 370
rect 134842 0 134902 310
rect 137326 0 137386 1395
rect 139531 1052 139597 1053
rect 139531 988 139532 1052
rect 139596 988 139597 1052
rect 139531 987 139597 988
rect 138795 780 138861 781
rect 138795 716 138796 780
rect 138860 716 138861 780
rect 138795 715 138861 716
rect 138059 644 138125 645
rect 138059 580 138060 644
rect 138124 580 138125 644
rect 138059 579 138125 580
rect 138062 0 138122 579
rect 138798 0 138858 715
rect 139534 0 139594 987
rect 140270 0 140330 1803
rect 141003 1460 141069 1461
rect 141003 1396 141004 1460
rect 141068 1396 141069 1460
rect 141003 1395 141069 1396
rect 141006 0 141066 1395
rect 141739 780 141805 781
rect 141739 716 141740 780
rect 141804 716 141805 780
rect 141739 715 141805 716
rect 142475 780 142541 781
rect 142475 716 142476 780
rect 142540 716 142541 780
rect 142475 715 142541 716
rect 141742 0 141802 715
rect 142478 0 142538 715
rect 143211 644 143277 645
rect 143211 580 143212 644
rect 143276 580 143277 644
rect 143211 579 143277 580
rect 143214 0 143274 579
rect 143947 508 144013 509
rect 143947 444 143948 508
rect 144012 444 144013 508
rect 143947 443 144013 444
rect 143950 0 144010 443
rect 144686 0 144746 3163
rect 149099 2956 149165 2957
rect 149099 2892 149100 2956
rect 149164 2892 149165 2956
rect 149099 2891 149165 2892
rect 145419 2820 145485 2821
rect 145419 2756 145420 2820
rect 145484 2756 145485 2820
rect 145419 2755 145485 2756
rect 145422 0 145482 2755
rect 146155 780 146221 781
rect 146155 716 146156 780
rect 146220 716 146221 780
rect 146155 715 146221 716
rect 148363 780 148429 781
rect 148363 716 148364 780
rect 148428 716 148429 780
rect 148363 715 148429 716
rect 146158 0 146218 715
rect 147627 644 147693 645
rect 147627 580 147628 644
rect 147692 580 147693 644
rect 147627 579 147693 580
rect 146891 372 146957 373
rect 146891 308 146892 372
rect 146956 308 146957 372
rect 146891 307 146957 308
rect 146894 0 146954 307
rect 147630 0 147690 579
rect 148366 0 148426 715
rect 149102 0 149162 2891
rect 151678 2413 151738 6563
rect 169936 6016 170256 7040
rect 169936 5952 169944 6016
rect 170008 5952 170024 6016
rect 170088 5952 170104 6016
rect 170168 5952 170184 6016
rect 170248 5952 170256 6016
rect 151859 5676 151925 5677
rect 151859 5612 151860 5676
rect 151924 5612 151925 5676
rect 151859 5611 151925 5612
rect 151675 2412 151741 2413
rect 151675 2348 151676 2412
rect 151740 2348 151741 2412
rect 151675 2347 151741 2348
rect 150571 1460 150637 1461
rect 150571 1396 150572 1460
rect 150636 1396 150637 1460
rect 150571 1395 150637 1396
rect 149835 780 149901 781
rect 149835 716 149836 780
rect 149900 716 149901 780
rect 149835 715 149901 716
rect 149838 0 149898 715
rect 150574 0 150634 1395
rect 151862 781 151922 5611
rect 169936 4928 170256 5952
rect 169936 4864 169944 4928
rect 170008 4864 170024 4928
rect 170088 4864 170104 4928
rect 170168 4864 170184 4928
rect 170248 4864 170256 4928
rect 153147 4044 153213 4045
rect 153147 3980 153148 4044
rect 153212 3980 153213 4044
rect 153147 3979 153213 3980
rect 152043 1460 152109 1461
rect 152043 1396 152044 1460
rect 152108 1396 152109 1460
rect 152043 1395 152109 1396
rect 151859 780 151925 781
rect 151859 716 151860 780
rect 151924 716 151925 780
rect 151859 715 151925 716
rect 151307 644 151373 645
rect 151307 580 151308 644
rect 151372 580 151373 644
rect 151307 579 151373 580
rect 151310 0 151370 579
rect 152046 0 152106 1395
rect 152779 1324 152845 1325
rect 152779 1260 152780 1324
rect 152844 1260 152845 1324
rect 152779 1259 152845 1260
rect 152782 0 152842 1259
rect 153150 237 153210 3979
rect 169936 3840 170256 4864
rect 169936 3776 169944 3840
rect 170008 3776 170024 3840
rect 170088 3776 170104 3840
rect 170168 3776 170184 3840
rect 170248 3776 170256 3840
rect 154251 3364 154317 3365
rect 154251 3300 154252 3364
rect 154316 3300 154317 3364
rect 154251 3299 154317 3300
rect 153515 2956 153581 2957
rect 153515 2892 153516 2956
rect 153580 2892 153581 2956
rect 153515 2891 153581 2892
rect 153147 236 153213 237
rect 153147 172 153148 236
rect 153212 172 153213 236
rect 153147 171 153213 172
rect 153518 0 153578 2891
rect 154254 0 154314 3299
rect 154987 2956 155053 2957
rect 154987 2892 154988 2956
rect 155052 2892 155053 2956
rect 154987 2891 155053 2892
rect 154990 0 155050 2891
rect 156459 2820 156525 2821
rect 156459 2756 156460 2820
rect 156524 2756 156525 2820
rect 156459 2755 156525 2756
rect 155723 1460 155789 1461
rect 155723 1396 155724 1460
rect 155788 1396 155789 1460
rect 155723 1395 155789 1396
rect 155726 0 155786 1395
rect 156462 0 156522 2755
rect 169936 2752 170256 3776
rect 203734 9824 204054 9840
rect 211475 9828 211476 9892
rect 211540 9828 211541 9892
rect 211475 9827 211541 9828
rect 203734 9760 203742 9824
rect 203806 9760 203822 9824
rect 203886 9760 203902 9824
rect 203966 9760 203982 9824
rect 204046 9760 204054 9824
rect 203734 8736 204054 9760
rect 215158 9621 215218 10880
rect 215894 10165 215954 10880
rect 215891 10164 215957 10165
rect 215891 10100 215892 10164
rect 215956 10100 215957 10164
rect 215891 10099 215957 10100
rect 216630 9893 216690 10880
rect 217366 10165 217426 10880
rect 218102 10573 218162 10880
rect 218099 10572 218165 10573
rect 218099 10508 218100 10572
rect 218164 10508 218165 10572
rect 218099 10507 218165 10508
rect 218838 10165 218898 10880
rect 219574 10165 219634 10880
rect 220310 10301 220370 10880
rect 221046 10437 221106 10880
rect 221043 10436 221109 10437
rect 221043 10372 221044 10436
rect 221108 10372 221109 10436
rect 221043 10371 221109 10372
rect 220307 10300 220373 10301
rect 220307 10236 220308 10300
rect 220372 10236 220373 10300
rect 220307 10235 220373 10236
rect 217363 10164 217429 10165
rect 217363 10100 217364 10164
rect 217428 10100 217429 10164
rect 217363 10099 217429 10100
rect 218835 10164 218901 10165
rect 218835 10100 218836 10164
rect 218900 10100 218901 10164
rect 218835 10099 218901 10100
rect 219571 10164 219637 10165
rect 219571 10100 219572 10164
rect 219636 10100 219637 10164
rect 219571 10099 219637 10100
rect 221782 9893 221842 10880
rect 222518 10165 222578 10880
rect 223254 10165 223314 10880
rect 222515 10164 222581 10165
rect 222515 10100 222516 10164
rect 222580 10100 222581 10164
rect 222515 10099 222581 10100
rect 223251 10164 223317 10165
rect 223251 10100 223252 10164
rect 223316 10100 223317 10164
rect 223251 10099 223317 10100
rect 216627 9892 216693 9893
rect 216627 9828 216628 9892
rect 216692 9828 216693 9892
rect 216627 9827 216693 9828
rect 221779 9892 221845 9893
rect 221779 9828 221780 9892
rect 221844 9828 221845 9892
rect 221779 9827 221845 9828
rect 215155 9620 215221 9621
rect 215155 9556 215156 9620
rect 215220 9556 215221 9620
rect 215155 9555 215221 9556
rect 223990 9485 224050 10880
rect 223987 9484 224053 9485
rect 223987 9420 223988 9484
rect 224052 9420 224053 9484
rect 223987 9419 224053 9420
rect 213867 9076 213933 9077
rect 213867 9012 213868 9076
rect 213932 9012 213933 9076
rect 213867 9011 213933 9012
rect 203734 8672 203742 8736
rect 203806 8672 203822 8736
rect 203886 8672 203902 8736
rect 203966 8672 203982 8736
rect 204046 8672 204054 8736
rect 203734 7648 204054 8672
rect 203734 7584 203742 7648
rect 203806 7584 203822 7648
rect 203886 7584 203902 7648
rect 203966 7584 203982 7648
rect 204046 7584 204054 7648
rect 203734 6560 204054 7584
rect 203734 6496 203742 6560
rect 203806 6496 203822 6560
rect 203886 6496 203902 6560
rect 203966 6496 203982 6560
rect 204046 6496 204054 6560
rect 203734 5472 204054 6496
rect 213870 5813 213930 9011
rect 224726 8669 224786 10880
rect 225462 8669 225522 10880
rect 226011 8804 226077 8805
rect 226011 8740 226012 8804
rect 226076 8740 226077 8804
rect 226011 8739 226077 8740
rect 224723 8668 224789 8669
rect 224723 8604 224724 8668
rect 224788 8604 224789 8668
rect 224723 8603 224789 8604
rect 225459 8668 225525 8669
rect 225459 8604 225460 8668
rect 225524 8604 225525 8668
rect 225459 8603 225525 8604
rect 224355 8396 224421 8397
rect 224355 8332 224356 8396
rect 224420 8332 224421 8396
rect 224355 8331 224421 8332
rect 219939 7580 220005 7581
rect 219939 7516 219940 7580
rect 220004 7516 220005 7580
rect 219939 7515 220005 7516
rect 213867 5812 213933 5813
rect 213867 5748 213868 5812
rect 213932 5748 213933 5812
rect 213867 5747 213933 5748
rect 203734 5408 203742 5472
rect 203806 5408 203822 5472
rect 203886 5408 203902 5472
rect 203966 5408 203982 5472
rect 204046 5408 204054 5472
rect 203734 4384 204054 5408
rect 219942 5269 220002 7515
rect 220859 6764 220925 6765
rect 220859 6700 220860 6764
rect 220924 6700 220925 6764
rect 220859 6699 220925 6700
rect 220862 5541 220922 6699
rect 220859 5540 220925 5541
rect 220859 5476 220860 5540
rect 220924 5476 220925 5540
rect 220859 5475 220925 5476
rect 219939 5268 220005 5269
rect 219939 5204 219940 5268
rect 220004 5204 220005 5268
rect 219939 5203 220005 5204
rect 203734 4320 203742 4384
rect 203806 4320 203822 4384
rect 203886 4320 203902 4384
rect 203966 4320 203982 4384
rect 204046 4320 204054 4384
rect 203734 3296 204054 4320
rect 215155 4044 215221 4045
rect 215155 3980 215156 4044
rect 215220 3980 215221 4044
rect 215155 3979 215221 3980
rect 223987 4044 224053 4045
rect 223987 3980 223988 4044
rect 224052 3980 224053 4044
rect 223987 3979 224053 3980
rect 203734 3232 203742 3296
rect 203806 3232 203822 3296
rect 203886 3232 203902 3296
rect 203966 3232 203982 3296
rect 204046 3232 204054 3296
rect 189947 2820 190013 2821
rect 189947 2756 189948 2820
rect 190012 2756 190013 2820
rect 189947 2755 190013 2756
rect 191419 2820 191485 2821
rect 191419 2756 191420 2820
rect 191484 2756 191485 2820
rect 191419 2755 191485 2756
rect 198043 2820 198109 2821
rect 198043 2756 198044 2820
rect 198108 2756 198109 2820
rect 198043 2755 198109 2756
rect 199515 2820 199581 2821
rect 199515 2756 199516 2820
rect 199580 2756 199581 2820
rect 199515 2755 199581 2756
rect 200987 2820 201053 2821
rect 200987 2756 200988 2820
rect 201052 2756 201053 2820
rect 200987 2755 201053 2756
rect 169936 2688 169944 2752
rect 170008 2688 170024 2752
rect 170088 2688 170104 2752
rect 170168 2688 170184 2752
rect 170248 2688 170256 2752
rect 169936 1664 170256 2688
rect 169936 1600 169944 1664
rect 170008 1600 170024 1664
rect 170088 1600 170104 1664
rect 170168 1600 170184 1664
rect 170248 1600 170256 1664
rect 157195 1460 157261 1461
rect 157195 1396 157196 1460
rect 157260 1396 157261 1460
rect 157195 1395 157261 1396
rect 168235 1460 168301 1461
rect 168235 1396 168236 1460
rect 168300 1396 168301 1460
rect 168235 1395 168301 1396
rect 157198 0 157258 1395
rect 157931 1324 157997 1325
rect 157931 1260 157932 1324
rect 157996 1260 157997 1324
rect 157931 1259 157997 1260
rect 157934 0 157994 1259
rect 158667 1188 158733 1189
rect 158667 1124 158668 1188
rect 158732 1124 158733 1188
rect 158667 1123 158733 1124
rect 160139 1188 160205 1189
rect 160139 1124 160140 1188
rect 160204 1124 160205 1188
rect 160139 1123 160205 1124
rect 161611 1188 161677 1189
rect 161611 1124 161612 1188
rect 161676 1124 161677 1188
rect 161611 1123 161677 1124
rect 163819 1188 163885 1189
rect 163819 1124 163820 1188
rect 163884 1124 163885 1188
rect 163819 1123 163885 1124
rect 165291 1188 165357 1189
rect 165291 1124 165292 1188
rect 165356 1124 165357 1188
rect 165291 1123 165357 1124
rect 166027 1188 166093 1189
rect 166027 1124 166028 1188
rect 166092 1124 166093 1188
rect 166027 1123 166093 1124
rect 166763 1188 166829 1189
rect 166763 1124 166764 1188
rect 166828 1124 166829 1188
rect 166763 1123 166829 1124
rect 158670 0 158730 1123
rect 159403 644 159469 645
rect 159403 580 159404 644
rect 159468 580 159469 644
rect 159403 579 159469 580
rect 159406 0 159466 579
rect 160142 0 160202 1123
rect 160875 372 160941 373
rect 160875 308 160876 372
rect 160940 308 160941 372
rect 160875 307 160941 308
rect 160878 0 160938 307
rect 161614 0 161674 1123
rect 162347 644 162413 645
rect 162347 580 162348 644
rect 162412 580 162413 644
rect 162347 579 162413 580
rect 163083 644 163149 645
rect 163083 580 163084 644
rect 163148 580 163149 644
rect 163083 579 163149 580
rect 162350 0 162410 579
rect 163086 0 163146 579
rect 163822 0 163882 1123
rect 164555 644 164621 645
rect 164555 580 164556 644
rect 164620 580 164621 644
rect 164555 579 164621 580
rect 164558 0 164618 579
rect 165294 0 165354 1123
rect 166030 0 166090 1123
rect 166766 0 166826 1123
rect 167499 372 167565 373
rect 167499 308 167500 372
rect 167564 308 167565 372
rect 167499 307 167565 308
rect 167502 0 167562 307
rect 168238 0 168298 1395
rect 169936 1040 170256 1600
rect 186267 1460 186333 1461
rect 186267 1396 186268 1460
rect 186332 1396 186333 1460
rect 186267 1395 186333 1396
rect 168971 644 169037 645
rect 168971 580 168972 644
rect 169036 580 169037 644
rect 168971 579 169037 580
rect 171455 644 171521 645
rect 171455 580 171456 644
rect 171520 580 171521 644
rect 171455 579 171521 580
rect 172191 644 172257 645
rect 172191 580 172192 644
rect 172256 580 172257 644
rect 172191 579 172257 580
rect 172927 644 172993 645
rect 172927 580 172928 644
rect 172992 580 172993 644
rect 172927 579 172993 580
rect 173663 644 173729 645
rect 173663 580 173664 644
rect 173728 580 173729 644
rect 173663 579 173729 580
rect 174399 644 174465 645
rect 174399 580 174400 644
rect 174464 580 174465 644
rect 174399 579 174465 580
rect 175135 644 175201 645
rect 175135 580 175136 644
rect 175200 580 175201 644
rect 175135 579 175201 580
rect 176607 644 176673 645
rect 176607 580 176608 644
rect 176672 580 176673 644
rect 176607 579 176673 580
rect 177343 644 177409 645
rect 177343 580 177344 644
rect 177408 580 177409 644
rect 177343 579 177409 580
rect 178079 644 178145 645
rect 178079 580 178080 644
rect 178144 580 178145 644
rect 178079 579 178145 580
rect 178815 644 178881 645
rect 178815 580 178816 644
rect 178880 580 178881 644
rect 178815 579 178881 580
rect 179551 644 179617 645
rect 179551 580 179552 644
rect 179616 580 179617 644
rect 179551 579 179617 580
rect 180287 644 180353 645
rect 180287 580 180288 644
rect 180352 580 180353 644
rect 180287 579 180353 580
rect 168974 0 169034 579
rect 171458 0 171518 579
rect 172194 0 172254 579
rect 172930 0 172990 579
rect 173666 0 173726 579
rect 174402 0 174462 579
rect 175138 0 175198 579
rect 175871 508 175937 509
rect 175871 444 175872 508
rect 175936 444 175937 508
rect 175871 443 175937 444
rect 175874 0 175934 443
rect 176610 0 176670 579
rect 177346 0 177406 579
rect 178082 0 178142 579
rect 178818 0 178878 579
rect 179554 0 179614 579
rect 180290 0 180350 579
rect 181759 508 181825 509
rect 181759 444 181760 508
rect 181824 444 181825 508
rect 181759 443 181825 444
rect 182495 508 182561 509
rect 182495 444 182496 508
rect 182560 444 182561 508
rect 182495 443 182561 444
rect 183231 508 183297 509
rect 183231 444 183232 508
rect 183296 444 183297 508
rect 183231 443 183297 444
rect 183967 508 184033 509
rect 183967 444 183968 508
rect 184032 444 184033 508
rect 183967 443 184033 444
rect 184703 508 184769 509
rect 184703 444 184704 508
rect 184768 444 184769 508
rect 184703 443 184769 444
rect 185439 508 185505 509
rect 185439 444 185440 508
rect 185504 444 185505 508
rect 185439 443 185505 444
rect 181023 372 181089 373
rect 181023 308 181024 372
rect 181088 308 181089 372
rect 181023 307 181089 308
rect 181026 0 181086 307
rect 181762 0 181822 443
rect 182498 0 182558 443
rect 183234 0 183294 443
rect 183970 0 184030 443
rect 184706 0 184766 443
rect 185442 0 185502 443
rect 186270 370 186330 1395
rect 186911 508 186977 509
rect 186911 444 186912 508
rect 186976 444 186977 508
rect 186911 443 186977 444
rect 187647 508 187713 509
rect 187647 444 187648 508
rect 187712 444 187713 508
rect 187647 443 187713 444
rect 188383 508 188449 509
rect 188383 444 188384 508
rect 188448 444 188449 508
rect 188383 443 188449 444
rect 189119 508 189185 509
rect 189119 444 189120 508
rect 189184 444 189185 508
rect 189119 443 189185 444
rect 186178 310 186330 370
rect 186178 0 186238 310
rect 186914 0 186974 443
rect 187650 0 187710 443
rect 188386 0 188446 443
rect 189122 0 189182 443
rect 189950 370 190010 2755
rect 190591 508 190657 509
rect 190591 444 190592 508
rect 190656 444 190657 508
rect 190591 443 190657 444
rect 189858 310 190010 370
rect 189858 0 189918 310
rect 190594 0 190654 443
rect 191422 370 191482 2755
rect 194363 1868 194429 1869
rect 194363 1804 194364 1868
rect 194428 1804 194429 1868
rect 194363 1803 194429 1804
rect 195835 1868 195901 1869
rect 195835 1804 195836 1868
rect 195900 1804 195901 1868
rect 195835 1803 195901 1804
rect 192799 508 192865 509
rect 192799 444 192800 508
rect 192864 444 192865 508
rect 192799 443 192865 444
rect 193535 508 193601 509
rect 193535 444 193536 508
rect 193600 444 193601 508
rect 193535 443 193601 444
rect 191330 310 191482 370
rect 192063 372 192129 373
rect 191330 0 191390 310
rect 192063 308 192064 372
rect 192128 308 192129 372
rect 192063 307 192129 308
rect 192066 0 192126 307
rect 192802 0 192862 443
rect 193538 0 193598 443
rect 194366 370 194426 1803
rect 195007 508 195073 509
rect 195007 444 195008 508
rect 195072 444 195073 508
rect 195007 443 195073 444
rect 194274 310 194426 370
rect 194274 0 194334 310
rect 195010 0 195070 443
rect 195838 370 195898 1803
rect 197307 1460 197373 1461
rect 197307 1396 197308 1460
rect 197372 1396 197373 1460
rect 197307 1395 197373 1396
rect 196479 508 196545 509
rect 196479 444 196480 508
rect 196544 444 196545 508
rect 196479 443 196545 444
rect 195746 310 195898 370
rect 195746 0 195806 310
rect 196482 0 196542 443
rect 197310 370 197370 1395
rect 198046 370 198106 2755
rect 198687 508 198753 509
rect 198687 444 198688 508
rect 198752 444 198753 508
rect 198687 443 198753 444
rect 197218 310 197370 370
rect 197954 310 198106 370
rect 197218 0 197278 310
rect 197954 0 198014 310
rect 198690 0 198750 443
rect 199518 370 199578 2755
rect 200159 508 200225 509
rect 200159 444 200160 508
rect 200224 444 200225 508
rect 200159 443 200225 444
rect 199426 310 199578 370
rect 199426 0 199486 310
rect 200162 0 200222 443
rect 200990 370 201050 2755
rect 203734 2208 204054 3232
rect 211475 3092 211541 3093
rect 211475 3028 211476 3092
rect 211540 3028 211541 3092
rect 211475 3027 211541 3028
rect 210739 2820 210805 2821
rect 210739 2756 210740 2820
rect 210804 2756 210805 2820
rect 210739 2755 210805 2756
rect 203734 2144 203742 2208
rect 203806 2144 203822 2208
rect 203886 2144 203902 2208
rect 203966 2144 203982 2208
rect 204046 2144 204054 2208
rect 201723 1460 201789 1461
rect 201723 1396 201724 1460
rect 201788 1396 201789 1460
rect 201723 1395 201789 1396
rect 201726 370 201786 1395
rect 203734 1120 204054 2144
rect 210003 1460 210069 1461
rect 210003 1396 210004 1460
rect 210068 1396 210069 1460
rect 210003 1395 210069 1396
rect 203734 1056 203742 1120
rect 203806 1056 203822 1120
rect 203886 1056 203902 1120
rect 203966 1056 203982 1120
rect 204046 1056 204054 1120
rect 203734 1040 204054 1056
rect 205587 916 205653 917
rect 205587 852 205588 916
rect 205652 852 205653 916
rect 205587 851 205653 852
rect 206323 916 206389 917
rect 206323 852 206324 916
rect 206388 852 206389 916
rect 206323 851 206389 852
rect 207059 916 207125 917
rect 207059 852 207060 916
rect 207124 852 207125 916
rect 207059 851 207125 852
rect 208531 916 208597 917
rect 208531 852 208532 916
rect 208596 852 208597 916
rect 208531 851 208597 852
rect 202367 508 202433 509
rect 202367 444 202368 508
rect 202432 444 202433 508
rect 202367 443 202433 444
rect 203103 508 203169 509
rect 203103 444 203104 508
rect 203168 444 203169 508
rect 203103 443 203169 444
rect 200898 310 201050 370
rect 201634 310 201786 370
rect 200898 0 200958 310
rect 201634 0 201694 310
rect 202370 0 202430 443
rect 203106 0 203166 443
rect 205590 0 205650 851
rect 206326 0 206386 851
rect 207062 0 207122 851
rect 207795 372 207861 373
rect 207795 308 207796 372
rect 207860 308 207861 372
rect 207795 307 207861 308
rect 207798 0 207858 307
rect 208534 0 208594 851
rect 209267 508 209333 509
rect 209267 444 209268 508
rect 209332 444 209333 508
rect 209267 443 209333 444
rect 209270 0 209330 443
rect 210006 0 210066 1395
rect 210742 0 210802 2755
rect 211478 0 211538 3027
rect 212211 1868 212277 1869
rect 212211 1804 212212 1868
rect 212276 1804 212277 1868
rect 212211 1803 212277 1804
rect 212214 0 212274 1803
rect 213683 508 213749 509
rect 213683 444 213684 508
rect 213748 444 213749 508
rect 213683 443 213749 444
rect 212947 372 213013 373
rect 212947 308 212948 372
rect 213012 308 213013 372
rect 212947 307 213013 308
rect 212950 0 213010 307
rect 213686 0 213746 443
rect 214419 372 214485 373
rect 214419 308 214420 372
rect 214484 308 214485 372
rect 214419 307 214485 308
rect 214422 0 214482 307
rect 215158 0 215218 3979
rect 218835 3772 218901 3773
rect 218835 3708 218836 3772
rect 218900 3708 218901 3772
rect 218835 3707 218901 3708
rect 223251 3772 223317 3773
rect 223251 3708 223252 3772
rect 223316 3708 223317 3772
rect 223251 3707 223317 3708
rect 217363 3228 217429 3229
rect 217363 3164 217364 3228
rect 217428 3164 217429 3228
rect 217363 3163 217429 3164
rect 216627 2956 216693 2957
rect 216627 2892 216628 2956
rect 216692 2892 216693 2956
rect 216627 2891 216693 2892
rect 215891 780 215957 781
rect 215891 716 215892 780
rect 215956 716 215957 780
rect 215891 715 215957 716
rect 215894 0 215954 715
rect 216630 0 216690 2891
rect 217366 0 217426 3163
rect 218099 1460 218165 1461
rect 218099 1396 218100 1460
rect 218164 1396 218165 1460
rect 218099 1395 218165 1396
rect 218102 0 218162 1395
rect 218838 0 218898 3707
rect 221043 3228 221109 3229
rect 221043 3164 221044 3228
rect 221108 3164 221109 3228
rect 221043 3163 221109 3164
rect 219571 1460 219637 1461
rect 219571 1396 219572 1460
rect 219636 1396 219637 1460
rect 219571 1395 219637 1396
rect 219574 0 219634 1395
rect 220307 372 220373 373
rect 220307 308 220308 372
rect 220372 308 220373 372
rect 220307 307 220373 308
rect 220310 0 220370 307
rect 221046 0 221106 3163
rect 222515 1460 222581 1461
rect 222515 1396 222516 1460
rect 222580 1396 222581 1460
rect 222515 1395 222581 1396
rect 221779 644 221845 645
rect 221779 580 221780 644
rect 221844 580 221845 644
rect 221779 579 221845 580
rect 221782 0 221842 579
rect 222518 0 222578 1395
rect 223254 0 223314 3707
rect 223990 3637 224050 3979
rect 223987 3636 224053 3637
rect 223987 3572 223988 3636
rect 224052 3572 224053 3636
rect 223987 3571 224053 3572
rect 224358 2821 224418 8331
rect 225091 4860 225157 4861
rect 225091 4796 225092 4860
rect 225156 4796 225157 4860
rect 225091 4795 225157 4796
rect 224355 2820 224421 2821
rect 224355 2756 224356 2820
rect 224420 2756 224421 2820
rect 224355 2755 224421 2756
rect 223987 1188 224053 1189
rect 223987 1124 223988 1188
rect 224052 1124 224053 1188
rect 223987 1123 224053 1124
rect 223990 0 224050 1123
rect 225094 781 225154 4795
rect 226014 3909 226074 8739
rect 226198 8669 226258 10880
rect 226934 8669 226994 10880
rect 227670 9485 227730 10880
rect 228406 9485 228466 10880
rect 227667 9484 227733 9485
rect 227667 9420 227668 9484
rect 227732 9420 227733 9484
rect 227667 9419 227733 9420
rect 228403 9484 228469 9485
rect 228403 9420 228404 9484
rect 228468 9420 228469 9484
rect 228403 9419 228469 9420
rect 227483 8940 227549 8941
rect 227483 8876 227484 8940
rect 227548 8876 227549 8940
rect 227483 8875 227549 8876
rect 226195 8668 226261 8669
rect 226195 8604 226196 8668
rect 226260 8604 226261 8668
rect 226195 8603 226261 8604
rect 226931 8668 226997 8669
rect 226931 8604 226932 8668
rect 226996 8604 226997 8668
rect 226931 8603 226997 8604
rect 227299 8532 227365 8533
rect 227299 8468 227300 8532
rect 227364 8468 227365 8532
rect 227299 8467 227365 8468
rect 226195 4588 226261 4589
rect 226195 4524 226196 4588
rect 226260 4524 226261 4588
rect 226195 4523 226261 4524
rect 226011 3908 226077 3909
rect 226011 3844 226012 3908
rect 226076 3844 226077 3908
rect 226011 3843 226077 3844
rect 226198 2957 226258 4523
rect 227302 3773 227362 8467
rect 227486 6765 227546 8875
rect 229142 8669 229202 10880
rect 229878 9485 229938 10880
rect 229875 9484 229941 9485
rect 229875 9420 229876 9484
rect 229940 9420 229941 9484
rect 229875 9419 229941 9420
rect 230614 8669 230674 10880
rect 231350 8669 231410 10880
rect 232086 9485 232146 10880
rect 232083 9484 232149 9485
rect 232083 9420 232084 9484
rect 232148 9420 232149 9484
rect 232083 9419 232149 9420
rect 232822 8669 232882 10880
rect 233558 9485 233618 10880
rect 233555 9484 233621 9485
rect 233555 9420 233556 9484
rect 233620 9420 233621 9484
rect 233555 9419 233621 9420
rect 234294 8669 234354 10880
rect 229139 8668 229205 8669
rect 229139 8604 229140 8668
rect 229204 8604 229205 8668
rect 229139 8603 229205 8604
rect 230611 8668 230677 8669
rect 230611 8604 230612 8668
rect 230676 8604 230677 8668
rect 230611 8603 230677 8604
rect 231347 8668 231413 8669
rect 231347 8604 231348 8668
rect 231412 8604 231413 8668
rect 231347 8603 231413 8604
rect 232819 8668 232885 8669
rect 232819 8604 232820 8668
rect 232884 8604 232885 8668
rect 232819 8603 232885 8604
rect 234291 8668 234357 8669
rect 234291 8604 234292 8668
rect 234356 8604 234357 8668
rect 234291 8603 234357 8604
rect 235030 8397 235090 10880
rect 235766 9485 235826 10880
rect 235763 9484 235829 9485
rect 235763 9420 235764 9484
rect 235828 9420 235829 9484
rect 235763 9419 235829 9420
rect 236502 9213 236562 10880
rect 236499 9212 236565 9213
rect 236499 9148 236500 9212
rect 236564 9148 236565 9212
rect 236499 9147 236565 9148
rect 237238 8669 237298 10880
rect 239722 10301 239782 10880
rect 240458 10301 240518 10880
rect 241194 10301 241254 10880
rect 241930 10301 241990 10880
rect 242666 10301 242726 10880
rect 243402 10301 243462 10880
rect 244138 10301 244198 10880
rect 244874 10301 244934 10880
rect 245610 10437 245670 10880
rect 245607 10436 245673 10437
rect 245607 10372 245608 10436
rect 245672 10372 245673 10436
rect 245607 10371 245673 10372
rect 246346 10301 246406 10880
rect 247082 10301 247142 10880
rect 247818 10301 247878 10880
rect 248554 10301 248614 10880
rect 249290 10301 249350 10880
rect 250026 10301 250086 10880
rect 250762 10301 250822 10880
rect 251498 10301 251558 10880
rect 252234 10301 252294 10880
rect 252970 10437 253030 10880
rect 252967 10436 253033 10437
rect 252967 10372 252968 10436
rect 253032 10372 253033 10436
rect 252967 10371 253033 10372
rect 253706 10301 253766 10880
rect 254442 10301 254502 10880
rect 255178 10301 255238 10880
rect 255914 10301 255974 10880
rect 256650 10301 256710 10880
rect 257386 10301 257446 10880
rect 258122 10301 258182 10880
rect 258858 10301 258918 10880
rect 259594 10301 259654 10880
rect 260330 10301 260390 10880
rect 261066 10437 261126 10880
rect 261063 10436 261129 10437
rect 261063 10372 261064 10436
rect 261128 10372 261129 10436
rect 261063 10371 261129 10372
rect 261802 10301 261862 10880
rect 262538 10301 262598 10880
rect 263274 10301 263334 10880
rect 264010 10301 264070 10880
rect 239719 10300 239785 10301
rect 239719 10236 239720 10300
rect 239784 10236 239785 10300
rect 239719 10235 239785 10236
rect 240455 10300 240521 10301
rect 240455 10236 240456 10300
rect 240520 10236 240521 10300
rect 240455 10235 240521 10236
rect 241191 10300 241257 10301
rect 241191 10236 241192 10300
rect 241256 10236 241257 10300
rect 241191 10235 241257 10236
rect 241927 10300 241993 10301
rect 241927 10236 241928 10300
rect 241992 10236 241993 10300
rect 241927 10235 241993 10236
rect 242663 10300 242729 10301
rect 242663 10236 242664 10300
rect 242728 10236 242729 10300
rect 242663 10235 242729 10236
rect 243399 10300 243465 10301
rect 243399 10236 243400 10300
rect 243464 10236 243465 10300
rect 243399 10235 243465 10236
rect 244135 10300 244201 10301
rect 244135 10236 244136 10300
rect 244200 10236 244201 10300
rect 244135 10235 244201 10236
rect 244871 10300 244937 10301
rect 244871 10236 244872 10300
rect 244936 10236 244937 10300
rect 244871 10235 244937 10236
rect 246343 10300 246409 10301
rect 246343 10236 246344 10300
rect 246408 10236 246409 10300
rect 246343 10235 246409 10236
rect 247079 10300 247145 10301
rect 247079 10236 247080 10300
rect 247144 10236 247145 10300
rect 247079 10235 247145 10236
rect 247815 10300 247881 10301
rect 247815 10236 247816 10300
rect 247880 10236 247881 10300
rect 247815 10235 247881 10236
rect 248551 10300 248617 10301
rect 248551 10236 248552 10300
rect 248616 10236 248617 10300
rect 248551 10235 248617 10236
rect 249287 10300 249353 10301
rect 249287 10236 249288 10300
rect 249352 10236 249353 10300
rect 249287 10235 249353 10236
rect 250023 10300 250089 10301
rect 250023 10236 250024 10300
rect 250088 10236 250089 10300
rect 250023 10235 250089 10236
rect 250759 10300 250825 10301
rect 250759 10236 250760 10300
rect 250824 10236 250825 10300
rect 250759 10235 250825 10236
rect 251495 10300 251561 10301
rect 251495 10236 251496 10300
rect 251560 10236 251561 10300
rect 251495 10235 251561 10236
rect 252231 10300 252297 10301
rect 252231 10236 252232 10300
rect 252296 10236 252297 10300
rect 252231 10235 252297 10236
rect 253703 10300 253769 10301
rect 253703 10236 253704 10300
rect 253768 10236 253769 10300
rect 253703 10235 253769 10236
rect 254439 10300 254505 10301
rect 254439 10236 254440 10300
rect 254504 10236 254505 10300
rect 254439 10235 254505 10236
rect 255175 10300 255241 10301
rect 255175 10236 255176 10300
rect 255240 10236 255241 10300
rect 255175 10235 255241 10236
rect 255911 10300 255977 10301
rect 255911 10236 255912 10300
rect 255976 10236 255977 10300
rect 255911 10235 255977 10236
rect 256647 10300 256713 10301
rect 256647 10236 256648 10300
rect 256712 10236 256713 10300
rect 256647 10235 256713 10236
rect 257383 10300 257449 10301
rect 257383 10236 257384 10300
rect 257448 10236 257449 10300
rect 257383 10235 257449 10236
rect 258119 10300 258185 10301
rect 258119 10236 258120 10300
rect 258184 10236 258185 10300
rect 258119 10235 258185 10236
rect 258855 10300 258921 10301
rect 258855 10236 258856 10300
rect 258920 10236 258921 10300
rect 258855 10235 258921 10236
rect 259591 10300 259657 10301
rect 259591 10236 259592 10300
rect 259656 10236 259657 10300
rect 259591 10235 259657 10236
rect 260327 10300 260393 10301
rect 260327 10236 260328 10300
rect 260392 10236 260393 10300
rect 260327 10235 260393 10236
rect 261799 10300 261865 10301
rect 261799 10236 261800 10300
rect 261864 10236 261865 10300
rect 261799 10235 261865 10236
rect 262535 10300 262601 10301
rect 262535 10236 262536 10300
rect 262600 10236 262601 10300
rect 262535 10235 262601 10236
rect 263271 10300 263337 10301
rect 263271 10236 263272 10300
rect 263336 10236 263337 10300
rect 263271 10235 263337 10236
rect 264007 10300 264073 10301
rect 264007 10236 264008 10300
rect 264072 10236 264073 10300
rect 264746 10298 264806 10880
rect 265482 10437 265542 10880
rect 265479 10436 265545 10437
rect 265479 10372 265480 10436
rect 265544 10372 265545 10436
rect 265479 10371 265545 10372
rect 266218 10301 266278 10880
rect 266215 10300 266281 10301
rect 264746 10238 264898 10298
rect 264007 10235 264073 10236
rect 237533 9280 237853 9840
rect 237533 9216 237541 9280
rect 237605 9216 237621 9280
rect 237685 9216 237701 9280
rect 237765 9216 237781 9280
rect 237845 9216 237853 9280
rect 237235 8668 237301 8669
rect 237235 8604 237236 8668
rect 237300 8604 237301 8668
rect 237235 8603 237301 8604
rect 235027 8396 235093 8397
rect 235027 8332 235028 8396
rect 235092 8332 235093 8396
rect 235027 8331 235093 8332
rect 237533 8192 237853 9216
rect 237533 8128 237541 8192
rect 237605 8128 237621 8192
rect 237685 8128 237701 8192
rect 237765 8128 237781 8192
rect 237845 8128 237853 8192
rect 237533 7104 237853 8128
rect 264838 8125 264898 10238
rect 266215 10236 266216 10300
rect 266280 10236 266281 10300
rect 266954 10298 267014 10880
rect 266215 10235 266281 10236
rect 266862 10238 267014 10298
rect 267690 10298 267750 10880
rect 268426 10298 268486 10880
rect 269162 10298 269222 10880
rect 269898 10298 269958 10880
rect 270634 10298 270694 10880
rect 271370 10298 271430 10880
rect 267690 10238 267842 10298
rect 268426 10238 268578 10298
rect 269162 10238 269314 10298
rect 269898 10238 270050 10298
rect 264835 8124 264901 8125
rect 264835 8060 264836 8124
rect 264900 8060 264901 8124
rect 264835 8059 264901 8060
rect 237533 7040 237541 7104
rect 237605 7040 237621 7104
rect 237685 7040 237701 7104
rect 237765 7040 237781 7104
rect 237845 7040 237853 7104
rect 227483 6764 227549 6765
rect 227483 6700 227484 6764
rect 227548 6700 227549 6764
rect 227483 6699 227549 6700
rect 237533 6016 237853 7040
rect 266862 6901 266922 10238
rect 267595 9484 267661 9485
rect 267595 9420 267596 9484
rect 267660 9420 267661 9484
rect 267595 9419 267661 9420
rect 266859 6900 266925 6901
rect 266859 6836 266860 6900
rect 266924 6836 266925 6900
rect 266859 6835 266925 6836
rect 249011 6764 249077 6765
rect 249011 6700 249012 6764
rect 249076 6700 249077 6764
rect 249011 6699 249077 6700
rect 237533 5952 237541 6016
rect 237605 5952 237621 6016
rect 237685 5952 237701 6016
rect 237765 5952 237781 6016
rect 237845 5952 237853 6016
rect 237533 4928 237853 5952
rect 249014 5405 249074 6699
rect 266307 5812 266373 5813
rect 266307 5748 266308 5812
rect 266372 5748 266373 5812
rect 266307 5747 266373 5748
rect 249011 5404 249077 5405
rect 249011 5340 249012 5404
rect 249076 5340 249077 5404
rect 249011 5339 249077 5340
rect 237533 4864 237541 4928
rect 237605 4864 237621 4928
rect 237685 4864 237701 4928
rect 237765 4864 237781 4928
rect 237845 4864 237853 4928
rect 237533 3840 237853 4864
rect 237533 3776 237541 3840
rect 237605 3776 237621 3840
rect 237685 3776 237701 3840
rect 237765 3776 237781 3840
rect 237845 3776 237853 3840
rect 227299 3772 227365 3773
rect 227299 3708 227300 3772
rect 227364 3708 227365 3772
rect 227299 3707 227365 3708
rect 226195 2956 226261 2957
rect 226195 2892 226196 2956
rect 226260 2892 226261 2956
rect 226195 2891 226261 2892
rect 237533 2752 237853 3776
rect 258947 3228 259013 3229
rect 258947 3164 258948 3228
rect 259012 3164 259013 3228
rect 258947 3163 259013 3164
rect 250851 3092 250917 3093
rect 250851 3028 250852 3092
rect 250916 3028 250917 3092
rect 250851 3027 250917 3028
rect 246435 2956 246501 2957
rect 246435 2892 246436 2956
rect 246500 2892 246501 2956
rect 246435 2891 246501 2892
rect 237533 2688 237541 2752
rect 237605 2688 237621 2752
rect 237685 2688 237701 2752
rect 237765 2688 237781 2752
rect 237845 2688 237853 2752
rect 237533 1664 237853 2688
rect 237533 1600 237541 1664
rect 237605 1600 237621 1664
rect 237685 1600 237701 1664
rect 237765 1600 237781 1664
rect 237845 1600 237853 1664
rect 237235 1596 237301 1597
rect 237235 1532 237236 1596
rect 237300 1532 237301 1596
rect 237235 1531 237301 1532
rect 226195 1460 226261 1461
rect 226195 1396 226196 1460
rect 226260 1396 226261 1460
rect 226195 1395 226261 1396
rect 225459 1188 225525 1189
rect 225459 1124 225460 1188
rect 225524 1124 225525 1188
rect 225459 1123 225525 1124
rect 224723 780 224789 781
rect 224723 716 224724 780
rect 224788 716 224789 780
rect 224723 715 224789 716
rect 225091 780 225157 781
rect 225091 716 225092 780
rect 225156 716 225157 780
rect 225091 715 225157 716
rect 224726 0 224786 715
rect 225462 0 225522 1123
rect 226198 0 226258 1395
rect 227667 1188 227733 1189
rect 227667 1124 227668 1188
rect 227732 1124 227733 1188
rect 227667 1123 227733 1124
rect 229875 1188 229941 1189
rect 229875 1124 229876 1188
rect 229940 1124 229941 1188
rect 229875 1123 229941 1124
rect 230611 1188 230677 1189
rect 230611 1124 230612 1188
rect 230676 1124 230677 1188
rect 230611 1123 230677 1124
rect 232083 1188 232149 1189
rect 232083 1124 232084 1188
rect 232148 1124 232149 1188
rect 232083 1123 232149 1124
rect 232819 1188 232885 1189
rect 232819 1124 232820 1188
rect 232884 1124 232885 1188
rect 232819 1123 232885 1124
rect 235027 1188 235093 1189
rect 235027 1124 235028 1188
rect 235092 1124 235093 1188
rect 235027 1123 235093 1124
rect 236499 1188 236565 1189
rect 236499 1124 236500 1188
rect 236564 1124 236565 1188
rect 236499 1123 236565 1124
rect 226931 644 226997 645
rect 226931 580 226932 644
rect 226996 580 226997 644
rect 226931 579 226997 580
rect 226934 0 226994 579
rect 227670 0 227730 1123
rect 228403 644 228469 645
rect 228403 580 228404 644
rect 228468 580 228469 644
rect 228403 579 228469 580
rect 229139 644 229205 645
rect 229139 580 229140 644
rect 229204 580 229205 644
rect 229139 579 229205 580
rect 228406 0 228466 579
rect 229142 0 229202 579
rect 229878 0 229938 1123
rect 230614 0 230674 1123
rect 231347 644 231413 645
rect 231347 580 231348 644
rect 231412 580 231413 644
rect 231347 579 231413 580
rect 231350 0 231410 579
rect 232086 0 232146 1123
rect 232822 0 232882 1123
rect 233555 644 233621 645
rect 233555 580 233556 644
rect 233620 580 233621 644
rect 233555 579 233621 580
rect 234291 644 234357 645
rect 234291 580 234292 644
rect 234356 580 234357 644
rect 234291 579 234357 580
rect 233558 0 233618 579
rect 234294 0 234354 579
rect 235030 0 235090 1123
rect 235763 644 235829 645
rect 235763 580 235764 644
rect 235828 580 235829 644
rect 235763 579 235829 580
rect 235766 0 235826 579
rect 236502 0 236562 1123
rect 237238 0 237298 1531
rect 237533 1040 237853 1600
rect 242755 1460 242821 1461
rect 242755 1396 242756 1460
rect 242820 1396 242821 1460
rect 242755 1395 242821 1396
rect 245699 1460 245765 1461
rect 245699 1396 245700 1460
rect 245764 1396 245765 1460
rect 245699 1395 245765 1396
rect 239719 644 239785 645
rect 239719 580 239720 644
rect 239784 580 239785 644
rect 239719 579 239785 580
rect 240455 644 240521 645
rect 240455 580 240456 644
rect 240520 580 240521 644
rect 240455 579 240521 580
rect 241191 644 241257 645
rect 241191 580 241192 644
rect 241256 580 241257 644
rect 241191 579 241257 580
rect 241927 644 241993 645
rect 241927 580 241928 644
rect 241992 580 241993 644
rect 241927 579 241993 580
rect 239722 0 239782 579
rect 240458 0 240518 579
rect 241194 0 241254 579
rect 241930 0 241990 579
rect 242758 370 242818 1395
rect 243399 644 243465 645
rect 243399 580 243400 644
rect 243464 580 243465 644
rect 243399 579 243465 580
rect 244135 644 244201 645
rect 244135 580 244136 644
rect 244200 580 244201 644
rect 244135 579 244201 580
rect 244871 644 244937 645
rect 244871 580 244872 644
rect 244936 580 244937 644
rect 244871 579 244937 580
rect 242666 310 242818 370
rect 242666 0 242726 310
rect 243402 0 243462 579
rect 244138 0 244198 579
rect 244874 0 244934 579
rect 245702 370 245762 1395
rect 246438 642 246498 2891
rect 249379 1596 249445 1597
rect 249379 1532 249380 1596
rect 249444 1532 249445 1596
rect 249379 1531 249445 1532
rect 248643 1460 248709 1461
rect 248643 1396 248644 1460
rect 248708 1396 248709 1460
rect 248643 1395 248709 1396
rect 245610 310 245762 370
rect 246346 582 246498 642
rect 247079 644 247145 645
rect 245610 0 245670 310
rect 246346 0 246406 582
rect 247079 580 247080 644
rect 247144 580 247145 644
rect 247079 579 247145 580
rect 247815 644 247881 645
rect 247815 580 247816 644
rect 247880 580 247881 644
rect 247815 579 247881 580
rect 247082 0 247142 579
rect 247818 0 247878 579
rect 248646 370 248706 1395
rect 249382 370 249442 1531
rect 250023 644 250089 645
rect 250023 580 250024 644
rect 250088 580 250089 644
rect 250854 642 250914 3027
rect 256003 2956 256069 2957
rect 256003 2892 256004 2956
rect 256068 2892 256069 2956
rect 256003 2891 256069 2892
rect 251587 1596 251653 1597
rect 251587 1532 251588 1596
rect 251652 1532 251653 1596
rect 251587 1531 251653 1532
rect 250023 579 250089 580
rect 250762 582 250914 642
rect 248554 310 248706 370
rect 249290 310 249442 370
rect 248554 0 248614 310
rect 249290 0 249350 310
rect 250026 0 250086 579
rect 250762 0 250822 582
rect 251590 370 251650 1531
rect 252323 1460 252389 1461
rect 252323 1396 252324 1460
rect 252388 1396 252389 1460
rect 252323 1395 252389 1396
rect 252326 370 252386 1395
rect 254439 644 254505 645
rect 254439 580 254440 644
rect 254504 580 254505 644
rect 254439 579 254505 580
rect 255175 644 255241 645
rect 255175 580 255176 644
rect 255240 580 255241 644
rect 256006 642 256066 2891
rect 256739 1596 256805 1597
rect 256739 1532 256740 1596
rect 256804 1532 256805 1596
rect 256739 1531 256805 1532
rect 255175 579 255241 580
rect 255914 582 256066 642
rect 252967 508 253033 509
rect 252967 444 252968 508
rect 253032 444 253033 508
rect 252967 443 253033 444
rect 251498 310 251650 370
rect 252234 310 252386 370
rect 251498 0 251558 310
rect 252234 0 252294 310
rect 252970 0 253030 443
rect 253703 372 253769 373
rect 253703 308 253704 372
rect 253768 308 253769 372
rect 253703 307 253769 308
rect 253706 0 253766 307
rect 254442 0 254502 579
rect 255178 0 255238 579
rect 255914 0 255974 582
rect 256742 370 256802 1531
rect 257475 1460 257541 1461
rect 257475 1396 257476 1460
rect 257540 1396 257541 1460
rect 257475 1395 257541 1396
rect 257478 370 257538 1395
rect 258119 644 258185 645
rect 258119 580 258120 644
rect 258184 580 258185 644
rect 258950 642 259010 3163
rect 259683 2820 259749 2821
rect 259683 2756 259684 2820
rect 259748 2756 259749 2820
rect 259683 2755 259749 2756
rect 260419 2820 260485 2821
rect 260419 2756 260420 2820
rect 260484 2756 260485 2820
rect 260419 2755 260485 2756
rect 261891 2820 261957 2821
rect 261891 2756 261892 2820
rect 261956 2756 261957 2820
rect 261891 2755 261957 2756
rect 259686 642 259746 2755
rect 260422 642 260482 2755
rect 258119 579 258185 580
rect 258858 582 259010 642
rect 259594 582 259746 642
rect 260330 582 260482 642
rect 261063 644 261129 645
rect 256650 310 256802 370
rect 257386 310 257538 370
rect 256650 0 256710 310
rect 257386 0 257446 310
rect 258122 0 258182 579
rect 258858 0 258918 582
rect 259594 0 259654 582
rect 260330 0 260390 582
rect 261063 580 261064 644
rect 261128 580 261129 644
rect 261894 642 261954 2755
rect 266310 1053 266370 5747
rect 267598 2141 267658 9419
rect 267782 7717 267842 10238
rect 267779 7716 267845 7717
rect 267779 7652 267780 7716
rect 267844 7652 267845 7716
rect 267779 7651 267845 7652
rect 268518 6221 268578 10238
rect 268515 6220 268581 6221
rect 268515 6156 268516 6220
rect 268580 6156 268581 6220
rect 268515 6155 268581 6156
rect 269254 5677 269314 10238
rect 269990 6221 270050 10238
rect 270542 10238 270694 10298
rect 271094 10238 271430 10298
rect 269987 6220 270053 6221
rect 269987 6156 269988 6220
rect 270052 6156 270053 6220
rect 269987 6155 270053 6156
rect 270542 5677 270602 10238
rect 271094 6357 271154 10238
rect 271331 9824 271651 9840
rect 271331 9760 271339 9824
rect 271403 9760 271419 9824
rect 271483 9760 271499 9824
rect 271563 9760 271579 9824
rect 271643 9760 271651 9824
rect 271331 8736 271651 9760
rect 271331 8672 271339 8736
rect 271403 8672 271419 8736
rect 271483 8672 271499 8736
rect 271563 8672 271579 8736
rect 271643 8672 271651 8736
rect 271331 7648 271651 8672
rect 271331 7584 271339 7648
rect 271403 7584 271419 7648
rect 271483 7584 271499 7648
rect 271563 7584 271579 7648
rect 271643 7584 271651 7648
rect 271331 6560 271651 7584
rect 271331 6496 271339 6560
rect 271403 6496 271419 6560
rect 271483 6496 271499 6560
rect 271563 6496 271579 6560
rect 271643 6496 271651 6560
rect 271091 6356 271157 6357
rect 271091 6292 271092 6356
rect 271156 6292 271157 6356
rect 271091 6291 271157 6292
rect 269251 5676 269317 5677
rect 269251 5612 269252 5676
rect 269316 5612 269317 5676
rect 269251 5611 269317 5612
rect 270539 5676 270605 5677
rect 270539 5612 270540 5676
rect 270604 5612 270605 5676
rect 270539 5611 270605 5612
rect 271331 5472 271651 6496
rect 271331 5408 271339 5472
rect 271403 5408 271419 5472
rect 271483 5408 271499 5472
rect 271563 5408 271579 5472
rect 271643 5408 271651 5472
rect 271331 4384 271651 5408
rect 271331 4320 271339 4384
rect 271403 4320 271419 4384
rect 271483 4320 271499 4384
rect 271563 4320 271579 4384
rect 271643 4320 271651 4384
rect 271331 3296 271651 4320
rect 271331 3232 271339 3296
rect 271403 3232 271419 3296
rect 271483 3232 271499 3296
rect 271563 3232 271579 3296
rect 271643 3232 271651 3296
rect 271091 2820 271157 2821
rect 271091 2756 271092 2820
rect 271156 2756 271157 2820
rect 271091 2755 271157 2756
rect 267595 2140 267661 2141
rect 267595 2076 267596 2140
rect 267660 2076 267661 2140
rect 267595 2075 267661 2076
rect 266307 1052 266373 1053
rect 266307 988 266308 1052
rect 266372 988 266373 1052
rect 266307 987 266373 988
rect 261063 579 261129 580
rect 261802 582 261954 642
rect 262535 644 262601 645
rect 261066 0 261126 579
rect 261802 0 261862 582
rect 262535 580 262536 644
rect 262600 580 262601 644
rect 262535 579 262601 580
rect 263271 644 263337 645
rect 263271 580 263272 644
rect 263336 580 263337 644
rect 263271 579 263337 580
rect 264007 644 264073 645
rect 264007 580 264008 644
rect 264072 580 264073 644
rect 264007 579 264073 580
rect 264743 644 264809 645
rect 264743 580 264744 644
rect 264808 580 264809 644
rect 264743 579 264809 580
rect 265479 644 265545 645
rect 265479 580 265480 644
rect 265544 580 265545 644
rect 265479 579 265545 580
rect 266215 644 266281 645
rect 266215 580 266216 644
rect 266280 580 266281 644
rect 266215 579 266281 580
rect 266951 644 267017 645
rect 266951 580 266952 644
rect 267016 580 267017 644
rect 266951 579 267017 580
rect 267687 644 267753 645
rect 267687 580 267688 644
rect 267752 580 267753 644
rect 267687 579 267753 580
rect 268423 644 268489 645
rect 268423 580 268424 644
rect 268488 580 268489 644
rect 268423 579 268489 580
rect 269159 644 269225 645
rect 269159 580 269160 644
rect 269224 580 269225 644
rect 269159 579 269225 580
rect 270631 644 270697 645
rect 270631 580 270632 644
rect 270696 580 270697 644
rect 271094 642 271154 2755
rect 271331 2208 271651 3232
rect 271331 2144 271339 2208
rect 271403 2144 271419 2208
rect 271483 2144 271499 2208
rect 271563 2144 271579 2208
rect 271643 2144 271651 2208
rect 271331 1120 271651 2144
rect 271331 1056 271339 1120
rect 271403 1056 271419 1120
rect 271483 1056 271499 1120
rect 271563 1056 271579 1120
rect 271643 1056 271651 1120
rect 271331 1040 271651 1056
rect 271094 582 271430 642
rect 270631 579 270697 580
rect 262538 0 262598 579
rect 263274 0 263334 579
rect 264010 0 264070 579
rect 264746 0 264806 579
rect 265482 0 265542 579
rect 266218 0 266278 579
rect 266954 0 267014 579
rect 267690 0 267750 579
rect 268426 0 268486 579
rect 269162 0 269222 579
rect 269895 372 269961 373
rect 269895 308 269896 372
rect 269960 308 269961 372
rect 269895 307 269961 308
rect 269898 0 269958 307
rect 270634 0 270694 579
rect 271370 0 271430 582
use sky130_fd_sc_hd__inv_2  _0303_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 270756 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0304_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 270388 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0305_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 256404 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0306_
timestamp 1676037725
transform 1 0 263672 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0307_
timestamp 1676037725
transform 1 0 270756 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0308_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 269652 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0309_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 255576 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0310_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 268732 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o221ai_4  _0311_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 269100 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  _0312_
timestamp 1676037725
transform 1 0 254288 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0313_
timestamp 1676037725
transform 1 0 269100 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0314_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 269376 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _0315_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 269560 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0316_
timestamp 1676037725
transform 1 0 255024 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__nor4_1  _0317_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 252540 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0318_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 254196 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0319_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 255668 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0320_
timestamp 1676037725
transform 1 0 254104 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0321_
timestamp 1676037725
transform 1 0 258244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0322_
timestamp 1676037725
transform 1 0 252816 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0323_
timestamp 1676037725
transform 1 0 254656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0324_
timestamp 1676037725
transform 1 0 255300 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0325_
timestamp 1676037725
transform 1 0 253644 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0326_
timestamp 1676037725
transform 1 0 258704 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0327_
timestamp 1676037725
transform 1 0 257140 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0328_
timestamp 1676037725
transform 1 0 258704 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0329_
timestamp 1676037725
transform 1 0 257692 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0330_
timestamp 1676037725
transform 1 0 257324 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0331_
timestamp 1676037725
transform 1 0 258796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0332_
timestamp 1676037725
transform 1 0 256220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0333_
timestamp 1676037725
transform 1 0 256404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0334_
timestamp 1676037725
transform 1 0 257416 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0335_
timestamp 1676037725
transform 1 0 253092 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0336_
timestamp 1676037725
transform 1 0 250976 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0337_
timestamp 1676037725
transform 1 0 250976 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0338_
timestamp 1676037725
transform 1 0 247296 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0339_
timestamp 1676037725
transform 1 0 247572 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0340_
timestamp 1676037725
transform 1 0 246652 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0341_
timestamp 1676037725
transform 1 0 244352 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0342_
timestamp 1676037725
transform 1 0 247756 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0343_
timestamp 1676037725
transform 1 0 247940 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0344_
timestamp 1676037725
transform 1 0 252540 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0345_
timestamp 1676037725
transform 1 0 247112 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0346_
timestamp 1676037725
transform 1 0 251252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0347_
timestamp 1676037725
transform 1 0 252540 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0348_
timestamp 1676037725
transform 1 0 246192 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0349_
timestamp 1676037725
transform 1 0 245916 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0350_
timestamp 1676037725
transform 1 0 245088 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0351_
timestamp 1676037725
transform 1 0 245364 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0352_
timestamp 1676037725
transform 1 0 244168 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0353_
timestamp 1676037725
transform 1 0 250424 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0354_
timestamp 1676037725
transform 1 0 246744 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0355_
timestamp 1676037725
transform 1 0 251712 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0356_
timestamp 1676037725
transform 1 0 243984 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0357_
timestamp 1676037725
transform 1 0 244720 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0358_
timestamp 1676037725
transform 1 0 247296 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0359_
timestamp 1676037725
transform 1 0 245272 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0360_
timestamp 1676037725
transform 1 0 248860 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0361_
timestamp 1676037725
transform 1 0 249136 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0362_
timestamp 1676037725
transform 1 0 249596 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0363_
timestamp 1676037725
transform 1 0 250516 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0364_
timestamp 1676037725
transform 1 0 259256 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0365_
timestamp 1676037725
transform 1 0 259624 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0366_
timestamp 1676037725
transform 1 0 247664 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0367_
timestamp 1676037725
transform 1 0 249780 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0368_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 116380 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0369_
timestamp 1676037725
transform 1 0 117300 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0370_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 139656 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0371_
timestamp 1676037725
transform 1 0 111320 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0372_
timestamp 1676037725
transform 1 0 132756 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0373_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 136068 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0374_
timestamp 1676037725
transform 1 0 127604 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  _0375_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 144072 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__or3_1  _0376_
timestamp 1676037725
transform 1 0 113436 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0377_
timestamp 1676037725
transform 1 0 112148 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0378_
timestamp 1676037725
transform 1 0 114080 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0379_
timestamp 1676037725
transform 1 0 113160 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0380_
timestamp 1676037725
transform 1 0 114264 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0381_
timestamp 1676037725
transform 1 0 112792 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0382_
timestamp 1676037725
transform 1 0 113804 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0383_
timestamp 1676037725
transform 1 0 113988 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0384_
timestamp 1676037725
transform 1 0 114724 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0385_
timestamp 1676037725
transform 1 0 113436 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0386_
timestamp 1676037725
transform 1 0 102672 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0387_
timestamp 1676037725
transform 1 0 108560 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0388_
timestamp 1676037725
transform 1 0 109572 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0389_
timestamp 1676037725
transform 1 0 108560 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0390_
timestamp 1676037725
transform 1 0 106260 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0391_
timestamp 1676037725
transform 1 0 108560 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0392_
timestamp 1676037725
transform 1 0 108836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0393_
timestamp 1676037725
transform 1 0 107732 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0394_
timestamp 1676037725
transform 1 0 109112 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0395_
timestamp 1676037725
transform 1 0 102764 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0396_
timestamp 1676037725
transform 1 0 100280 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0397_
timestamp 1676037725
transform 1 0 101108 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0398_
timestamp 1676037725
transform 1 0 101844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0399_
timestamp 1676037725
transform 1 0 101936 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0400_
timestamp 1676037725
transform 1 0 101108 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0401_
timestamp 1676037725
transform 1 0 100924 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0402_
timestamp 1676037725
transform 1 0 102488 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0403_
timestamp 1676037725
transform 1 0 102304 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0404_
timestamp 1676037725
transform 1 0 103132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0405_
timestamp 1676037725
transform 1 0 101844 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0406_
timestamp 1676037725
transform 1 0 103408 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0407_
timestamp 1676037725
transform 1 0 101844 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0408_
timestamp 1676037725
transform 1 0 100464 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0409_
timestamp 1676037725
transform 1 0 112148 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0410_
timestamp 1676037725
transform 1 0 98348 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0411_
timestamp 1676037725
transform 1 0 99268 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0412_
timestamp 1676037725
transform 1 0 96968 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0413_
timestamp 1676037725
transform 1 0 92552 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0414_
timestamp 1676037725
transform 1 0 96692 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0415_
timestamp 1676037725
transform 1 0 92736 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0416_
timestamp 1676037725
transform 1 0 98256 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0417_
timestamp 1676037725
transform 1 0 95128 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0418_
timestamp 1676037725
transform 1 0 97336 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0419_
timestamp 1676037725
transform 1 0 93380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0420_
timestamp 1676037725
transform 1 0 97428 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0421_
timestamp 1676037725
transform 1 0 94484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0422_
timestamp 1676037725
transform 1 0 95772 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0423_
timestamp 1676037725
transform 1 0 95956 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0424_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 117576 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0425_
timestamp 1676037725
transform 1 0 118220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _0426_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 140484 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0427_
timestamp 1676037725
transform 1 0 119876 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _0428_
timestamp 1676037725
transform 1 0 145452 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0429_
timestamp 1676037725
transform 1 0 122452 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0430_
timestamp 1676037725
transform 1 0 122452 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0431_
timestamp 1676037725
transform 1 0 121256 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0432_
timestamp 1676037725
transform 1 0 121624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0433_
timestamp 1676037725
transform 1 0 120428 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0434_
timestamp 1676037725
transform 1 0 122268 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0435_
timestamp 1676037725
transform 1 0 120244 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0436_
timestamp 1676037725
transform 1 0 118680 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0437_
timestamp 1676037725
transform 1 0 120612 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0438_
timestamp 1676037725
transform 1 0 119876 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0439_
timestamp 1676037725
transform 1 0 106996 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0440_
timestamp 1676037725
transform 1 0 106996 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_1  _0441_
timestamp 1676037725
transform 1 0 110216 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0442_
timestamp 1676037725
transform 1 0 111412 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0443_
timestamp 1676037725
transform 1 0 109756 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0444_
timestamp 1676037725
transform 1 0 109572 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0445_
timestamp 1676037725
transform 1 0 110216 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0446_
timestamp 1676037725
transform 1 0 109572 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0447_
timestamp 1676037725
transform 1 0 108468 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0448_
timestamp 1676037725
transform 1 0 111872 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0449_
timestamp 1676037725
transform 1 0 109388 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _0450_
timestamp 1676037725
transform 1 0 108008 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0451_
timestamp 1676037725
transform 1 0 105248 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0452_
timestamp 1676037725
transform 1 0 106996 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0453_
timestamp 1676037725
transform 1 0 107916 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0454_
timestamp 1676037725
transform 1 0 107088 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0455_
timestamp 1676037725
transform 1 0 104604 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0456_
timestamp 1676037725
transform 1 0 105892 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0457_
timestamp 1676037725
transform 1 0 105616 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0458_
timestamp 1676037725
transform 1 0 105892 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0459_
timestamp 1676037725
transform 1 0 106076 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0460_
timestamp 1676037725
transform 1 0 104696 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0461_
timestamp 1676037725
transform 1 0 104972 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0462_
timestamp 1676037725
transform 1 0 121440 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0463_
timestamp 1676037725
transform 1 0 108100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0464_
timestamp 1676037725
transform 1 0 100740 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0465_
timestamp 1676037725
transform 1 0 99636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0466_
timestamp 1676037725
transform 1 0 101292 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0467_
timestamp 1676037725
transform 1 0 99912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0468_
timestamp 1676037725
transform 1 0 99452 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0469_
timestamp 1676037725
transform 1 0 93380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0470_
timestamp 1676037725
transform 1 0 100280 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0471_
timestamp 1676037725
transform 1 0 98440 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0472_
timestamp 1676037725
transform 1 0 99728 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0473_
timestamp 1676037725
transform 1 0 94668 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0474_
timestamp 1676037725
transform 1 0 99820 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0475_
timestamp 1676037725
transform 1 0 97704 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0476_
timestamp 1676037725
transform 1 0 99268 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0477_
timestamp 1676037725
transform 1 0 96692 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0478_
timestamp 1676037725
transform 1 0 168820 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0479_
timestamp 1676037725
transform 1 0 168820 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _0480_
timestamp 1676037725
transform 1 0 148212 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0481_
timestamp 1676037725
transform 1 0 155940 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0482_
timestamp 1676037725
transform 1 0 148212 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0483_
timestamp 1676037725
transform 1 0 154652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0484_
timestamp 1676037725
transform 1 0 147016 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0485_
timestamp 1676037725
transform 1 0 146464 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_1  _0486_
timestamp 1676037725
transform 1 0 149684 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0487_
timestamp 1676037725
transform 1 0 153364 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0488_
timestamp 1676037725
transform 1 0 142140 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _0489_
timestamp 1676037725
transform 1 0 150972 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0490_
timestamp 1676037725
transform 1 0 153364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0491_
timestamp 1676037725
transform 1 0 149960 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0492_
timestamp 1676037725
transform 1 0 154376 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0493_
timestamp 1676037725
transform 1 0 151800 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0494_
timestamp 1676037725
transform 1 0 150052 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0495_
timestamp 1676037725
transform 1 0 150788 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0496_
timestamp 1676037725
transform 1 0 149316 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0497_
timestamp 1676037725
transform 1 0 152260 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0498_
timestamp 1676037725
transform 1 0 150052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0499_
timestamp 1676037725
transform 1 0 151248 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0500_
timestamp 1676037725
transform 1 0 153088 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0501_
timestamp 1676037725
transform 1 0 149132 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0502_
timestamp 1676037725
transform 1 0 153732 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0503_
timestamp 1676037725
transform 1 0 148948 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0504_
timestamp 1676037725
transform 1 0 152536 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0505_
timestamp 1676037725
transform 1 0 147936 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0506_
timestamp 1676037725
transform 1 0 148212 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0507_
timestamp 1676037725
transform 1 0 141404 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0508_
timestamp 1676037725
transform 1 0 140484 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_1  _0509_
timestamp 1676037725
transform 1 0 143060 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0510_
timestamp 1676037725
transform 1 0 144164 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0511_
timestamp 1676037725
transform 1 0 138644 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _0512_
timestamp 1676037725
transform 1 0 142140 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0513_
timestamp 1676037725
transform 1 0 144808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0514_
timestamp 1676037725
transform 1 0 143152 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0515_
timestamp 1676037725
transform 1 0 144808 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0516_
timestamp 1676037725
transform 1 0 143796 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0517_
timestamp 1676037725
transform 1 0 143060 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0518_
timestamp 1676037725
transform 1 0 142784 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0519_
timestamp 1676037725
transform 1 0 138644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0520_
timestamp 1676037725
transform 1 0 141588 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0521_
timestamp 1676037725
transform 1 0 138184 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0522_
timestamp 1676037725
transform 1 0 141864 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0523_
timestamp 1676037725
transform 1 0 138828 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0524_
timestamp 1676037725
transform 1 0 138368 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0525_
timestamp 1676037725
transform 1 0 138276 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0526_
timestamp 1676037725
transform 1 0 139380 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0527_
timestamp 1676037725
transform 1 0 138920 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0528_
timestamp 1676037725
transform 1 0 139380 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0529_
timestamp 1676037725
transform 1 0 139472 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_4  _0530_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 212704 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  _0531_
timestamp 1676037725
transform 1 0 215464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0532_
timestamp 1676037725
transform 1 0 216568 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0533_
timestamp 1676037725
transform 1 0 215648 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_2  _0534_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 221352 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nand3b_2  _0535_
timestamp 1676037725
transform 1 0 221536 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__nand3b_2  _0536_
timestamp 1676037725
transform 1 0 223376 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nand3b_1  _0537_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 221536 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _0538_
timestamp 1676037725
transform 1 0 220432 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_2  _0539_
timestamp 1676037725
transform 1 0 218132 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nand3b_1  _0540_
timestamp 1676037725
transform 1 0 217764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _0541_
timestamp 1676037725
transform 1 0 216384 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _0542_
timestamp 1676037725
transform 1 0 217764 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _0543_
timestamp 1676037725
transform 1 0 220432 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0544_
timestamp 1676037725
transform 1 0 205712 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0545_
timestamp 1676037725
transform 1 0 209760 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0546_
timestamp 1676037725
transform 1 0 210036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_2  _0547_
timestamp 1676037725
transform 1 0 211232 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nand3b_2  _0548_
timestamp 1676037725
transform 1 0 212520 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nand3b_2  _0549_
timestamp 1676037725
transform 1 0 211324 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nand3b_2  _0550_
timestamp 1676037725
transform 1 0 211416 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nand3b_2  _0551_
timestamp 1676037725
transform 1 0 211232 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__nand3b_2  _0552_
timestamp 1676037725
transform 1 0 210128 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nand3b_2  _0553_
timestamp 1676037725
transform 1 0 208748 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__nand3b_2  _0554_
timestamp 1676037725
transform 1 0 207552 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nand3b_1  _0555_
timestamp 1676037725
transform 1 0 208748 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _0556_
timestamp 1676037725
transform 1 0 206448 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _0557_
timestamp 1676037725
transform 1 0 206448 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _0558_
timestamp 1676037725
transform 1 0 205528 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0559_
timestamp 1676037725
transform 1 0 248676 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0560_
timestamp 1676037725
transform 1 0 248492 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _0561_
timestamp 1676037725
transform 1 0 215740 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _0562_
timestamp 1676037725
transform 1 0 137448 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0563_
timestamp 1676037725
transform 1 0 138920 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0564_
timestamp 1676037725
transform 1 0 113436 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0565_
timestamp 1676037725
transform 1 0 112792 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0566_
timestamp 1676037725
transform 1 0 110216 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0567_
timestamp 1676037725
transform 1 0 111044 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_4  _0568_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 117300 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0569_
timestamp 1676037725
transform 1 0 68724 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0570_
timestamp 1676037725
transform 1 0 136988 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0571_
timestamp 1676037725
transform 1 0 116104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0572_
timestamp 1676037725
transform 1 0 135332 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0573_
timestamp 1676037725
transform 1 0 152168 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_2  _0574_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 115000 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0575_
timestamp 1676037725
transform 1 0 78660 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_2  _0576_
timestamp 1676037725
transform 1 0 115092 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0577_
timestamp 1676037725
transform 1 0 66700 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _0578_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 114908 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0579_
timestamp 1676037725
transform 1 0 76360 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_2  _0580_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 115828 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0581_
timestamp 1676037725
transform 1 0 91908 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0582_
timestamp 1676037725
transform 1 0 118036 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0583_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 116012 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0584_
timestamp 1676037725
transform 1 0 101292 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0585_
timestamp 1676037725
transform 1 0 119600 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0586_
timestamp 1676037725
transform 1 0 120796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0587_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 118588 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0588_
timestamp 1676037725
transform 1 0 119876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0589_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 167624 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0590_
timestamp 1676037725
transform 1 0 167624 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0591_
timestamp 1676037725
transform 1 0 169832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0592_
timestamp 1676037725
transform 1 0 168360 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0593_
timestamp 1676037725
transform 1 0 168544 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0594_
timestamp 1676037725
transform 1 0 189428 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0595_
timestamp 1676037725
transform 1 0 190256 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0596_
timestamp 1676037725
transform 1 0 189152 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0597_
timestamp 1676037725
transform 1 0 190164 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0598_
timestamp 1676037725
transform 1 0 223376 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0599_
timestamp 1676037725
transform 1 0 224572 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0600_
timestamp 1676037725
transform 1 0 217304 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0601_
timestamp 1676037725
transform 1 0 216752 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0602_
timestamp 1676037725
transform 1 0 221444 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0603_
timestamp 1676037725
transform 1 0 216108 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0604_
timestamp 1676037725
transform 1 0 236532 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _0605_
timestamp 1676037725
transform 1 0 216292 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0606_
timestamp 1676037725
transform 1 0 218408 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0643_
timestamp 1676037725
transform 1 0 62928 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0644_
timestamp 1676037725
transform 1 0 62192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0645_
timestamp 1676037725
transform 1 0 61456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0646_
timestamp 1676037725
transform 1 0 60720 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0647_
timestamp 1676037725
transform 1 0 59800 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0648_
timestamp 1676037725
transform 1 0 59248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0649_
timestamp 1676037725
transform 1 0 58052 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0650_
timestamp 1676037725
transform 1 0 57776 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0651_
timestamp 1676037725
transform 1 0 56948 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0652_
timestamp 1676037725
transform 1 0 56212 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0653_
timestamp 1676037725
transform 1 0 55476 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0654_
timestamp 1676037725
transform 1 0 55476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0655_
timestamp 1676037725
transform 1 0 54280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0656_
timestamp 1676037725
transform 1 0 52716 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0657_
timestamp 1676037725
transform 1 0 66056 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0658_
timestamp 1676037725
transform 1 0 65320 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0659_
timestamp 1676037725
transform 1 0 64492 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0660_
timestamp 1676037725
transform 1 0 63756 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0661_
timestamp 1676037725
transform 1 0 63204 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0662_
timestamp 1676037725
transform 1 0 62284 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0663_
timestamp 1676037725
transform 1 0 61548 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0664_
timestamp 1676037725
transform 1 0 60812 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0665_
timestamp 1676037725
transform 1 0 60076 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0666_
timestamp 1676037725
transform 1 0 59340 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0667_
timestamp 1676037725
transform 1 0 58604 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0668_
timestamp 1676037725
transform 1 0 58052 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0669_
timestamp 1676037725
transform 1 0 57132 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0670_
timestamp 1676037725
transform 1 0 56304 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0671_
timestamp 1676037725
transform 1 0 55476 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0672_
timestamp 1676037725
transform 1 0 55476 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0673_
timestamp 1676037725
transform 1 0 53636 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0674_
timestamp 1676037725
transform 1 0 53084 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0675_
timestamp 1676037725
transform 1 0 98624 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0676_
timestamp 1676037725
transform 1 0 101660 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0677_
timestamp 1676037725
transform 1 0 93564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0678_
timestamp 1676037725
transform 1 0 96692 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0679_
timestamp 1676037725
transform 1 0 94116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0680_
timestamp 1676037725
transform 1 0 92828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0681_
timestamp 1676037725
transform 1 0 93288 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0682_
timestamp 1676037725
transform 1 0 92368 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0683_
timestamp 1676037725
transform 1 0 93196 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0684_
timestamp 1676037725
transform 1 0 92552 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0685_
timestamp 1676037725
transform 1 0 91632 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0686_
timestamp 1676037725
transform 1 0 91816 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0687_
timestamp 1676037725
transform 1 0 90712 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0688_
timestamp 1676037725
transform 1 0 90620 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0689_
timestamp 1676037725
transform 1 0 89976 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0690_
timestamp 1676037725
transform 1 0 89332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0691_
timestamp 1676037725
transform 1 0 88136 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0692_
timestamp 1676037725
transform 1 0 88136 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0693_
timestamp 1676037725
transform 1 0 100280 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0694_
timestamp 1676037725
transform 1 0 99636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0695_
timestamp 1676037725
transform 1 0 99268 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0696_
timestamp 1676037725
transform 1 0 98072 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0697_
timestamp 1676037725
transform 1 0 97336 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0698_
timestamp 1676037725
transform 1 0 96692 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0699_
timestamp 1676037725
transform 1 0 95864 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0700_
timestamp 1676037725
transform 1 0 94852 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0701_
timestamp 1676037725
transform 1 0 94392 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0702_
timestamp 1676037725
transform 1 0 93288 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0703_
timestamp 1676037725
transform 1 0 92552 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0704_
timestamp 1676037725
transform 1 0 91540 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0705_
timestamp 1676037725
transform 1 0 91540 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0706_
timestamp 1676037725
transform 1 0 90620 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0707_
timestamp 1676037725
transform 1 0 90160 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0708_
timestamp 1676037725
transform 1 0 89516 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0709_
timestamp 1676037725
transform 1 0 88228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0710_
timestamp 1676037725
transform 1 0 88780 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0711_
timestamp 1676037725
transform 1 0 134320 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0712_
timestamp 1676037725
transform 1 0 133768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0713_
timestamp 1676037725
transform 1 0 133032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0714_
timestamp 1676037725
transform 1 0 131928 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0715_
timestamp 1676037725
transform 1 0 131468 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0716_
timestamp 1676037725
transform 1 0 130640 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0717_
timestamp 1676037725
transform 1 0 130548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0718_
timestamp 1676037725
transform 1 0 128984 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0719_
timestamp 1676037725
transform 1 0 128248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0720_
timestamp 1676037725
transform 1 0 127604 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0721_
timestamp 1676037725
transform 1 0 126776 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0722_
timestamp 1676037725
transform 1 0 126040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0723_
timestamp 1676037725
transform 1 0 125396 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0724_
timestamp 1676037725
transform 1 0 124200 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0725_
timestamp 1676037725
transform 1 0 124016 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0726_
timestamp 1676037725
transform 1 0 123188 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0727_
timestamp 1676037725
transform 1 0 122452 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0728_
timestamp 1676037725
transform 1 0 121624 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0729_
timestamp 1676037725
transform 1 0 133952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0730_
timestamp 1676037725
transform 1 0 133216 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0731_
timestamp 1676037725
transform 1 0 132756 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0732_
timestamp 1676037725
transform 1 0 131928 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0733_
timestamp 1676037725
transform 1 0 131284 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0734_
timestamp 1676037725
transform 1 0 130548 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0735_
timestamp 1676037725
transform 1 0 129352 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0736_
timestamp 1676037725
transform 1 0 129076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0737_
timestamp 1676037725
transform 1 0 128064 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0738_
timestamp 1676037725
transform 1 0 127512 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0739_
timestamp 1676037725
transform 1 0 126776 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0740_
timestamp 1676037725
transform 1 0 126132 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0741_
timestamp 1676037725
transform 1 0 125396 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0742_
timestamp 1676037725
transform 1 0 125028 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0743_
timestamp 1676037725
transform 1 0 123832 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0744_
timestamp 1676037725
transform 1 0 123004 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0745_
timestamp 1676037725
transform 1 0 122176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0746_
timestamp 1676037725
transform 1 0 121532 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0747_
timestamp 1676037725
transform 1 0 168728 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0748_
timestamp 1676037725
transform 1 0 167716 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0749_
timestamp 1676037725
transform 1 0 166612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0750_
timestamp 1676037725
transform 1 0 165784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0751_
timestamp 1676037725
transform 1 0 165048 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0752_
timestamp 1676037725
transform 1 0 164404 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0753_
timestamp 1676037725
transform 1 0 163668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0754_
timestamp 1676037725
transform 1 0 163668 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0755_
timestamp 1676037725
transform 1 0 161920 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0756_
timestamp 1676037725
transform 1 0 161460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0757_
timestamp 1676037725
transform 1 0 161092 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0758_
timestamp 1676037725
transform 1 0 160632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0759_
timestamp 1676037725
transform 1 0 160172 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0760_
timestamp 1676037725
transform 1 0 159160 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0761_
timestamp 1676037725
transform 1 0 158424 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0762_
timestamp 1676037725
transform 1 0 157688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0763_
timestamp 1676037725
transform 1 0 155572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0764_
timestamp 1676037725
transform 1 0 155756 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0765_
timestamp 1676037725
transform 1 0 170016 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0766_
timestamp 1676037725
transform 1 0 168820 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0767_
timestamp 1676037725
transform 1 0 166704 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0768_
timestamp 1676037725
transform 1 0 166612 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0769_
timestamp 1676037725
transform 1 0 165876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0770_
timestamp 1676037725
transform 1 0 165140 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0771_
timestamp 1676037725
transform 1 0 164404 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0772_
timestamp 1676037725
transform 1 0 163668 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0773_
timestamp 1676037725
transform 1 0 162932 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0774_
timestamp 1676037725
transform 1 0 162196 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0775_
timestamp 1676037725
transform 1 0 161460 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0776_
timestamp 1676037725
transform 1 0 160724 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0777_
timestamp 1676037725
transform 1 0 159988 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0778_
timestamp 1676037725
transform 1 0 159252 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0779_
timestamp 1676037725
transform 1 0 158516 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0780_
timestamp 1676037725
transform 1 0 157044 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0781_
timestamp 1676037725
transform 1 0 156492 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0782_
timestamp 1676037725
transform 1 0 155940 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0783_
timestamp 1676037725
transform 1 0 203688 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0784_
timestamp 1676037725
transform 1 0 203964 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0785_
timestamp 1676037725
transform 1 0 201756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0786_
timestamp 1676037725
transform 1 0 201020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0787_
timestamp 1676037725
transform 1 0 200192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0788_
timestamp 1676037725
transform 1 0 199732 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0789_
timestamp 1676037725
transform 1 0 198536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0790_
timestamp 1676037725
transform 1 0 197800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0791_
timestamp 1676037725
transform 1 0 196972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0792_
timestamp 1676037725
transform 1 0 196144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0793_
timestamp 1676037725
transform 1 0 195408 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0794_
timestamp 1676037725
transform 1 0 194672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0795_
timestamp 1676037725
transform 1 0 194580 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0796_
timestamp 1676037725
transform 1 0 193108 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0797_
timestamp 1676037725
transform 1 0 192372 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0798_
timestamp 1676037725
transform 1 0 191820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0799_
timestamp 1676037725
transform 1 0 190900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0800_
timestamp 1676037725
transform 1 0 190348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0801_
timestamp 1676037725
transform 1 0 203044 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0802_
timestamp 1676037725
transform 1 0 202308 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0803_
timestamp 1676037725
transform 1 0 201296 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0804_
timestamp 1676037725
transform 1 0 200560 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0805_
timestamp 1676037725
transform 1 0 199732 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0806_
timestamp 1676037725
transform 1 0 198996 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0807_
timestamp 1676037725
transform 1 0 198904 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0808_
timestamp 1676037725
transform 1 0 198260 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0809_
timestamp 1676037725
transform 1 0 196328 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0810_
timestamp 1676037725
transform 1 0 196052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0811_
timestamp 1676037725
transform 1 0 195316 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0812_
timestamp 1676037725
transform 1 0 194580 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0813_
timestamp 1676037725
transform 1 0 193844 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0814_
timestamp 1676037725
transform 1 0 193108 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0815_
timestamp 1676037725
transform 1 0 192740 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0816_
timestamp 1676037725
transform 1 0 192004 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0817_
timestamp 1676037725
transform 1 0 191084 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0818_
timestamp 1676037725
transform 1 0 190348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0819_
timestamp 1676037725
transform 1 0 236624 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0820_
timestamp 1676037725
transform 1 0 236624 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0821_
timestamp 1676037725
transform 1 0 234968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0822_
timestamp 1676037725
transform 1 0 234416 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0823_
timestamp 1676037725
transform 1 0 233680 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0824_
timestamp 1676037725
transform 1 0 232944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0825_
timestamp 1676037725
transform 1 0 232208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0826_
timestamp 1676037725
transform 1 0 232116 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0827_
timestamp 1676037725
transform 1 0 231380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0828_
timestamp 1676037725
transform 1 0 229816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0829_
timestamp 1676037725
transform 1 0 229264 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0830_
timestamp 1676037725
transform 1 0 228528 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0831_
timestamp 1676037725
transform 1 0 227792 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0832_
timestamp 1676037725
transform 1 0 227240 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0833_
timestamp 1676037725
transform 1 0 226228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0834_
timestamp 1676037725
transform 1 0 225492 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0835_
timestamp 1676037725
transform 1 0 225492 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0836_
timestamp 1676037725
transform 1 0 224020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0837_
timestamp 1676037725
transform 1 0 236624 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0838_
timestamp 1676037725
transform 1 0 235796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0839_
timestamp 1676037725
transform 1 0 234692 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0840_
timestamp 1676037725
transform 1 0 234232 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0841_
timestamp 1676037725
transform 1 0 233220 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0842_
timestamp 1676037725
transform 1 0 232392 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0843_
timestamp 1676037725
transform 1 0 231748 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0844_
timestamp 1676037725
transform 1 0 231472 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0845_
timestamp 1676037725
transform 1 0 230736 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0846_
timestamp 1676037725
transform 1 0 229632 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0847_
timestamp 1676037725
transform 1 0 228988 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0848_
timestamp 1676037725
transform 1 0 228804 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0849_
timestamp 1676037725
transform 1 0 228068 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0850_
timestamp 1676037725
transform 1 0 226780 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0851_
timestamp 1676037725
transform 1 0 226044 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0852_
timestamp 1676037725
transform 1 0 225308 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0853_
timestamp 1676037725
transform 1 0 224480 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0854_
timestamp 1676037725
transform 1 0 223836 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0855_
timestamp 1676037725
transform 1 0 270572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0856_
timestamp 1676037725
transform 1 0 270112 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0857_
timestamp 1676037725
transform 1 0 270112 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0858_
timestamp 1676037725
transform 1 0 268180 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0859_
timestamp 1676037725
transform 1 0 267444 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0860_
timestamp 1676037725
transform 1 0 266708 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0861_
timestamp 1676037725
transform 1 0 266708 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0862_
timestamp 1676037725
transform 1 0 265604 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0863_
timestamp 1676037725
transform 1 0 264868 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0864_
timestamp 1676037725
transform 1 0 264132 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0865_
timestamp 1676037725
transform 1 0 263120 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0866_
timestamp 1676037725
transform 1 0 263120 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0867_
timestamp 1676037725
transform 1 0 262384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0868_
timestamp 1676037725
transform 1 0 262384 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0869_
timestamp 1676037725
transform 1 0 261832 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0870_
timestamp 1676037725
transform 1 0 261096 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0871_
timestamp 1676037725
transform 1 0 260360 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0872_
timestamp 1676037725
transform 1 0 255576 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0873_
timestamp 1676037725
transform 1 0 270020 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0874_
timestamp 1676037725
transform 1 0 270480 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0875_
timestamp 1676037725
transform 1 0 269284 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0876_
timestamp 1676037725
transform 1 0 270296 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0877_
timestamp 1676037725
transform 1 0 265236 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0878_
timestamp 1676037725
transform 1 0 265880 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0879_
timestamp 1676037725
transform 1 0 265972 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0880_
timestamp 1676037725
transform 1 0 266064 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0881_
timestamp 1676037725
transform 1 0 264776 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0882_
timestamp 1676037725
transform 1 0 264132 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0883_
timestamp 1676037725
transform 1 0 263120 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0884_
timestamp 1676037725
transform 1 0 262292 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0885_
timestamp 1676037725
transform 1 0 262108 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0886_
timestamp 1676037725
transform 1 0 261556 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0887_
timestamp 1676037725
transform 1 0 260268 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0888_
timestamp 1676037725
transform 1 0 259716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0889_
timestamp 1676037725
transform 1 0 258980 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0890_
timestamp 1676037725
transform 1 0 258060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0891_
timestamp 1676037725
transform 1 0 33120 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0892_
timestamp 1676037725
transform 1 0 32844 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0893_
timestamp 1676037725
transform 1 0 67068 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0894_
timestamp 1676037725
transform 1 0 66976 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0895_
timestamp 1676037725
transform 1 0 102580 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0896_
timestamp 1676037725
transform 1 0 101016 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0897_
timestamp 1676037725
transform 1 0 135332 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0898_
timestamp 1676037725
transform 1 0 134504 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0899_
timestamp 1676037725
transform 1 0 168820 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0900_
timestamp 1676037725
transform 1 0 169556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0901_
timestamp 1676037725
transform 1 0 203872 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0902_
timestamp 1676037725
transform 1 0 203872 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0903_
timestamp 1676037725
transform 1 0 237360 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0904_
timestamp 1676037725
transform 1 0 236072 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0905_
timestamp 1676037725
transform 1 0 269836 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0906_
timestamp 1676037725
transform 1 0 269836 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0907_
timestamp 1676037725
transform 1 0 32292 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0908_
timestamp 1676037725
transform 1 0 31004 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0909_
timestamp 1676037725
transform 1 0 30268 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0910_
timestamp 1676037725
transform 1 0 29716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0911_
timestamp 1676037725
transform 1 0 28796 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0912_
timestamp 1676037725
transform 1 0 27968 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0913_
timestamp 1676037725
transform 1 0 27416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0914_
timestamp 1676037725
transform 1 0 26312 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0915_
timestamp 1676037725
transform 1 0 25576 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0916_
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0917_
timestamp 1676037725
transform 1 0 23644 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0918_
timestamp 1676037725
transform 1 0 23368 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0919_
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0920_
timestamp 1676037725
transform 1 0 21160 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0921_
timestamp 1676037725
transform 1 0 22080 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0922_
timestamp 1676037725
transform 1 0 23920 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0923_
timestamp 1676037725
transform 1 0 24840 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0924_
timestamp 1676037725
transform 1 0 25760 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0925_
timestamp 1676037725
transform 1 0 32292 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0926_
timestamp 1676037725
transform 1 0 30820 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0927_
timestamp 1676037725
transform 1 0 30176 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0928_
timestamp 1676037725
transform 1 0 28888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0929_
timestamp 1676037725
transform 1 0 28704 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0930_
timestamp 1676037725
transform 1 0 27968 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0931_
timestamp 1676037725
transform 1 0 27232 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0932_
timestamp 1676037725
transform 1 0 27140 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0933_
timestamp 1676037725
transform 1 0 26312 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0934_
timestamp 1676037725
transform 1 0 25024 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0935_
timestamp 1676037725
transform 1 0 23736 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0936_
timestamp 1676037725
transform 1 0 23460 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0937_
timestamp 1676037725
transform 1 0 22724 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0938_
timestamp 1676037725
transform 1 0 20240 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0939_
timestamp 1676037725
transform 1 0 21160 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0940_
timestamp 1676037725
transform 1 0 21712 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0941_
timestamp 1676037725
transform 1 0 22816 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0942_
timestamp 1676037725
transform 1 0 24564 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0943_
timestamp 1676037725
transform 1 0 66792 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0944_
timestamp 1676037725
transform 1 0 65780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0945_
timestamp 1676037725
transform 1 0 64400 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0946_
timestamp 1676037725
transform 1 0 63664 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_8  _0947_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 248676 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0948_
timestamp 1676037725
transform 1 0 253368 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0949_
timestamp 1676037725
transform 1 0 255024 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0950_
timestamp 1676037725
transform 1 0 255116 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0951_
timestamp 1676037725
transform 1 0 256404 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0952_
timestamp 1676037725
transform 1 0 256404 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0953_
timestamp 1676037725
transform 1 0 255484 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0954_
timestamp 1676037725
transform 1 0 255116 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0955_
timestamp 1676037725
transform 1 0 256404 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0956_
timestamp 1676037725
transform 1 0 254012 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0957_
timestamp 1676037725
transform 1 0 244996 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0958_
timestamp 1676037725
transform 1 0 248676 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0959_
timestamp 1676037725
transform 1 0 248768 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0960_
timestamp 1676037725
transform 1 0 250976 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0961_
timestamp 1676037725
transform 1 0 244904 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0962_
timestamp 1676037725
transform 1 0 244812 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0963_
timestamp 1676037725
transform 1 0 251252 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0964_
timestamp 1676037725
transform 1 0 248768 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0965_
timestamp 1676037725
transform 1 0 248676 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0966_
timestamp 1676037725
transform 1 0 246100 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0967_
timestamp 1676037725
transform 1 0 248492 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0968_
timestamp 1676037725
transform 1 0 248676 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0969_
timestamp 1676037725
transform 1 0 259624 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0970_
timestamp 1676037725
transform 1 0 248860 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0971_
timestamp 1676037725
transform 1 0 110768 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0972_
timestamp 1676037725
transform 1 0 116932 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0973_
timestamp 1676037725
transform 1 0 114816 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0974_
timestamp 1676037725
transform 1 0 115000 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0975_
timestamp 1676037725
transform 1 0 114908 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0976_
timestamp 1676037725
transform 1 0 114724 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0977_
timestamp 1676037725
transform 1 0 114908 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0978_
timestamp 1676037725
transform 1 0 109020 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0979_
timestamp 1676037725
transform 1 0 109112 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0980_
timestamp 1676037725
transform 1 0 109572 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0981_
timestamp 1676037725
transform 1 0 109296 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0982_
timestamp 1676037725
transform 1 0 101844 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0983_
timestamp 1676037725
transform 1 0 101844 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0984_
timestamp 1676037725
transform 1 0 101936 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0985_
timestamp 1676037725
transform 1 0 102304 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0986_
timestamp 1676037725
transform 1 0 102028 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0987_
timestamp 1676037725
transform 1 0 99544 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0988_
timestamp 1676037725
transform 1 0 99084 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0989_
timestamp 1676037725
transform 1 0 99268 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0990_
timestamp 1676037725
transform 1 0 96876 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0991_
timestamp 1676037725
transform 1 0 97428 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0992_
timestamp 1676037725
transform 1 0 94300 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0993_
timestamp 1676037725
transform 1 0 96600 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0994_
timestamp 1676037725
transform 1 0 94300 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0995_
timestamp 1676037725
transform 1 0 113712 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0996_
timestamp 1676037725
transform 1 0 117300 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0997_
timestamp 1676037725
transform 1 0 121440 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0998_
timestamp 1676037725
transform 1 0 120704 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0999_
timestamp 1676037725
transform 1 0 120060 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1000_
timestamp 1676037725
transform 1 0 119508 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1001_
timestamp 1676037725
transform 1 0 117484 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1002_
timestamp 1676037725
transform 1 0 111596 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1003_
timestamp 1676037725
transform 1 0 112148 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1004_
timestamp 1676037725
transform 1 0 111780 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1005_
timestamp 1676037725
transform 1 0 112148 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1006_
timestamp 1676037725
transform 1 0 106996 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1007_
timestamp 1676037725
transform 1 0 107180 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1008_
timestamp 1676037725
transform 1 0 107180 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1009_
timestamp 1676037725
transform 1 0 106996 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1010_
timestamp 1676037725
transform 1 0 105708 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1011_
timestamp 1676037725
transform 1 0 104604 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1012_
timestamp 1676037725
transform 1 0 99452 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1013_
timestamp 1676037725
transform 1 0 99268 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1014_
timestamp 1676037725
transform 1 0 97152 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1015_
timestamp 1676037725
transform 1 0 96876 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1016_
timestamp 1676037725
transform 1 0 94576 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1017_
timestamp 1676037725
transform 1 0 97520 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1018_
timestamp 1676037725
transform 1 0 95312 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1019_
timestamp 1676037725
transform 1 0 140576 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1020_
timestamp 1676037725
transform 1 0 168084 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1021_
timestamp 1676037725
transform 1 0 158240 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1022_
timestamp 1676037725
transform 1 0 156124 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1023_
timestamp 1676037725
transform 1 0 155940 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1024_
timestamp 1676037725
transform 1 0 155664 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1025_
timestamp 1676037725
transform 1 0 155940 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1026_
timestamp 1676037725
transform 1 0 153364 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1027_
timestamp 1676037725
transform 1 0 153088 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1028_
timestamp 1676037725
transform 1 0 150788 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1029_
timestamp 1676037725
transform 1 0 150788 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1030_
timestamp 1676037725
transform 1 0 150236 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1031_
timestamp 1676037725
transform 1 0 150880 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1032_
timestamp 1676037725
transform 1 0 148580 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1033_
timestamp 1676037725
transform 1 0 145636 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1034_
timestamp 1676037725
transform 1 0 145360 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1035_
timestamp 1676037725
transform 1 0 145636 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1036_
timestamp 1676037725
transform 1 0 145360 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1037_
timestamp 1676037725
transform 1 0 142876 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1038_
timestamp 1676037725
transform 1 0 143060 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1039_
timestamp 1676037725
transform 1 0 143060 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1040_
timestamp 1676037725
transform 1 0 140484 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1041_
timestamp 1676037725
transform 1 0 140484 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1042_
timestamp 1676037725
transform 1 0 139564 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1043_
timestamp 1676037725
transform 1 0 220340 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1044_
timestamp 1676037725
transform 1 0 222732 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1045_
timestamp 1676037725
transform 1 0 225216 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1046_
timestamp 1676037725
transform 1 0 225216 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1047_
timestamp 1676037725
transform 1 0 225492 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1048_
timestamp 1676037725
transform 1 0 222916 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1049_
timestamp 1676037725
transform 1 0 221076 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1050_
timestamp 1676037725
transform 1 0 220156 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1051_
timestamp 1676037725
transform 1 0 217948 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1052_
timestamp 1676037725
transform 1 0 217396 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1053_
timestamp 1676037725
transform 1 0 218132 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1054_
timestamp 1676037725
transform 1 0 221352 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1055_
timestamp 1676037725
transform 1 0 215188 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1056_
timestamp 1676037725
transform 1 0 214912 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1057_
timestamp 1676037725
transform 1 0 213164 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1058_
timestamp 1676037725
transform 1 0 215188 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1059_
timestamp 1676037725
transform 1 0 212612 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1060_
timestamp 1676037725
transform 1 0 212336 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1061_
timestamp 1676037725
transform 1 0 210036 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1062_
timestamp 1676037725
transform 1 0 208932 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1063_
timestamp 1676037725
transform 1 0 209760 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1064_
timestamp 1676037725
transform 1 0 207460 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1065_
timestamp 1676037725
transform 1 0 207276 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1066_
timestamp 1676037725
transform 1 0 206448 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 66332 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 248124 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 260820 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 158424 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 159528 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 156308 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1676037725
transform 1 0 259716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1676037725
transform 1 0 156124 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1676037725
transform 1 0 257600 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1676037725
transform 1 0 166888 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1676037725
transform 1 0 270020 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1676037725
transform 1 0 269284 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1676037725
transform 1 0 164588 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1676037725
transform 1 0 266064 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1676037725
transform 1 0 165876 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1676037725
transform 1 0 265696 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1676037725
transform 1 0 163208 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1676037725
transform 1 0 265236 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1676037725
transform 1 0 163024 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1676037725
transform 1 0 161644 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1676037725
transform 1 0 264868 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1676037725
transform 1 0 161460 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1676037725
transform 1 0 264868 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1676037725
transform 1 0 260912 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1676037725
transform 1 0 259808 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1676037725
transform 1 0 261096 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1676037725
transform 1 0 263488 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1676037725
transform 1 0 151800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1676037725
transform 1 0 167624 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1676037725
transform 1 0 216016 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1676037725
transform 1 0 51060 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1676037725
transform 1 0 109572 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1676037725
transform 1 0 103776 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1676037725
transform 1 0 96048 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1676037725
transform 1 0 117300 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1676037725
transform 1 0 117668 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 1676037725
transform 1 0 44620 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp 1676037725
transform 1 0 103408 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp 1676037725
transform 1 0 40204 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp 1676037725
transform 1 0 50416 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_41
timestamp 1676037725
transform 1 0 35144 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_42
timestamp 1676037725
transform 1 0 165876 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_43
timestamp 1676037725
transform 1 0 148028 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_44
timestamp 1676037725
transform 1 0 142416 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_45
timestamp 1676037725
transform 1 0 155848 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_46
timestamp 1676037725
transform 1 0 165508 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_47
timestamp 1676037725
transform 1 0 227608 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_48
timestamp 1676037725
transform 1 0 225032 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_49
timestamp 1676037725
transform 1 0 212428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_50
timestamp 1676037725
transform 1 0 209392 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_51
timestamp 1676037725
transform 1 0 208564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_52
timestamp 1676037725
transform 1 0 224848 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_53
timestamp 1676037725
transform 1 0 214544 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_54
timestamp 1676037725
transform 1 0 40940 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_55
timestamp 1676037725
transform 1 0 39652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_56
timestamp 1676037725
transform 1 0 49588 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_57
timestamp 1676037725
transform 1 0 111504 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_58
timestamp 1676037725
transform 1 0 105248 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_59
timestamp 1676037725
transform 1 0 53452 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_60
timestamp 1676037725
transform 1 0 53636 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_61
timestamp 1676037725
transform 1 0 30636 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_62
timestamp 1676037725
transform 1 0 64676 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_63
timestamp 1676037725
transform 1 0 94852 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_64
timestamp 1676037725
transform 1 0 24932 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_65
timestamp 1676037725
transform 1 0 53636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_66
timestamp 1676037725
transform 1 0 88504 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_67
timestamp 1676037725
transform 1 0 190532 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_68
timestamp 1676037725
transform 1 0 224388 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_69
timestamp 1676037725
transform 1 0 20792 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_70
timestamp 1676037725
transform 1 0 54188 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_71
timestamp 1676037725
transform 1 0 89332 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_72
timestamp 1676037725
transform 1 0 123188 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_73
timestamp 1676037725
transform 1 0 23736 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_74
timestamp 1676037725
transform 1 0 54280 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_75
timestamp 1676037725
transform 1 0 89516 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_76
timestamp 1676037725
transform 1 0 31372 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_77
timestamp 1676037725
transform 1 0 66700 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_78
timestamp 1676037725
transform 1 0 99820 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_79
timestamp 1676037725
transform 1 0 133308 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_80
timestamp 1676037725
transform 1 0 167992 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_81
timestamp 1676037725
transform 1 0 190348 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_82
timestamp 1676037725
transform 1 0 216384 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_83
timestamp 1676037725
transform 1 0 215740 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_84
timestamp 1676037725
transform 1 0 188784 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_85
timestamp 1676037725
transform 1 0 188784 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_86
timestamp 1676037725
transform 1 0 217028 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_87
timestamp 1676037725
transform 1 0 215924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_88
timestamp 1676037725
transform 1 0 248032 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_89
timestamp 1676037725
transform 1 0 259256 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_90
timestamp 1676037725
transform 1 0 262660 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_91
timestamp 1676037725
transform 1 0 117116 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_92
timestamp 1676037725
transform 1 0 103132 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_93
timestamp 1676037725
transform 1 0 213072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_94
timestamp 1676037725
transform 1 0 219972 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_95
timestamp 1676037725
transform 1 0 47932 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_96
timestamp 1676037725
transform 1 0 189980 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_97
timestamp 1676037725
transform 1 0 24288 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_98
timestamp 1676037725
transform 1 0 58512 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_99
timestamp 1676037725
transform 1 0 92920 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_100
timestamp 1676037725
transform 1 0 25116 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_101
timestamp 1676037725
transform 1 0 61272 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_102
timestamp 1676037725
transform 1 0 95588 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_103
timestamp 1676037725
transform 1 0 25760 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_104
timestamp 1676037725
transform 1 0 61640 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_105
timestamp 1676037725
transform 1 0 95956 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_106
timestamp 1676037725
transform 1 0 121072 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_107
timestamp 1676037725
transform 1 0 190164 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_108
timestamp 1676037725
transform 1 0 223376 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_109
timestamp 1676037725
transform 1 0 22724 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_110
timestamp 1676037725
transform 1 0 53268 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_111
timestamp 1676037725
transform 1 0 192464 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_112
timestamp 1676037725
transform 1 0 226044 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_113
timestamp 1676037725
transform 1 0 262292 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_114
timestamp 1676037725
transform 1 0 39284 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_115
timestamp 1676037725
transform 1 0 51428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_116
timestamp 1676037725
transform 1 0 36800 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_117
timestamp 1676037725
transform 1 0 127880 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_118
timestamp 1676037725
transform 1 0 128616 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_119
timestamp 1676037725
transform 1 0 130824 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_120
timestamp 1676037725
transform 1 0 26588 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_121
timestamp 1676037725
transform 1 0 61456 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_122
timestamp 1676037725
transform 1 0 95404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_123
timestamp 1676037725
transform 1 0 122728 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_124
timestamp 1676037725
transform 1 0 21620 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_125
timestamp 1676037725
transform 1 0 56580 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_126
timestamp 1676037725
transform 1 0 91172 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_127
timestamp 1676037725
transform 1 0 124660 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_128
timestamp 1676037725
transform 1 0 195224 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_129
timestamp 1676037725
transform 1 0 23276 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_130
timestamp 1676037725
transform 1 0 57500 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[0\].cell0_I openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 51796 0 1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[1\].cell0_I
timestamp 1676037725
transform 1 0 50784 0 -1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[2\].cell0_I
timestamp 1676037725
transform 1 0 50324 0 -1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[3\].cell0_I
timestamp 1676037725
transform 1 0 50324 0 1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[4\].cell0_I
timestamp 1676037725
transform 1 0 48300 0 -1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[5\].cell0_I
timestamp 1676037725
transform 1 0 48024 0 1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[6\].cell0_I
timestamp 1676037725
transform 1 0 47748 0 -1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[7\].cell0_I
timestamp 1676037725
transform 1 0 46552 0 1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[8\].cell0_I
timestamp 1676037725
transform 1 0 45632 0 -1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[9\].cell0_I
timestamp 1676037725
transform 1 0 45172 0 1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[10\].cell0_I
timestamp 1676037725
transform 1 0 44252 0 -1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[11\].cell0_I
timestamp 1676037725
transform 1 0 43056 0 1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[12\].cell0_I
timestamp 1676037725
transform 1 0 42780 0 -1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[13\].cell0_I
timestamp 1676037725
transform 1 0 42044 0 1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[14\].cell0_I
timestamp 1676037725
transform 1 0 41308 0 1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[15\].cell0_I
timestamp 1676037725
transform 1 0 40572 0 1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[16\].cell0_I
timestamp 1676037725
transform 1 0 40020 0 1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[17\].cell0_I
timestamp 1676037725
transform 1 0 38916 0 -1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[18\].cell0_I
timestamp 1676037725
transform 1 0 37904 0 1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[19\].cell0_I
timestamp 1676037725
transform 1 0 37444 0 -1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[20\].cell0_I
timestamp 1676037725
transform 1 0 37444 0 -1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[21\].cell0_I
timestamp 1676037725
transform 1 0 36156 0 1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[22\].cell0_I
timestamp 1676037725
transform 1 0 35328 0 -1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[23\].cell0_I
timestamp 1676037725
transform 1 0 35512 0 1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  col\[0\].zbuf_bot_ena_I.genblk1.cell0_I_536 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32292 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_ena_I.genblk1.cell0_I openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31832 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 32292 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 31004 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 29992 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 29348 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 28520 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 27692 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 27140 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 25852 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 25024 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 24380 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 23368 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 22816 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 22632 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 22540 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 22080 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 23092 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 23644 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 25300 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 32752 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[0\].zbuf_top_ena_I.genblk1.cell0_I_537
timestamp 1676037725
transform 1 0 32844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 31740 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 30728 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 29992 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 29440 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 28612 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 27784 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 26956 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 26128 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 25484 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 24656 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 23644 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 22632 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 21988 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 22356 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 21988 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 20976 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 23276 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 24472 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[1\].zbuf_bot_ena_I.genblk1.cell0_I_538
timestamp 1676037725
transform 1 0 66332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 66240 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 65964 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 65044 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 64032 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 63388 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 62284 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 62008 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 61272 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 60444 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 59616 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 58788 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 58328 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 57132 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 56304 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 55476 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 54648 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 53636 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 54280 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 54004 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[1\].zbuf_top_ena_I.genblk1.cell0_I_539
timestamp 1676037725
transform 1 0 67712 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 66884 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 66056 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 64860 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 64032 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 63204 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 62376 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 62192 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 61824 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 60628 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 59708 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 58880 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 57868 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 56856 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 56948 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 56212 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 55476 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 54556 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 54464 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 54280 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[0\].cell0_I openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 111872 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[1\].cell0_I
timestamp 1676037725
transform 1 0 115000 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[2\].cell0_I
timestamp 1676037725
transform 1 0 117760 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[3\].cell0_I
timestamp 1676037725
transform 1 0 117484 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[4\].cell0_I
timestamp 1676037725
transform 1 0 117024 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[5\].cell0_I
timestamp 1676037725
transform 1 0 115000 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[6\].cell0_I
timestamp 1676037725
transform 1 0 114908 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[7\].cell0_I
timestamp 1676037725
transform 1 0 109756 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[8\].cell0_I
timestamp 1676037725
transform 1 0 110676 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[9\].cell0_I
timestamp 1676037725
transform 1 0 109756 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[10\].cell0_I
timestamp 1676037725
transform 1 0 112148 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[11\].cell0_I
timestamp 1676037725
transform 1 0 107180 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[12\].cell0_I
timestamp 1676037725
transform 1 0 104880 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[13\].cell0_I
timestamp 1676037725
transform 1 0 104604 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[14\].cell0_I
timestamp 1676037725
transform 1 0 104420 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[15\].cell0_I
timestamp 1676037725
transform 1 0 103500 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[16\].cell0_I
timestamp 1676037725
transform 1 0 99636 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[17\].cell0_I
timestamp 1676037725
transform 1 0 96876 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[18\].cell0_I
timestamp 1676037725
transform 1 0 96692 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[19\].cell0_I
timestamp 1676037725
transform 1 0 94300 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[20\].cell0_I
timestamp 1676037725
transform 1 0 93932 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[21\].cell0_I
timestamp 1676037725
transform 1 0 91540 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[22\].cell0_I
timestamp 1676037725
transform 1 0 94760 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[23\].cell0_I
timestamp 1676037725
transform 1 0 91724 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  col\[2\].zbuf_bot_ena_I.genblk1.cell0_I_540
timestamp 1676037725
transform 1 0 97796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 96048 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 99176 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 95220 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 95404 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 96048 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 94208 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 94944 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 94852 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 94116 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 93196 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 93104 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 92368 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 91540 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 90712 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 90528 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 89884 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 88872 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 89056 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 88872 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[2\].zbuf_top_ena_I.genblk1.cell0_I_541
timestamp 1676037725
transform 1 0 101936 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 100464 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 100188 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 99176 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 98532 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 97704 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 96876 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 96508 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 95772 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 94944 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 94116 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 93288 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 93012 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 92276 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 91540 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 90620 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 89792 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 89700 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 88964 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 89148 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[3\].zbuf_bot_ena_I.genblk1.cell0_I_542
timestamp 1676037725
transform 1 0 135332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 134596 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 134136 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 133308 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 133124 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 132296 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 131376 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 130456 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 129720 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 128892 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 127972 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 127144 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 126316 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 126132 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 125396 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 124752 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 123924 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 123096 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 122084 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 121440 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 134136 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[3\].zbuf_top_ena_I.genblk1.cell0_I_543
timestamp 1676037725
transform 1 0 134228 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 133676 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 132664 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 132664 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 131836 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 131008 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 130180 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 130180 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 128984 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 128248 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 127604 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 126684 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 125856 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 125028 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 124016 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 123372 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 122544 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 121532 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 121256 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_2  col\[4\].genblk1.mux4_I\[0\].cell0_I
timestamp 1676037725
transform 1 0 156216 0 1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[1\].cell0_I
timestamp 1676037725
transform 1 0 166244 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[2\].cell0_I
timestamp 1676037725
transform 1 0 158516 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[3\].cell0_I
timestamp 1676037725
transform 1 0 155664 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[4\].cell0_I
timestamp 1676037725
transform 1 0 153732 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[5\].cell0_I
timestamp 1676037725
transform 1 0 153180 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[6\].cell0_I
timestamp 1676037725
transform 1 0 153364 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[7\].cell0_I
timestamp 1676037725
transform 1 0 150972 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[8\].cell0_I
timestamp 1676037725
transform 1 0 150788 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[9\].cell0_I
timestamp 1676037725
transform 1 0 148948 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[10\].cell0_I
timestamp 1676037725
transform 1 0 148396 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[11\].cell0_I
timestamp 1676037725
transform 1 0 150788 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[12\].cell0_I
timestamp 1676037725
transform 1 0 148212 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[13\].cell0_I
timestamp 1676037725
transform 1 0 147936 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[14\].cell0_I
timestamp 1676037725
transform 1 0 145636 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[15\].cell0_I
timestamp 1676037725
transform 1 0 144440 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[16\].cell0_I
timestamp 1676037725
transform 1 0 145636 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[17\].cell0_I
timestamp 1676037725
transform 1 0 143060 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[18\].cell0_I
timestamp 1676037725
transform 1 0 142784 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[19\].cell0_I
timestamp 1676037725
transform 1 0 140300 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[20\].cell0_I
timestamp 1676037725
transform 1 0 140484 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[21\].cell0_I
timestamp 1676037725
transform 1 0 139288 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[22\].cell0_I
timestamp 1676037725
transform 1 0 140484 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[23\].cell0_I
timestamp 1676037725
transform 1 0 138184 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  col\[4\].zbuf_bot_ena_I.genblk1.cell0_I_544
timestamp 1676037725
transform 1 0 167900 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 167808 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 167900 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 166888 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 167072 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 166244 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 165232 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 164404 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 163576 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 162656 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 162748 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 161920 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 161092 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 159804 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 159344 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 159896 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 159068 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 158516 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 157228 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 156400 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[4\].zbuf_top_ena_I.genblk1.cell0_I_545
timestamp 1676037725
transform 1 0 169924 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 168820 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 167808 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 167256 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 166428 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 166244 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 165324 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 164496 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 163668 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 162748 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 161920 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 161092 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 161000 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 159988 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 158792 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 157780 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 157228 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 156676 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 156952 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 156124 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[5\].zbuf_bot_ena_I.genblk1.cell0_I_546
timestamp 1676037725
transform 1 0 203136 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 203044 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 202860 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 203136 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 202308 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 201296 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 201020 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 200192 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 199364 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 197892 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 197156 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 196236 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 196144 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 195316 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 194488 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 193660 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 192832 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 191820 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 190900 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 190532 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 203136 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[5\].zbuf_top_ena_I.genblk1.cell0_I_547
timestamp 1676037725
transform 1 0 202952 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 203044 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 202308 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 202216 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 201388 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 200560 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 199732 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 198168 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 197432 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 197156 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 196236 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 195224 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 195408 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 194580 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 193200 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 192280 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 192372 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 191544 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 190716 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[0\].cell0_I
timestamp 1676037725
transform 1 0 225216 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[1\].cell0_I
timestamp 1676037725
transform 1 0 223100 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[2\].cell0_I
timestamp 1676037725
transform 1 0 223376 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[3\].cell0_I
timestamp 1676037725
transform 1 0 225492 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[4\].cell0_I
timestamp 1676037725
transform 1 0 222916 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[5\].cell0_I
timestamp 1676037725
transform 1 0 221076 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[6\].cell0_I
timestamp 1676037725
transform 1 0 220064 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[7\].cell0_I
timestamp 1676037725
transform 1 0 218776 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[8\].cell0_I
timestamp 1676037725
transform 1 0 217856 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[9\].cell0_I
timestamp 1676037725
transform 1 0 217764 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[10\].cell0_I
timestamp 1676037725
transform 1 0 217488 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[11\].cell0_I
timestamp 1676037725
transform 1 0 220064 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[12\].cell0_I
timestamp 1676037725
transform 1 0 217764 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[13\].cell0_I
timestamp 1676037725
transform 1 0 215188 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[14\].cell0_I
timestamp 1676037725
transform 1 0 213440 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[15\].cell0_I
timestamp 1676037725
transform 1 0 212796 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[16\].cell0_I
timestamp 1676037725
transform 1 0 214912 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[17\].cell0_I
timestamp 1676037725
transform 1 0 212428 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[18\].cell0_I
timestamp 1676037725
transform 1 0 212612 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[19\].cell0_I
timestamp 1676037725
transform 1 0 210036 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[20\].cell0_I
timestamp 1676037725
transform 1 0 208932 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[21\].cell0_I
timestamp 1676037725
transform 1 0 207000 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[22\].cell0_I
timestamp 1676037725
transform 1 0 208196 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[23\].cell0_I
timestamp 1676037725
transform 1 0 207460 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  col\[6\].zbuf_bot_ena_I.genblk1.cell0_I_548
timestamp 1676037725
transform 1 0 235704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 235796 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 236532 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 235796 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 235704 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 234876 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 234048 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 233220 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 232208 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 231288 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 231380 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 230552 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 229724 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 228896 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 228068 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 226872 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 226412 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 225400 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 224756 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 223744 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 235060 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[6\].zbuf_top_ena_I.genblk1.cell0_I_549
timestamp 1676037725
transform 1 0 235796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 235796 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 234600 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 234416 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 233404 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 233588 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 232760 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 231932 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 230644 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 229908 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 229632 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 228804 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 228068 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 227976 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 227148 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 226320 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 225492 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 224204 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 223376 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[7\].zbuf_bot_ena_I.genblk1.cell0_I_550
timestamp 1676037725
transform 1 0 266616 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 269744 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 269284 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 268916 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 269284 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 268272 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 267444 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 266616 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 265788 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 264960 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 263948 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 264132 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 262936 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 262108 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 261556 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 261556 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 260268 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 261280 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 260268 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 257968 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 268548 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[7\].zbuf_top_ena_I.genblk1.cell0_I_551
timestamp 1676037725
transform 1 0 268548 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 270480 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 267076 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 267444 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 267720 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 266892 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 266524 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 265512 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 265052 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 263948 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 263212 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 263396 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 262384 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 260636 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 261556 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 260636 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 259808 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 258980 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 257876 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  fanout419
timestamp 1676037725
transform 1 0 190716 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout420
timestamp 1676037725
transform 1 0 197616 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout421
timestamp 1676037725
transform 1 0 191084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout422
timestamp 1676037725
transform 1 0 198076 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout423
timestamp 1676037725
transform 1 0 162196 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout424
timestamp 1676037725
transform 1 0 168636 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout425
timestamp 1676037725
transform 1 0 120796 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout426
timestamp 1676037725
transform 1 0 128524 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout427
timestamp 1676037725
transform 1 0 122452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout428
timestamp 1676037725
transform 1 0 128800 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout429
timestamp 1676037725
transform 1 0 94668 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout430
timestamp 1676037725
transform 1 0 100648 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout431
timestamp 1676037725
transform 1 0 60628 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout432
timestamp 1676037725
transform 1 0 66976 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout433
timestamp 1676037725
transform 1 0 60628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout434
timestamp 1676037725
transform 1 0 66516 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout435
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout436
timestamp 1676037725
transform 1 0 33580 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout437
timestamp 1676037725
transform 1 0 258980 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout438
timestamp 1676037725
transform 1 0 264224 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout439
timestamp 1676037725
transform 1 0 259624 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout440
timestamp 1676037725
transform 1 0 264868 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout441
timestamp 1676037725
transform 1 0 223560 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout442
timestamp 1676037725
transform 1 0 230644 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout443
timestamp 1676037725
transform 1 0 162196 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout444
timestamp 1676037725
transform 1 0 168820 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout445
timestamp 1676037725
transform 1 0 92092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout446
timestamp 1676037725
transform 1 0 97796 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout447
timestamp 1676037725
transform 1 0 26128 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout448
timestamp 1676037725
transform 1 0 32660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout449
timestamp 1676037725
transform 1 0 230644 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout450
timestamp 1676037725
transform 1 0 224112 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout451
timestamp 1676037725
transform 1 0 41584 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout452
timestamp 1676037725
transform 1 0 48116 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout453
timestamp 1676037725
transform 1 0 52900 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout454
timestamp 1676037725
transform 1 0 116196 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout455
timestamp 1676037725
transform 1 0 119876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout456
timestamp 1676037725
transform 1 0 105616 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout457
timestamp 1676037725
transform 1 0 152720 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout458
timestamp 1676037725
transform 1 0 153732 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout459
timestamp 1676037725
transform 1 0 167992 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout460
timestamp 1676037725
transform 1 0 223284 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout461
timestamp 1676037725
transform 1 0 225492 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout462
timestamp 1676037725
transform 1 0 225492 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout463 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 225860 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout464
timestamp 1676037725
transform 1 0 42596 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout465
timestamp 1676037725
transform 1 0 47196 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout466
timestamp 1676037725
transform 1 0 52900 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout467
timestamp 1676037725
transform 1 0 109572 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout468
timestamp 1676037725
transform 1 0 117300 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout469
timestamp 1676037725
transform 1 0 119324 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout470
timestamp 1676037725
transform 1 0 151800 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout471
timestamp 1676037725
transform 1 0 152812 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout472
timestamp 1676037725
transform 1 0 169464 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout473
timestamp 1676037725
transform 1 0 224020 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout474
timestamp 1676037725
transform 1 0 225492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout475
timestamp 1676037725
transform 1 0 224296 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout476 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 224388 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout477
timestamp 1676037725
transform 1 0 161828 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout478
timestamp 1676037725
transform 1 0 264132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout479
timestamp 1676037725
transform 1 0 162012 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout480
timestamp 1676037725
transform 1 0 264132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout481
timestamp 1676037725
transform 1 0 163668 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout482
timestamp 1676037725
transform 1 0 265512 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout483
timestamp 1676037725
transform 1 0 163576 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout484
timestamp 1676037725
transform 1 0 265604 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout485
timestamp 1676037725
transform 1 0 164864 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout486
timestamp 1676037725
transform 1 0 266708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout487
timestamp 1676037725
transform 1 0 164956 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout488
timestamp 1676037725
transform 1 0 267628 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout489
timestamp 1676037725
transform 1 0 166060 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout490
timestamp 1676037725
transform 1 0 268548 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout491
timestamp 1676037725
transform 1 0 167256 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout492
timestamp 1676037725
transform 1 0 269468 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout493
timestamp 1676037725
transform 1 0 167256 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout494
timestamp 1676037725
transform 1 0 270388 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout495
timestamp 1676037725
transform 1 0 156492 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout496
timestamp 1676037725
transform 1 0 257968 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout497
timestamp 1676037725
transform 1 0 156676 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout498
timestamp 1676037725
transform 1 0 258980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout499
timestamp 1676037725
transform 1 0 157872 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout500
timestamp 1676037725
transform 1 0 259992 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout501
timestamp 1676037725
transform 1 0 158516 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout502
timestamp 1676037725
transform 1 0 260360 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout503
timestamp 1676037725
transform 1 0 158516 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout504
timestamp 1676037725
transform 1 0 261556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout505
timestamp 1676037725
transform 1 0 158792 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout506
timestamp 1676037725
transform 1 0 261188 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout507
timestamp 1676037725
transform 1 0 159620 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout508
timestamp 1676037725
transform 1 0 262476 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout509
timestamp 1676037725
transform 1 0 160172 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  fanout510
timestamp 1676037725
transform 1 0 262844 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout511
timestamp 1676037725
transform 1 0 168820 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout512
timestamp 1676037725
transform 1 0 268272 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout513
timestamp 1676037725
transform 1 0 265696 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout514
timestamp 1676037725
transform 1 0 265696 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout515
timestamp 1676037725
transform 1 0 261556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout516
timestamp 1676037725
transform 1 0 253000 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_3 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_7 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1748 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_12
timestamp 1676037725
transform 1 0 2208 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3496 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_41 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4876 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_54
timestamp 1676037725
transform 1 0 6072 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1676037725
transform 1 0 6348 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_69
timestamp 1676037725
transform 1 0 7452 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_82
timestamp 1676037725
transform 1 0 8648 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1676037725
transform 1 0 8924 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_97
timestamp 1676037725
transform 1 0 10028 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_110
timestamp 1676037725
transform 1 0 11224 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_113
timestamp 1676037725
transform 1 0 11500 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_125 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12604 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1676037725
transform 1 0 13708 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1676037725
transform 1 0 14076 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_153
timestamp 1676037725
transform 1 0 15180 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_166
timestamp 1676037725
transform 1 0 16376 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_169
timestamp 1676037725
transform 1 0 16652 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_183 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17940 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1676037725
transform 1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1676037725
transform 1 0 19228 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1676037725
transform 1 0 20332 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1676037725
transform 1 0 21436 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_225
timestamp 1676037725
transform 1 0 21804 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_232
timestamp 1676037725
transform 1 0 22448 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_241
timestamp 1676037725
transform 1 0 23276 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_250
timestamp 1676037725
transform 1 0 24104 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_253
timestamp 1676037725
transform 1 0 24380 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_259
timestamp 1676037725
transform 1 0 24932 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_265
timestamp 1676037725
transform 1 0 25484 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_274
timestamp 1676037725
transform 1 0 26312 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_281
timestamp 1676037725
transform 1 0 26956 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_288
timestamp 1676037725
transform 1 0 27600 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_296
timestamp 1676037725
transform 1 0 28336 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_300
timestamp 1676037725
transform 1 0 28704 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1676037725
transform 1 0 29164 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_309
timestamp 1676037725
transform 1 0 29532 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_321
timestamp 1676037725
transform 1 0 30636 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_329
timestamp 1676037725
transform 1 0 31372 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_335
timestamp 1676037725
transform 1 0 31924 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_337
timestamp 1676037725
transform 1 0 32108 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_343
timestamp 1676037725
transform 1 0 32660 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_355
timestamp 1676037725
transform 1 0 33764 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_363
timestamp 1676037725
transform 1 0 34500 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_365
timestamp 1676037725
transform 1 0 34684 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_376
timestamp 1676037725
transform 1 0 35696 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_383
timestamp 1676037725
transform 1 0 36340 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_390
timestamp 1676037725
transform 1 0 36984 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_393
timestamp 1676037725
transform 1 0 37260 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_404
timestamp 1676037725
transform 1 0 38272 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_411
timestamp 1676037725
transform 1 0 38916 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_418
timestamp 1676037725
transform 1 0 39560 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_421
timestamp 1676037725
transform 1 0 39836 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_432
timestamp 1676037725
transform 1 0 40848 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_439
timestamp 1676037725
transform 1 0 41492 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_446
timestamp 1676037725
transform 1 0 42136 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_449
timestamp 1676037725
transform 1 0 42412 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_455
timestamp 1676037725
transform 1 0 42964 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_459
timestamp 1676037725
transform 1 0 43332 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_463
timestamp 1676037725
transform 1 0 43700 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_467
timestamp 1676037725
transform 1 0 44068 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_474
timestamp 1676037725
transform 1 0 44712 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_477
timestamp 1676037725
transform 1 0 44988 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_488
timestamp 1676037725
transform 1 0 46000 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_495
timestamp 1676037725
transform 1 0 46644 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_502
timestamp 1676037725
transform 1 0 47288 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_505
timestamp 1676037725
transform 1 0 47564 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_511
timestamp 1676037725
transform 1 0 48116 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_515
timestamp 1676037725
transform 1 0 48484 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_519
timestamp 1676037725
transform 1 0 48852 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_523
timestamp 1676037725
transform 1 0 49220 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_530
timestamp 1676037725
transform 1 0 49864 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_533
timestamp 1676037725
transform 1 0 50140 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_539
timestamp 1676037725
transform 1 0 50692 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_543
timestamp 1676037725
transform 1 0 51060 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_547
timestamp 1676037725
transform 1 0 51428 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_551
timestamp 1676037725
transform 1 0 51796 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_555
timestamp 1676037725
transform 1 0 52164 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_559
timestamp 1676037725
transform 1 0 52532 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_561
timestamp 1676037725
transform 1 0 52716 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_566
timestamp 1676037725
transform 1 0 53176 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_583
timestamp 1676037725
transform 1 0 54740 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_587
timestamp 1676037725
transform 1 0 55108 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_589
timestamp 1676037725
transform 1 0 55292 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_595
timestamp 1676037725
transform 1 0 55844 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_603
timestamp 1676037725
transform 1 0 56580 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_611
timestamp 1676037725
transform 1 0 57316 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_615
timestamp 1676037725
transform 1 0 57684 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_617
timestamp 1676037725
transform 1 0 57868 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_621
timestamp 1676037725
transform 1 0 58236 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_627
timestamp 1676037725
transform 1 0 58788 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_635
timestamp 1676037725
transform 1 0 59524 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_642
timestamp 1676037725
transform 1 0 60168 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_645
timestamp 1676037725
transform 1 0 60444 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_652
timestamp 1676037725
transform 1 0 61088 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_660
timestamp 1676037725
transform 1 0 61824 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_667
timestamp 1676037725
transform 1 0 62468 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_671
timestamp 1676037725
transform 1 0 62836 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_673
timestamp 1676037725
transform 1 0 63020 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_679
timestamp 1676037725
transform 1 0 63572 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_684
timestamp 1676037725
transform 1 0 64032 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_692
timestamp 1676037725
transform 1 0 64768 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_701
timestamp 1676037725
transform 1 0 65596 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_710
timestamp 1676037725
transform 1 0 66424 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_718
timestamp 1676037725
transform 1 0 67160 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_726
timestamp 1676037725
transform 1 0 67896 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_729
timestamp 1676037725
transform 1 0 68172 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_740
timestamp 1676037725
transform 1 0 69184 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_754
timestamp 1676037725
transform 1 0 70472 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_757
timestamp 1676037725
transform 1 0 70748 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_769
timestamp 1676037725
transform 1 0 71852 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_777
timestamp 1676037725
transform 1 0 72588 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_782
timestamp 1676037725
transform 1 0 73048 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_785
timestamp 1676037725
transform 1 0 73324 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_796
timestamp 1676037725
transform 1 0 74336 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_810
timestamp 1676037725
transform 1 0 75624 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_813
timestamp 1676037725
transform 1 0 75900 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_825
timestamp 1676037725
transform 1 0 77004 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_838
timestamp 1676037725
transform 1 0 78200 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_841
timestamp 1676037725
transform 1 0 78476 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_853
timestamp 1676037725
transform 1 0 79580 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_866
timestamp 1676037725
transform 1 0 80776 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_869
timestamp 1676037725
transform 1 0 81052 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_881
timestamp 1676037725
transform 1 0 82156 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_894
timestamp 1676037725
transform 1 0 83352 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_897
timestamp 1676037725
transform 1 0 83628 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_909
timestamp 1676037725
transform 1 0 84732 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_922
timestamp 1676037725
transform 1 0 85928 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_925
timestamp 1676037725
transform 1 0 86204 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_941
timestamp 1676037725
transform 1 0 87676 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_945
timestamp 1676037725
transform 1 0 88044 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_950
timestamp 1676037725
transform 1 0 88504 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_953
timestamp 1676037725
transform 1 0 88780 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_961
timestamp 1676037725
transform 1 0 89516 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_969
timestamp 1676037725
transform 1 0 90252 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_977
timestamp 1676037725
transform 1 0 90988 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_981
timestamp 1676037725
transform 1 0 91356 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_988
timestamp 1676037725
transform 1 0 92000 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_996
timestamp 1676037725
transform 1 0 92736 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1005
timestamp 1676037725
transform 1 0 93564 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1009
timestamp 1676037725
transform 1 0 93932 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1016
timestamp 1676037725
transform 1 0 94576 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1030
timestamp 1676037725
transform 1 0 95864 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1034
timestamp 1676037725
transform 1 0 96232 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1037
timestamp 1676037725
transform 1 0 96508 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1065
timestamp 1676037725
transform 1 0 99084 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1097
timestamp 1676037725
transform 1 0 102028 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1109
timestamp 1676037725
transform 1 0 103132 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1114
timestamp 1676037725
transform 1 0 103592 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1118
timestamp 1676037725
transform 1 0 103960 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1121
timestamp 1676037725
transform 1 0 104236 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1146
timestamp 1676037725
transform 1 0 106536 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1149
timestamp 1676037725
transform 1 0 106812 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1174
timestamp 1676037725
transform 1 0 109112 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1177
timestamp 1676037725
transform 1 0 109388 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1202
timestamp 1676037725
transform 1 0 111688 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1205
timestamp 1676037725
transform 1 0 111964 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1228
timestamp 1676037725
transform 1 0 114080 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1233
timestamp 1676037725
transform 1 0 114540 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1258
timestamp 1676037725
transform 1 0 116840 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1261
timestamp 1676037725
transform 1 0 117116 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1265
timestamp 1676037725
transform 1 0 117484 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1272
timestamp 1676037725
transform 1 0 118128 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1279
timestamp 1676037725
transform 1 0 118772 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1286
timestamp 1676037725
transform 1 0 119416 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1289
timestamp 1676037725
transform 1 0 119692 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1293
timestamp 1676037725
transform 1 0 120060 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1297
timestamp 1676037725
transform 1 0 120428 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1301
timestamp 1676037725
transform 1 0 120796 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1305
timestamp 1676037725
transform 1 0 121164 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1309
timestamp 1676037725
transform 1 0 121532 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1314
timestamp 1676037725
transform 1 0 121992 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1317
timestamp 1676037725
transform 1 0 122268 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1323
timestamp 1676037725
transform 1 0 122820 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_1331
timestamp 1676037725
transform 1 0 123556 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1337
timestamp 1676037725
transform 1 0 124108 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1342
timestamp 1676037725
transform 1 0 124568 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_1345
timestamp 1676037725
transform 1 0 124844 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1355
timestamp 1676037725
transform 1 0 125764 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1364
timestamp 1676037725
transform 1 0 126592 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1373
timestamp 1676037725
transform 1 0 127420 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1379
timestamp 1676037725
transform 1 0 127972 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1387
timestamp 1676037725
transform 1 0 128708 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_1394
timestamp 1676037725
transform 1 0 129352 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_1401
timestamp 1676037725
transform 1 0 129996 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1407
timestamp 1676037725
transform 1 0 130548 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1412
timestamp 1676037725
transform 1 0 131008 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1420
timestamp 1676037725
transform 1 0 131744 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1426
timestamp 1676037725
transform 1 0 132296 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_1429
timestamp 1676037725
transform 1 0 132572 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1440
timestamp 1676037725
transform 1 0 133584 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1452
timestamp 1676037725
transform 1 0 134688 0 1 1088
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1457
timestamp 1676037725
transform 1 0 135148 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1469
timestamp 1676037725
transform 1 0 136252 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1481
timestamp 1676037725
transform 1 0 137356 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1485
timestamp 1676037725
transform 1 0 137724 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1490
timestamp 1676037725
transform 1 0 138184 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1497
timestamp 1676037725
transform 1 0 138828 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1504
timestamp 1676037725
transform 1 0 139472 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1534
timestamp 1676037725
transform 1 0 142232 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1538
timestamp 1676037725
transform 1 0 142600 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1541
timestamp 1676037725
transform 1 0 142876 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1564
timestamp 1676037725
transform 1 0 144992 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1569
timestamp 1676037725
transform 1 0 145452 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1574
timestamp 1676037725
transform 1 0 145912 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1581
timestamp 1676037725
transform 1 0 146556 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1588
timestamp 1676037725
transform 1 0 147200 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1597
timestamp 1676037725
transform 1 0 148028 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1620
timestamp 1676037725
transform 1 0 150144 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1625
timestamp 1676037725
transform 1 0 150604 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1630
timestamp 1676037725
transform 1 0 151064 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1637
timestamp 1676037725
transform 1 0 151708 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1644
timestamp 1676037725
transform 1 0 152352 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1653
timestamp 1676037725
transform 1 0 153180 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1658
timestamp 1676037725
transform 1 0 153640 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1665
timestamp 1676037725
transform 1 0 154284 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1672
timestamp 1676037725
transform 1 0 154928 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_1681
timestamp 1676037725
transform 1 0 155756 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1687
timestamp 1676037725
transform 1 0 156308 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1693
timestamp 1676037725
transform 1 0 156860 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_1702
timestamp 1676037725
transform 1 0 157688 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1709
timestamp 1676037725
transform 1 0 158332 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1716
timestamp 1676037725
transform 1 0 158976 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1725
timestamp 1676037725
transform 1 0 159804 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1733
timestamp 1676037725
transform 1 0 160540 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1737
timestamp 1676037725
transform 1 0 160908 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1743
timestamp 1676037725
transform 1 0 161460 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1747
timestamp 1676037725
transform 1 0 161828 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1752
timestamp 1676037725
transform 1 0 162288 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1761
timestamp 1676037725
transform 1 0 163116 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1765
timestamp 1676037725
transform 1 0 163484 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1771
timestamp 1676037725
transform 1 0 164036 0 1 1088
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1779
timestamp 1676037725
transform 1 0 164772 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1791
timestamp 1676037725
transform 1 0 165876 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1793
timestamp 1676037725
transform 1 0 166060 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1801
timestamp 1676037725
transform 1 0 166796 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1807
timestamp 1676037725
transform 1 0 167348 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1815
timestamp 1676037725
transform 1 0 168084 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1819
timestamp 1676037725
transform 1 0 168452 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1821
timestamp 1676037725
transform 1 0 168636 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1827
timestamp 1676037725
transform 1 0 169188 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1839
timestamp 1676037725
transform 1 0 170292 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1847
timestamp 1676037725
transform 1 0 171028 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1849
timestamp 1676037725
transform 1 0 171212 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1855
timestamp 1676037725
transform 1 0 171764 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1859
timestamp 1676037725
transform 1 0 172132 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_1870
timestamp 1676037725
transform 1 0 173144 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1877
timestamp 1676037725
transform 1 0 173788 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1889
timestamp 1676037725
transform 1 0 174892 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1901
timestamp 1676037725
transform 1 0 175996 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1905
timestamp 1676037725
transform 1 0 176364 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1917
timestamp 1676037725
transform 1 0 177468 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1929
timestamp 1676037725
transform 1 0 178572 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1933
timestamp 1676037725
transform 1 0 178940 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1945
timestamp 1676037725
transform 1 0 180044 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1957
timestamp 1676037725
transform 1 0 181148 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1961
timestamp 1676037725
transform 1 0 181516 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1973
timestamp 1676037725
transform 1 0 182620 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1985
timestamp 1676037725
transform 1 0 183724 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1989
timestamp 1676037725
transform 1 0 184092 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_2001
timestamp 1676037725
transform 1 0 185196 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_2013
timestamp 1676037725
transform 1 0 186300 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2017
timestamp 1676037725
transform 1 0 186668 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_2029
timestamp 1676037725
transform 1 0 187772 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2035
timestamp 1676037725
transform 1 0 188324 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2039
timestamp 1676037725
transform 1 0 188692 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2043
timestamp 1676037725
transform 1 0 189060 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2045
timestamp 1676037725
transform 1 0 189244 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2057
timestamp 1676037725
transform 1 0 190348 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2061
timestamp 1676037725
transform 1 0 190716 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2068
timestamp 1676037725
transform 1 0 191360 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_2073
timestamp 1676037725
transform 1 0 191820 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2083
timestamp 1676037725
transform 1 0 192740 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2091
timestamp 1676037725
transform 1 0 193476 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2099
timestamp 1676037725
transform 1 0 194212 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2101
timestamp 1676037725
transform 1 0 194396 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2107
timestamp 1676037725
transform 1 0 194948 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2111
timestamp 1676037725
transform 1 0 195316 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2116
timestamp 1676037725
transform 1 0 195776 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2120
timestamp 1676037725
transform 1 0 196144 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2126
timestamp 1676037725
transform 1 0 196696 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2129
timestamp 1676037725
transform 1 0 196972 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2137
timestamp 1676037725
transform 1 0 197708 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_2144
timestamp 1676037725
transform 1 0 198352 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2157
timestamp 1676037725
transform 1 0 199548 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_2163
timestamp 1676037725
transform 1 0 200100 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2175
timestamp 1676037725
transform 1 0 201204 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_2181
timestamp 1676037725
transform 1 0 201756 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2185
timestamp 1676037725
transform 1 0 202124 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2198
timestamp 1676037725
transform 1 0 203320 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_2206
timestamp 1676037725
transform 1 0 204056 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2213
timestamp 1676037725
transform 1 0 204700 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2221
timestamp 1676037725
transform 1 0 205436 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2226
timestamp 1676037725
transform 1 0 205896 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2230
timestamp 1676037725
transform 1 0 206264 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_2234
timestamp 1676037725
transform 1 0 206632 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2241
timestamp 1676037725
transform 1 0 207276 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2246
timestamp 1676037725
transform 1 0 207736 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2253
timestamp 1676037725
transform 1 0 208380 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2260
timestamp 1676037725
transform 1 0 209024 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2266
timestamp 1676037725
transform 1 0 209576 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2269
timestamp 1676037725
transform 1 0 209852 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2292
timestamp 1676037725
transform 1 0 211968 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2318
timestamp 1676037725
transform 1 0 214360 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2322
timestamp 1676037725
transform 1 0 214728 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2325
timestamp 1676037725
transform 1 0 215004 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2348
timestamp 1676037725
transform 1 0 217120 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2353
timestamp 1676037725
transform 1 0 217580 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2361
timestamp 1676037725
transform 1 0 218316 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2368
timestamp 1676037725
transform 1 0 218960 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2375
timestamp 1676037725
transform 1 0 219604 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2379
timestamp 1676037725
transform 1 0 219972 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2381
timestamp 1676037725
transform 1 0 220156 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2386
timestamp 1676037725
transform 1 0 220616 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2394
timestamp 1676037725
transform 1 0 221352 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_2405
timestamp 1676037725
transform 1 0 222364 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2409
timestamp 1676037725
transform 1 0 222732 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2414
timestamp 1676037725
transform 1 0 223192 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2422
timestamp 1676037725
transform 1 0 223928 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2428
timestamp 1676037725
transform 1 0 224480 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2437
timestamp 1676037725
transform 1 0 225308 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2443
timestamp 1676037725
transform 1 0 225860 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2450
timestamp 1676037725
transform 1 0 226504 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2459
timestamp 1676037725
transform 1 0 227332 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2463
timestamp 1676037725
transform 1 0 227700 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_2465
timestamp 1676037725
transform 1 0 227884 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2471
timestamp 1676037725
transform 1 0 228436 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2476
timestamp 1676037725
transform 1 0 228896 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2484
timestamp 1676037725
transform 1 0 229632 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2493
timestamp 1676037725
transform 1 0 230460 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2501
timestamp 1676037725
transform 1 0 231196 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2507
timestamp 1676037725
transform 1 0 231748 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2515
timestamp 1676037725
transform 1 0 232484 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2519
timestamp 1676037725
transform 1 0 232852 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_2521
timestamp 1676037725
transform 1 0 233036 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2527
timestamp 1676037725
transform 1 0 233588 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2532
timestamp 1676037725
transform 1 0 234048 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2540
timestamp 1676037725
transform 1 0 234784 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2549
timestamp 1676037725
transform 1 0 235612 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2556
timestamp 1676037725
transform 1 0 236256 0 1 1088
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_2564
timestamp 1676037725
transform 1 0 236992 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_2577
timestamp 1676037725
transform 1 0 238188 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2589
timestamp 1676037725
transform 1 0 239292 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2593
timestamp 1676037725
transform 1 0 239660 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_2597
timestamp 1676037725
transform 1 0 240028 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2603
timestamp 1676037725
transform 1 0 240580 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2605
timestamp 1676037725
transform 1 0 240764 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_2617
timestamp 1676037725
transform 1 0 241868 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_2629
timestamp 1676037725
transform 1 0 242972 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2633
timestamp 1676037725
transform 1 0 243340 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2645
timestamp 1676037725
transform 1 0 244444 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2653
timestamp 1676037725
transform 1 0 245180 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_2657
timestamp 1676037725
transform 1 0 245548 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2661
timestamp 1676037725
transform 1 0 245916 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_2673
timestamp 1676037725
transform 1 0 247020 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2682
timestamp 1676037725
transform 1 0 247848 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2686
timestamp 1676037725
transform 1 0 248216 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_2689
timestamp 1676037725
transform 1 0 248492 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_2713
timestamp 1676037725
transform 1 0 250700 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2717
timestamp 1676037725
transform 1 0 251068 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2729
timestamp 1676037725
transform 1 0 252172 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2736
timestamp 1676037725
transform 1 0 252816 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2745
timestamp 1676037725
transform 1 0 253644 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2757
timestamp 1676037725
transform 1 0 254748 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2765
timestamp 1676037725
transform 1 0 255484 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2770
timestamp 1676037725
transform 1 0 255944 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2773
timestamp 1676037725
transform 1 0 256220 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_2785
timestamp 1676037725
transform 1 0 257324 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2791
timestamp 1676037725
transform 1 0 257876 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_2797
timestamp 1676037725
transform 1 0 258428 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2801
timestamp 1676037725
transform 1 0 258796 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2813
timestamp 1676037725
transform 1 0 259900 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_2822
timestamp 1676037725
transform 1 0 260728 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2829
timestamp 1676037725
transform 1 0 261372 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2836
timestamp 1676037725
transform 1 0 262016 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2844
timestamp 1676037725
transform 1 0 262752 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2852
timestamp 1676037725
transform 1 0 263488 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2857
timestamp 1676037725
transform 1 0 263948 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2863
timestamp 1676037725
transform 1 0 264500 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2871
timestamp 1676037725
transform 1 0 265236 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2879
timestamp 1676037725
transform 1 0 265972 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2883
timestamp 1676037725
transform 1 0 266340 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2885
timestamp 1676037725
transform 1 0 266524 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2891
timestamp 1676037725
transform 1 0 267076 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2899
timestamp 1676037725
transform 1 0 267812 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2907
timestamp 1676037725
transform 1 0 268548 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2911
timestamp 1676037725
transform 1 0 268916 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2913
timestamp 1676037725
transform 1 0 269100 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2920
timestamp 1676037725
transform 1 0 269744 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2928
timestamp 1676037725
transform 1 0 270480 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_9
timestamp 1676037725
transform 1 0 1932 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_21
timestamp 1676037725
transform 1 0 3036 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_43
timestamp 1676037725
transform 1 0 5060 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 1676037725
transform 1 0 6072 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_75
timestamp 1676037725
transform 1 0 8004 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_89
timestamp 1676037725
transform 1 0 9292 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_103
timestamp 1676037725
transform 1 0 10580 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_121
timestamp 1676037725
transform 1 0 12236 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_129
timestamp 1676037725
transform 1 0 12972 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_151
timestamp 1676037725
transform 1 0 14996 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_155
timestamp 1676037725
transform 1 0 15364 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_166
timestamp 1676037725
transform 1 0 16376 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_185
timestamp 1676037725
transform 1 0 18124 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_197
timestamp 1676037725
transform 1 0 19228 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_209
timestamp 1676037725
transform 1 0 20332 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_217
timestamp 1676037725
transform 1 0 21068 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_222
timestamp 1676037725
transform 1 0 21528 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_233
timestamp 1676037725
transform 1 0 22540 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_244
timestamp 1676037725
transform 1 0 23552 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_254
timestamp 1676037725
transform 1 0 24472 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_264
timestamp 1676037725
transform 1 0 25392 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_274
timestamp 1676037725
transform 1 0 26312 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_294
timestamp 1676037725
transform 1 0 28152 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_303
timestamp 1676037725
transform 1 0 28980 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_312
timestamp 1676037725
transform 1 0 29808 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_319
timestamp 1676037725
transform 1 0 30452 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_323
timestamp 1676037725
transform 1 0 30820 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_330
timestamp 1676037725
transform 1 0 31464 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_344
timestamp 1676037725
transform 1 0 32752 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_352
timestamp 1676037725
transform 1 0 33488 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_364
timestamp 1676037725
transform 1 0 34592 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_371
timestamp 1676037725
transform 1 0 35236 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_383
timestamp 1676037725
transform 1 0 36340 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_399
timestamp 1676037725
transform 1 0 37812 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_403
timestamp 1676037725
transform 1 0 38180 0 -1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_429
timestamp 1676037725
transform 1 0 40572 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_441
timestamp 1676037725
transform 1 0 41676 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_447
timestamp 1676037725
transform 1 0 42228 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_461
timestamp 1676037725
transform 1 0 43516 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_473
timestamp 1676037725
transform 1 0 44620 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_479
timestamp 1676037725
transform 1 0 45172 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_483
timestamp 1676037725
transform 1 0 45540 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_495
timestamp 1676037725
transform 1 0 46644 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_503
timestamp 1676037725
transform 1 0 47380 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_505
timestamp 1676037725
transform 1 0 47564 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_517
timestamp 1676037725
transform 1 0 48668 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_529
timestamp 1676037725
transform 1 0 49772 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_541
timestamp 1676037725
transform 1 0 50876 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_553
timestamp 1676037725
transform 1 0 51980 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_559
timestamp 1676037725
transform 1 0 52532 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_565
timestamp 1676037725
transform 1 0 53084 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_569
timestamp 1676037725
transform 1 0 53452 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_576
timestamp 1676037725
transform 1 0 54096 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_580
timestamp 1676037725
transform 1 0 54464 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_587
timestamp 1676037725
transform 1 0 55108 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_596
timestamp 1676037725
transform 1 0 55936 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_605
timestamp 1676037725
transform 1 0 56764 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_614
timestamp 1676037725
transform 1 0 57592 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_617
timestamp 1676037725
transform 1 0 57868 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_623
timestamp 1676037725
transform 1 0 58420 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_632
timestamp 1676037725
transform 1 0 59248 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_641
timestamp 1676037725
transform 1 0 60076 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_650
timestamp 1676037725
transform 1 0 60904 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_659
timestamp 1676037725
transform 1 0 61732 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_670
timestamp 1676037725
transform 1 0 62744 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_673
timestamp 1676037725
transform 1 0 63020 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_682
timestamp 1676037725
transform 1 0 63848 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_689
timestamp 1676037725
transform 1 0 64492 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_693
timestamp 1676037725
transform 1 0 64860 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_700
timestamp 1676037725
transform 1 0 65504 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_713
timestamp 1676037725
transform 1 0 66700 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_721
timestamp 1676037725
transform 1 0 67436 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_727
timestamp 1676037725
transform 1 0 67988 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_729
timestamp 1676037725
transform 1 0 68172 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_741
timestamp 1676037725
transform 1 0 69276 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_753
timestamp 1676037725
transform 1 0 70380 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_761
timestamp 1676037725
transform 1 0 71116 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_766
timestamp 1676037725
transform 1 0 71576 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_770
timestamp 1676037725
transform 1 0 71944 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_774
timestamp 1676037725
transform 1 0 72312 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_782
timestamp 1676037725
transform 1 0 73048 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_785
timestamp 1676037725
transform 1 0 73324 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_790
timestamp 1676037725
transform 1 0 73784 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_802
timestamp 1676037725
transform 1 0 74888 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_810
timestamp 1676037725
transform 1 0 75624 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_821
timestamp 1676037725
transform 1 0 76636 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_837
timestamp 1676037725
transform 1 0 78108 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_841
timestamp 1676037725
transform 1 0 78476 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_849
timestamp 1676037725
transform 1 0 79212 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_861
timestamp 1676037725
transform 1 0 80316 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_877
timestamp 1676037725
transform 1 0 81788 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_893
timestamp 1676037725
transform 1 0 83260 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_897
timestamp 1676037725
transform 1 0 83628 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_905
timestamp 1676037725
transform 1 0 84364 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_917
timestamp 1676037725
transform 1 0 85468 0 -1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_933
timestamp 1676037725
transform 1 0 86940 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_945
timestamp 1676037725
transform 1 0 88044 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_950
timestamp 1676037725
transform 1 0 88504 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_953
timestamp 1676037725
transform 1 0 88780 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_959
timestamp 1676037725
transform 1 0 89332 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_963
timestamp 1676037725
transform 1 0 89700 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_970
timestamp 1676037725
transform 1 0 90344 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_979
timestamp 1676037725
transform 1 0 91172 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_988
timestamp 1676037725
transform 1 0 92000 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_997
timestamp 1676037725
transform 1 0 92828 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1006
timestamp 1676037725
transform 1 0 93656 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_1009
timestamp 1676037725
transform 1 0 93932 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1017
timestamp 1676037725
transform 1 0 94668 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1021
timestamp 1676037725
transform 1 0 95036 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1028
timestamp 1676037725
transform 1 0 95680 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1037
timestamp 1676037725
transform 1 0 96508 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1062
timestamp 1676037725
transform 1 0 98808 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1065
timestamp 1676037725
transform 1 0 99084 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_1088
timestamp 1676037725
transform 1 0 101200 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_1094
timestamp 1676037725
transform 1 0 101752 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1116
timestamp 1676037725
transform 1 0 103776 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_1121
timestamp 1676037725
transform 1 0 104236 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_1127
timestamp 1676037725
transform 1 0 104788 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1149
timestamp 1676037725
transform 1 0 106812 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1174
timestamp 1676037725
transform 1 0 109112 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1177
timestamp 1676037725
transform 1 0 109388 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_1185
timestamp 1676037725
transform 1 0 110124 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_1212
timestamp 1676037725
transform 1 0 112608 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1223
timestamp 1676037725
transform 1 0 113620 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1230
timestamp 1676037725
transform 1 0 114264 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1233
timestamp 1676037725
transform 1 0 114540 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_1237
timestamp 1676037725
transform 1 0 114908 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1259
timestamp 1676037725
transform 1 0 116932 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1263
timestamp 1676037725
transform 1 0 117300 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1286
timestamp 1676037725
transform 1 0 119416 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1289
timestamp 1676037725
transform 1 0 119692 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1294
timestamp 1676037725
transform 1 0 120152 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_1301
timestamp 1676037725
transform 1 0 120796 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1306
timestamp 1676037725
transform 1 0 121256 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1313
timestamp 1676037725
transform 1 0 121900 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1320
timestamp 1676037725
transform 1 0 122544 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1324
timestamp 1676037725
transform 1 0 122912 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1331
timestamp 1676037725
transform 1 0 123556 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1340
timestamp 1676037725
transform 1 0 124384 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_1345
timestamp 1676037725
transform 1 0 124844 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1356
timestamp 1676037725
transform 1 0 125856 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_1360
timestamp 1676037725
transform 1 0 126224 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1366
timestamp 1676037725
transform 1 0 126776 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1375
timestamp 1676037725
transform 1 0 127604 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1384
timestamp 1676037725
transform 1 0 128432 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1398
timestamp 1676037725
transform 1 0 129720 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1401
timestamp 1676037725
transform 1 0 129996 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_1405
timestamp 1676037725
transform 1 0 130364 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1411
timestamp 1676037725
transform 1 0 130916 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_1415
timestamp 1676037725
transform 1 0 131284 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1421
timestamp 1676037725
transform 1 0 131836 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_1425
timestamp 1676037725
transform 1 0 132204 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_1431
timestamp 1676037725
transform 1 0 132756 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1442
timestamp 1676037725
transform 1 0 133768 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1451
timestamp 1676037725
transform 1 0 134596 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_1455
timestamp 1676037725
transform 1 0 134964 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1457
timestamp 1676037725
transform 1 0 135148 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1463
timestamp 1676037725
transform 1 0 135700 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1475
timestamp 1676037725
transform 1 0 136804 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1487
timestamp 1676037725
transform 1 0 137908 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1494
timestamp 1676037725
transform 1 0 138552 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1501
timestamp 1676037725
transform 1 0 139196 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1508
timestamp 1676037725
transform 1 0 139840 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1513
timestamp 1676037725
transform 1 0 140300 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1536
timestamp 1676037725
transform 1 0 142416 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_1561
timestamp 1676037725
transform 1 0 144716 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_1567
timestamp 1676037725
transform 1 0 145268 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1569
timestamp 1676037725
transform 1 0 145452 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1592
timestamp 1676037725
transform 1 0 147568 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_1617
timestamp 1676037725
transform 1 0 149868 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_1623
timestamp 1676037725
transform 1 0 150420 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1625
timestamp 1676037725
transform 1 0 150604 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1648
timestamp 1676037725
transform 1 0 152720 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1655
timestamp 1676037725
transform 1 0 153364 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1662
timestamp 1676037725
transform 1 0 154008 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1669
timestamp 1676037725
transform 1 0 154652 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1676
timestamp 1676037725
transform 1 0 155296 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1685
timestamp 1676037725
transform 1 0 156124 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1689
timestamp 1676037725
transform 1 0 156492 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1700
timestamp 1676037725
transform 1 0 157504 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1713
timestamp 1676037725
transform 1 0 158700 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1722
timestamp 1676037725
transform 1 0 159528 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1731
timestamp 1676037725
transform 1 0 160356 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_1735
timestamp 1676037725
transform 1 0 160724 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1737
timestamp 1676037725
transform 1 0 160908 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1744
timestamp 1676037725
transform 1 0 161552 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1753
timestamp 1676037725
transform 1 0 162380 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1762
timestamp 1676037725
transform 1 0 163208 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1771
timestamp 1676037725
transform 1 0 164036 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1780
timestamp 1676037725
transform 1 0 164864 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_1789
timestamp 1676037725
transform 1 0 165692 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1793
timestamp 1676037725
transform 1 0 166060 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1800
timestamp 1676037725
transform 1 0 166704 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1809
timestamp 1676037725
transform 1 0 167532 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1818
timestamp 1676037725
transform 1 0 168360 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1826
timestamp 1676037725
transform 1 0 169096 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_1838
timestamp 1676037725
transform 1 0 170200 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1846
timestamp 1676037725
transform 1 0 170936 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1849
timestamp 1676037725
transform 1 0 171212 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_1861
timestamp 1676037725
transform 1 0 172316 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_1867
timestamp 1676037725
transform 1 0 172868 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_1878
timestamp 1676037725
transform 1 0 173880 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_1894
timestamp 1676037725
transform 1 0 175352 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1902
timestamp 1676037725
transform 1 0 176088 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1905
timestamp 1676037725
transform 1 0 176364 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1917
timestamp 1676037725
transform 1 0 177468 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1931
timestamp 1676037725
transform 1 0 178756 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1945
timestamp 1676037725
transform 1 0 180044 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_1957
timestamp 1676037725
transform 1 0 181148 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1961
timestamp 1676037725
transform 1 0 181516 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1973
timestamp 1676037725
transform 1 0 182620 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1987
timestamp 1676037725
transform 1 0 183908 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_2001
timestamp 1676037725
transform 1 0 185196 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_2013
timestamp 1676037725
transform 1 0 186300 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2017
timestamp 1676037725
transform 1 0 186668 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2029
timestamp 1676037725
transform 1 0 187772 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_2043
timestamp 1676037725
transform 1 0 189060 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2057
timestamp 1676037725
transform 1 0 190348 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_2064
timestamp 1676037725
transform 1 0 190992 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2078
timestamp 1676037725
transform 1 0 192280 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2082
timestamp 1676037725
transform 1 0 192648 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2089
timestamp 1676037725
transform 1 0 193292 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2098
timestamp 1676037725
transform 1 0 194120 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2107
timestamp 1676037725
transform 1 0 194948 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2116
timestamp 1676037725
transform 1 0 195776 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_2125
timestamp 1676037725
transform 1 0 196604 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2129
timestamp 1676037725
transform 1 0 196972 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2136
timestamp 1676037725
transform 1 0 197616 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_2140
timestamp 1676037725
transform 1 0 197984 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2151
timestamp 1676037725
transform 1 0 198996 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2160
timestamp 1676037725
transform 1 0 199824 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2169
timestamp 1676037725
transform 1 0 200652 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_2178
timestamp 1676037725
transform 1 0 201480 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2185
timestamp 1676037725
transform 1 0 202124 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2192
timestamp 1676037725
transform 1 0 202768 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2201
timestamp 1676037725
transform 1 0 203596 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_2209
timestamp 1676037725
transform 1 0 204332 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_2221
timestamp 1676037725
transform 1 0 205436 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_2233
timestamp 1676037725
transform 1 0 206540 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_2239
timestamp 1676037725
transform 1 0 207092 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2241
timestamp 1676037725
transform 1 0 207276 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2248
timestamp 1676037725
transform 1 0 207920 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2255
timestamp 1676037725
transform 1 0 208564 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2280
timestamp 1676037725
transform 1 0 210864 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_2293
timestamp 1676037725
transform 1 0 212060 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2297
timestamp 1676037725
transform 1 0 212428 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2320
timestamp 1676037725
transform 1 0 214544 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_2345
timestamp 1676037725
transform 1 0 216844 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_2351
timestamp 1676037725
transform 1 0 217396 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2353
timestamp 1676037725
transform 1 0 217580 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2376
timestamp 1676037725
transform 1 0 219696 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_2401
timestamp 1676037725
transform 1 0 221996 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_2407
timestamp 1676037725
transform 1 0 222548 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2409
timestamp 1676037725
transform 1 0 222732 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2414
timestamp 1676037725
transform 1 0 223192 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2418
timestamp 1676037725
transform 1 0 223560 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2425
timestamp 1676037725
transform 1 0 224204 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2429
timestamp 1676037725
transform 1 0 224572 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2436
timestamp 1676037725
transform 1 0 225216 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2443
timestamp 1676037725
transform 1 0 225860 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2447
timestamp 1676037725
transform 1 0 226228 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2454
timestamp 1676037725
transform 1 0 226872 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2462
timestamp 1676037725
transform 1 0 227608 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2465
timestamp 1676037725
transform 1 0 227884 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2472
timestamp 1676037725
transform 1 0 228528 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2481
timestamp 1676037725
transform 1 0 229356 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2490
timestamp 1676037725
transform 1 0 230184 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2499
timestamp 1676037725
transform 1 0 231012 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2508
timestamp 1676037725
transform 1 0 231840 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_2517
timestamp 1676037725
transform 1 0 232668 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2521
timestamp 1676037725
transform 1 0 233036 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2528
timestamp 1676037725
transform 1 0 233680 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2537
timestamp 1676037725
transform 1 0 234508 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2546
timestamp 1676037725
transform 1 0 235336 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2555
timestamp 1676037725
transform 1 0 236164 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2564
timestamp 1676037725
transform 1 0 236992 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2572
timestamp 1676037725
transform 1 0 237728 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_2577
timestamp 1676037725
transform 1 0 238188 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_2589
timestamp 1676037725
transform 1 0 239292 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_2601
timestamp 1676037725
transform 1 0 240396 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_2609
timestamp 1676037725
transform 1 0 241132 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_2620
timestamp 1676037725
transform 1 0 242144 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2633
timestamp 1676037725
transform 1 0 243340 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2645
timestamp 1676037725
transform 1 0 244444 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2670
timestamp 1676037725
transform 1 0 246744 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2684
timestamp 1676037725
transform 1 0 248032 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2689
timestamp 1676037725
transform 1 0 248492 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2712
timestamp 1676037725
transform 1 0 250608 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2726
timestamp 1676037725
transform 1 0 251896 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2740
timestamp 1676037725
transform 1 0 253184 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2745
timestamp 1676037725
transform 1 0 253644 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_2757
timestamp 1676037725
transform 1 0 254748 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2786
timestamp 1676037725
transform 1 0 257416 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2790
timestamp 1676037725
transform 1 0 257784 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2798
timestamp 1676037725
transform 1 0 258520 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2801
timestamp 1676037725
transform 1 0 258796 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2813
timestamp 1676037725
transform 1 0 259900 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_2817
timestamp 1676037725
transform 1 0 260268 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2824
timestamp 1676037725
transform 1 0 260912 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2833
timestamp 1676037725
transform 1 0 261740 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2842
timestamp 1676037725
transform 1 0 262568 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2851
timestamp 1676037725
transform 1 0 263396 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_2855
timestamp 1676037725
transform 1 0 263764 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2857
timestamp 1676037725
transform 1 0 263948 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2864
timestamp 1676037725
transform 1 0 264592 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2873
timestamp 1676037725
transform 1 0 265420 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2882
timestamp 1676037725
transform 1 0 266248 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2891
timestamp 1676037725
transform 1 0 267076 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2900
timestamp 1676037725
transform 1 0 267904 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_2909
timestamp 1676037725
transform 1 0 268732 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2913
timestamp 1676037725
transform 1 0 269100 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2920
timestamp 1676037725
transform 1 0 269744 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_2928
timestamp 1676037725
transform 1 0 270480 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_3
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_8
timestamp 1676037725
transform 1 0 1840 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_20
timestamp 1676037725
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_47
timestamp 1676037725
transform 1 0 5428 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_59
timestamp 1676037725
transform 1 0 6532 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_71
timestamp 1676037725
transform 1 0 7636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1676037725
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1676037725
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1676037725
transform 1 0 11132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1676037725
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1676037725
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1676037725
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_159
timestamp 1676037725
transform 1 0 15732 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_171
timestamp 1676037725
transform 1 0 16836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_183
timestamp 1676037725
transform 1 0 17940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1676037725
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1676037725
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_221
timestamp 1676037725
transform 1 0 21436 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_229
timestamp 1676037725
transform 1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_238
timestamp 1676037725
transform 1 0 23000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_247
timestamp 1676037725
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1676037725
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_257
timestamp 1676037725
transform 1 0 24748 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_261
timestamp 1676037725
transform 1 0 25116 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_268
timestamp 1676037725
transform 1 0 25760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_282
timestamp 1676037725
transform 1 0 27048 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_290
timestamp 1676037725
transform 1 0 27784 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_302
timestamp 1676037725
transform 1 0 28888 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_315
timestamp 1676037725
transform 1 0 30084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_327
timestamp 1676037725
transform 1 0 31188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_333
timestamp 1676037725
transform 1 0 31740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_339
timestamp 1676037725
transform 1 0 32292 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_347
timestamp 1676037725
transform 1 0 33028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_359
timestamp 1676037725
transform 1 0 34132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1676037725
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1676037725
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_389
timestamp 1676037725
transform 1 0 36892 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_397
timestamp 1676037725
transform 1 0 37628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_418
timestamp 1676037725
transform 1 0 39560 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_441
timestamp 1676037725
transform 1 0 41676 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_463
timestamp 1676037725
transform 1 0 43700 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_475
timestamp 1676037725
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_477
timestamp 1676037725
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_489
timestamp 1676037725
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_501
timestamp 1676037725
transform 1 0 47196 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_513
timestamp 1676037725
transform 1 0 48300 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_525
timestamp 1676037725
transform 1 0 49404 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_531
timestamp 1676037725
transform 1 0 49956 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_533
timestamp 1676037725
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_545
timestamp 1676037725
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_557
timestamp 1676037725
transform 1 0 52348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_569
timestamp 1676037725
transform 1 0 53452 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_573
timestamp 1676037725
transform 1 0 53820 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_580
timestamp 1676037725
transform 1 0 54464 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_589
timestamp 1676037725
transform 1 0 55292 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_595
timestamp 1676037725
transform 1 0 55844 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_607
timestamp 1676037725
transform 1 0 56948 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_615
timestamp 1676037725
transform 1 0 57684 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_620
timestamp 1676037725
transform 1 0 58144 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_636
timestamp 1676037725
transform 1 0 59616 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_645
timestamp 1676037725
transform 1 0 60444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_651
timestamp 1676037725
transform 1 0 60996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_655
timestamp 1676037725
transform 1 0 61364 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_660
timestamp 1676037725
transform 1 0 61824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_668
timestamp 1676037725
transform 1 0 62560 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_676
timestamp 1676037725
transform 1 0 63296 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_688
timestamp 1676037725
transform 1 0 64400 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_701
timestamp 1676037725
transform 1 0 65596 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_707
timestamp 1676037725
transform 1 0 66148 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_721
timestamp 1676037725
transform 1 0 67436 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_733
timestamp 1676037725
transform 1 0 68540 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_745
timestamp 1676037725
transform 1 0 69644 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_753
timestamp 1676037725
transform 1 0 70380 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_757
timestamp 1676037725
transform 1 0 70748 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_769
timestamp 1676037725
transform 1 0 71852 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_781
timestamp 1676037725
transform 1 0 72956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_793
timestamp 1676037725
transform 1 0 74060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_805
timestamp 1676037725
transform 1 0 75164 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_811
timestamp 1676037725
transform 1 0 75716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_813
timestamp 1676037725
transform 1 0 75900 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_829
timestamp 1676037725
transform 1 0 77372 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_841
timestamp 1676037725
transform 1 0 78476 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_853
timestamp 1676037725
transform 1 0 79580 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_865
timestamp 1676037725
transform 1 0 80684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_869
timestamp 1676037725
transform 1 0 81052 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_885
timestamp 1676037725
transform 1 0 82524 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_897
timestamp 1676037725
transform 1 0 83628 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_909
timestamp 1676037725
transform 1 0 84732 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_921
timestamp 1676037725
transform 1 0 85836 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_925
timestamp 1676037725
transform 1 0 86204 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_937
timestamp 1676037725
transform 1 0 87308 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_949
timestamp 1676037725
transform 1 0 88412 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_952
timestamp 1676037725
transform 1 0 88688 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_959
timestamp 1676037725
transform 1 0 89332 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_965
timestamp 1676037725
transform 1 0 89884 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_970
timestamp 1676037725
transform 1 0 90344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_978
timestamp 1676037725
transform 1 0 91080 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_981
timestamp 1676037725
transform 1 0 91356 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_993
timestamp 1676037725
transform 1 0 92460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1001
timestamp 1676037725
transform 1 0 93196 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1009
timestamp 1676037725
transform 1 0 93932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1034
timestamp 1676037725
transform 1 0 96232 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_1037
timestamp 1676037725
transform 1 0 96508 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1043
timestamp 1676037725
transform 1 0 97060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1065
timestamp 1676037725
transform 1 0 99084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1090
timestamp 1676037725
transform 1 0 101384 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_1093
timestamp 1676037725
transform 1 0 101660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_1117
timestamp 1676037725
transform 1 0 103868 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1146
timestamp 1676037725
transform 1 0 106536 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1149
timestamp 1676037725
transform 1 0 106812 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1172
timestamp 1676037725
transform 1 0 108928 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_1197
timestamp 1676037725
transform 1 0 111228 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1203
timestamp 1676037725
transform 1 0 111780 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1205
timestamp 1676037725
transform 1 0 111964 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_1228
timestamp 1676037725
transform 1 0 114080 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_1257
timestamp 1676037725
transform 1 0 116748 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1261
timestamp 1676037725
transform 1 0 117116 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1266
timestamp 1676037725
transform 1 0 117576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1273
timestamp 1676037725
transform 1 0 118220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_1280
timestamp 1676037725
transform 1 0 118864 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1286
timestamp 1676037725
transform 1 0 119416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_1308
timestamp 1676037725
transform 1 0 121440 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1317
timestamp 1676037725
transform 1 0 122268 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1323
timestamp 1676037725
transform 1 0 122820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1335
timestamp 1676037725
transform 1 0 123924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1340
timestamp 1676037725
transform 1 0 124384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_1349
timestamp 1676037725
transform 1 0 125212 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1357
timestamp 1676037725
transform 1 0 125948 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1362
timestamp 1676037725
transform 1 0 126408 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1370
timestamp 1676037725
transform 1 0 127144 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_1373
timestamp 1676037725
transform 1 0 127420 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1381
timestamp 1676037725
transform 1 0 128156 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1386
timestamp 1676037725
transform 1 0 128616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1394
timestamp 1676037725
transform 1 0 129352 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1403
timestamp 1676037725
transform 1 0 130180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_1411
timestamp 1676037725
transform 1 0 130916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_1421
timestamp 1676037725
transform 1 0 131836 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1427
timestamp 1676037725
transform 1 0 132388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1429
timestamp 1676037725
transform 1 0 132572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1433
timestamp 1676037725
transform 1 0 132940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1438
timestamp 1676037725
transform 1 0 133400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1446
timestamp 1676037725
transform 1 0 134136 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1450
timestamp 1676037725
transform 1 0 134504 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1456
timestamp 1676037725
transform 1 0 135056 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1468
timestamp 1676037725
transform 1 0 136160 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1480
timestamp 1676037725
transform 1 0 137264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_1485
timestamp 1676037725
transform 1 0 137724 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1493
timestamp 1676037725
transform 1 0 138460 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1498
timestamp 1676037725
transform 1 0 138920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1523
timestamp 1676037725
transform 1 0 141220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_1534
timestamp 1676037725
transform 1 0 142232 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1541
timestamp 1676037725
transform 1 0 142876 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1564
timestamp 1676037725
transform 1 0 144992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_1589
timestamp 1676037725
transform 1 0 147292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1595
timestamp 1676037725
transform 1 0 147844 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_1597
timestamp 1676037725
transform 1 0 148028 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1624
timestamp 1676037725
transform 1 0 150512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_1649
timestamp 1676037725
transform 1 0 152812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1653
timestamp 1676037725
transform 1 0 153180 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1658
timestamp 1676037725
transform 1 0 153640 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1665
timestamp 1676037725
transform 1 0 154284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_1672
timestamp 1676037725
transform 1 0 154928 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1678
timestamp 1676037725
transform 1 0 155480 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1683
timestamp 1676037725
transform 1 0 155940 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1687
timestamp 1676037725
transform 1 0 156308 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1698
timestamp 1676037725
transform 1 0 157320 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1706
timestamp 1676037725
transform 1 0 158056 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1709
timestamp 1676037725
transform 1 0 158332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1720
timestamp 1676037725
transform 1 0 159344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1724
timestamp 1676037725
transform 1 0 159712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1730
timestamp 1676037725
transform 1 0 160264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1738
timestamp 1676037725
transform 1 0 161000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1742
timestamp 1676037725
transform 1 0 161368 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1747
timestamp 1676037725
transform 1 0 161828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_1755
timestamp 1676037725
transform 1 0 162564 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1763
timestamp 1676037725
transform 1 0 163300 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1765
timestamp 1676037725
transform 1 0 163484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_1771
timestamp 1676037725
transform 1 0 164036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_1779
timestamp 1676037725
transform 1 0 164772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1786
timestamp 1676037725
transform 1 0 165416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1794
timestamp 1676037725
transform 1 0 166152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1798
timestamp 1676037725
transform 1 0 166520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_1803
timestamp 1676037725
transform 1 0 166980 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1811
timestamp 1676037725
transform 1 0 167716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_1817
timestamp 1676037725
transform 1 0 168268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1821
timestamp 1676037725
transform 1 0 168636 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1833
timestamp 1676037725
transform 1 0 169740 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1845
timestamp 1676037725
transform 1 0 170844 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1857
timestamp 1676037725
transform 1 0 171948 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_1869
timestamp 1676037725
transform 1 0 173052 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1875
timestamp 1676037725
transform 1 0 173604 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1877
timestamp 1676037725
transform 1 0 173788 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1889
timestamp 1676037725
transform 1 0 174892 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_1901
timestamp 1676037725
transform 1 0 175996 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1907
timestamp 1676037725
transform 1 0 176548 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1918
timestamp 1676037725
transform 1 0 177560 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1930
timestamp 1676037725
transform 1 0 178664 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_1933
timestamp 1676037725
transform 1 0 178940 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1939
timestamp 1676037725
transform 1 0 179492 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1950
timestamp 1676037725
transform 1 0 180504 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1962
timestamp 1676037725
transform 1 0 181608 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1974
timestamp 1676037725
transform 1 0 182712 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1986
timestamp 1676037725
transform 1 0 183816 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_1989
timestamp 1676037725
transform 1 0 184092 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1995
timestamp 1676037725
transform 1 0 184644 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2006
timestamp 1676037725
transform 1 0 185656 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2018
timestamp 1676037725
transform 1 0 186760 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2030
timestamp 1676037725
transform 1 0 187864 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2042
timestamp 1676037725
transform 1 0 188968 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2045
timestamp 1676037725
transform 1 0 189244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2061
timestamp 1676037725
transform 1 0 190716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2069
timestamp 1676037725
transform 1 0 191452 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2077
timestamp 1676037725
transform 1 0 192188 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_2089
timestamp 1676037725
transform 1 0 193292 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_2097
timestamp 1676037725
transform 1 0 194028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_2101
timestamp 1676037725
transform 1 0 194396 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2108
timestamp 1676037725
transform 1 0 195040 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2124
timestamp 1676037725
transform 1 0 196512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2128
timestamp 1676037725
transform 1 0 196880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2133
timestamp 1676037725
transform 1 0 197340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2137
timestamp 1676037725
transform 1 0 197708 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2142
timestamp 1676037725
transform 1 0 198168 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_2150
timestamp 1676037725
transform 1 0 198904 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_2157
timestamp 1676037725
transform 1 0 199548 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2163
timestamp 1676037725
transform 1 0 200100 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2168
timestamp 1676037725
transform 1 0 200560 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2172
timestamp 1676037725
transform 1 0 200928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2177
timestamp 1676037725
transform 1 0 201388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_2185
timestamp 1676037725
transform 1 0 202124 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2193
timestamp 1676037725
transform 1 0 202860 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2200
timestamp 1676037725
transform 1 0 203504 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2208
timestamp 1676037725
transform 1 0 204240 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2213
timestamp 1676037725
transform 1 0 204700 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2225
timestamp 1676037725
transform 1 0 205804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2237
timestamp 1676037725
transform 1 0 206908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2249
timestamp 1676037725
transform 1 0 208012 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2253
timestamp 1676037725
transform 1 0 208380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2266
timestamp 1676037725
transform 1 0 209576 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2269
timestamp 1676037725
transform 1 0 209852 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2292
timestamp 1676037725
transform 1 0 211968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_2317
timestamp 1676037725
transform 1 0 214268 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2323
timestamp 1676037725
transform 1 0 214820 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2325
timestamp 1676037725
transform 1 0 215004 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2348
timestamp 1676037725
transform 1 0 217120 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_2373
timestamp 1676037725
transform 1 0 219420 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2379
timestamp 1676037725
transform 1 0 219972 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_2381
timestamp 1676037725
transform 1 0 220156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2390
timestamp 1676037725
transform 1 0 220984 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_2415
timestamp 1676037725
transform 1 0 223284 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2427
timestamp 1676037725
transform 1 0 224388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2434
timestamp 1676037725
transform 1 0 225032 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2437
timestamp 1676037725
transform 1 0 225308 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2443
timestamp 1676037725
transform 1 0 225860 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2451
timestamp 1676037725
transform 1 0 226596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_2458
timestamp 1676037725
transform 1 0 227240 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2468
timestamp 1676037725
transform 1 0 228160 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_2480
timestamp 1676037725
transform 1 0 229264 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2490
timestamp 1676037725
transform 1 0 230184 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2493
timestamp 1676037725
transform 1 0 230460 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2499
timestamp 1676037725
transform 1 0 231012 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2507
timestamp 1676037725
transform 1 0 231748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2511
timestamp 1676037725
transform 1 0 232116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2516
timestamp 1676037725
transform 1 0 232576 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2524
timestamp 1676037725
transform 1 0 233312 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_2536
timestamp 1676037725
transform 1 0 234416 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2546
timestamp 1676037725
transform 1 0 235336 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2549
timestamp 1676037725
transform 1 0 235612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2556
timestamp 1676037725
transform 1 0 236256 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2564
timestamp 1676037725
transform 1 0 236992 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2576
timestamp 1676037725
transform 1 0 238096 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2588
timestamp 1676037725
transform 1 0 239200 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2600
timestamp 1676037725
transform 1 0 240304 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2605
timestamp 1676037725
transform 1 0 240764 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2617
timestamp 1676037725
transform 1 0 241868 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2629
timestamp 1676037725
transform 1 0 242972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2633
timestamp 1676037725
transform 1 0 243340 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2644
timestamp 1676037725
transform 1 0 244352 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2658
timestamp 1676037725
transform 1 0 245640 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2661
timestamp 1676037725
transform 1 0 245916 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_2684
timestamp 1676037725
transform 1 0 248032 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_2713
timestamp 1676037725
transform 1 0 250700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2717
timestamp 1676037725
transform 1 0 251068 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2740
timestamp 1676037725
transform 1 0 253184 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2754
timestamp 1676037725
transform 1 0 254472 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2768
timestamp 1676037725
transform 1 0 255760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2773
timestamp 1676037725
transform 1 0 256220 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2796
timestamp 1676037725
transform 1 0 258336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2810
timestamp 1676037725
transform 1 0 259624 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_2820
timestamp 1676037725
transform 1 0 260544 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2829
timestamp 1676037725
transform 1 0 261372 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2836
timestamp 1676037725
transform 1 0 262016 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2844
timestamp 1676037725
transform 1 0 262752 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2852
timestamp 1676037725
transform 1 0 263488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2856
timestamp 1676037725
transform 1 0 263856 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2862
timestamp 1676037725
transform 1 0 264408 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2866
timestamp 1676037725
transform 1 0 264776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_2877
timestamp 1676037725
transform 1 0 265788 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2883
timestamp 1676037725
transform 1 0 266340 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2885
timestamp 1676037725
transform 1 0 266524 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_2891
timestamp 1676037725
transform 1 0 267076 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2900
timestamp 1676037725
transform 1 0 267904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2907
timestamp 1676037725
transform 1 0 268548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2916
timestamp 1676037725
transform 1 0 269376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2925
timestamp 1676037725
transform 1 0 270204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_2933
timestamp 1676037725
transform 1 0 270940 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_233
timestamp 1676037725
transform 1 0 22540 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_239
timestamp 1676037725
transform 1 0 23092 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_249
timestamp 1676037725
transform 1 0 24012 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_258
timestamp 1676037725
transform 1 0 24840 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_270
timestamp 1676037725
transform 1 0 25944 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_278
timestamp 1676037725
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1676037725
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1676037725
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1676037725
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_342
timestamp 1676037725
transform 1 0 32568 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_354
timestamp 1676037725
transform 1 0 33672 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_366
timestamp 1676037725
transform 1 0 34776 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_378
timestamp 1676037725
transform 1 0 35880 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_390
timestamp 1676037725
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_413
timestamp 1676037725
transform 1 0 39100 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_425
timestamp 1676037725
transform 1 0 40204 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_437
timestamp 1676037725
transform 1 0 41308 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_445
timestamp 1676037725
transform 1 0 42044 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_471
timestamp 1676037725
transform 1 0 44436 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_475
timestamp 1676037725
transform 1 0 44804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_487
timestamp 1676037725
transform 1 0 45908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_499
timestamp 1676037725
transform 1 0 47012 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_503
timestamp 1676037725
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_505
timestamp 1676037725
transform 1 0 47564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_525
timestamp 1676037725
transform 1 0 49404 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_529
timestamp 1676037725
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_541
timestamp 1676037725
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_553
timestamp 1676037725
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_559
timestamp 1676037725
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_561
timestamp 1676037725
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_573
timestamp 1676037725
transform 1 0 53820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_577
timestamp 1676037725
transform 1 0 54188 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_582
timestamp 1676037725
transform 1 0 54648 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_594
timestamp 1676037725
transform 1 0 55752 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_606
timestamp 1676037725
transform 1 0 56856 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_614
timestamp 1676037725
transform 1 0 57592 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_617
timestamp 1676037725
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_629
timestamp 1676037725
transform 1 0 58972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_641
timestamp 1676037725
transform 1 0 60076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_653
timestamp 1676037725
transform 1 0 61180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_665
timestamp 1676037725
transform 1 0 62284 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_671
timestamp 1676037725
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_673
timestamp 1676037725
transform 1 0 63020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_685
timestamp 1676037725
transform 1 0 64124 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_697
timestamp 1676037725
transform 1 0 65228 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_712
timestamp 1676037725
transform 1 0 66608 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_724
timestamp 1676037725
transform 1 0 67712 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_729
timestamp 1676037725
transform 1 0 68172 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_741
timestamp 1676037725
transform 1 0 69276 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_753
timestamp 1676037725
transform 1 0 70380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_765
timestamp 1676037725
transform 1 0 71484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_777
timestamp 1676037725
transform 1 0 72588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_783
timestamp 1676037725
transform 1 0 73140 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_785
timestamp 1676037725
transform 1 0 73324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_797
timestamp 1676037725
transform 1 0 74428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_809
timestamp 1676037725
transform 1 0 75532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_821
timestamp 1676037725
transform 1 0 76636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_833
timestamp 1676037725
transform 1 0 77740 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_839
timestamp 1676037725
transform 1 0 78292 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_841
timestamp 1676037725
transform 1 0 78476 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_853
timestamp 1676037725
transform 1 0 79580 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_865
timestamp 1676037725
transform 1 0 80684 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_877
timestamp 1676037725
transform 1 0 81788 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_889
timestamp 1676037725
transform 1 0 82892 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_895
timestamp 1676037725
transform 1 0 83444 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_897
timestamp 1676037725
transform 1 0 83628 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_909
timestamp 1676037725
transform 1 0 84732 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_921
timestamp 1676037725
transform 1 0 85836 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_933
timestamp 1676037725
transform 1 0 86940 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_945
timestamp 1676037725
transform 1 0 88044 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_951
timestamp 1676037725
transform 1 0 88596 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_953
timestamp 1676037725
transform 1 0 88780 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_963
timestamp 1676037725
transform 1 0 89700 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_971
timestamp 1676037725
transform 1 0 90436 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_977
timestamp 1676037725
transform 1 0 90988 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_985
timestamp 1676037725
transform 1 0 91724 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_990
timestamp 1676037725
transform 1 0 92184 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_998
timestamp 1676037725
transform 1 0 92920 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1006
timestamp 1676037725
transform 1 0 93656 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1009
timestamp 1676037725
transform 1 0 93932 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1015
timestamp 1676037725
transform 1 0 94484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_1024
timestamp 1676037725
transform 1 0 95312 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1037
timestamp 1676037725
transform 1 0 96508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1062
timestamp 1676037725
transform 1 0 98808 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1065
timestamp 1676037725
transform 1 0 99084 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_1069
timestamp 1676037725
transform 1 0 99452 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1091
timestamp 1676037725
transform 1 0 101476 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1116
timestamp 1676037725
transform 1 0 103776 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1121
timestamp 1676037725
transform 1 0 104236 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_1144
timestamp 1676037725
transform 1 0 106352 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_1152
timestamp 1676037725
transform 1 0 107088 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1174
timestamp 1676037725
transform 1 0 109112 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1177
timestamp 1676037725
transform 1 0 109388 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1182
timestamp 1676037725
transform 1 0 109848 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_1193
timestamp 1676037725
transform 1 0 110860 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1201
timestamp 1676037725
transform 1 0 111596 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_1224
timestamp 1676037725
transform 1 0 113712 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1233
timestamp 1676037725
transform 1 0 114540 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_1237
timestamp 1676037725
transform 1 0 114908 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_1259
timestamp 1676037725
transform 1 0 116932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1286
timestamp 1676037725
transform 1 0 119416 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1289
timestamp 1676037725
transform 1 0 119692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1295
timestamp 1676037725
transform 1 0 120244 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_1299
timestamp 1676037725
transform 1 0 120612 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1321
timestamp 1676037725
transform 1 0 122636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_1333
timestamp 1676037725
transform 1 0 123740 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_1341
timestamp 1676037725
transform 1 0 124476 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1345
timestamp 1676037725
transform 1 0 124844 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1357
timestamp 1676037725
transform 1 0 125948 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1369
timestamp 1676037725
transform 1 0 127052 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1381
timestamp 1676037725
transform 1 0 128156 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_1393
timestamp 1676037725
transform 1 0 129260 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_1399
timestamp 1676037725
transform 1 0 129812 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1401
timestamp 1676037725
transform 1 0 129996 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1413
timestamp 1676037725
transform 1 0 131100 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1425
timestamp 1676037725
transform 1 0 132204 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1437
timestamp 1676037725
transform 1 0 133308 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_1449
timestamp 1676037725
transform 1 0 134412 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_1455
timestamp 1676037725
transform 1 0 134964 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1457
timestamp 1676037725
transform 1 0 135148 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1462
timestamp 1676037725
transform 1 0 135608 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1474
timestamp 1676037725
transform 1 0 136712 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1486
timestamp 1676037725
transform 1 0 137816 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1493
timestamp 1676037725
transform 1 0 138460 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1500
timestamp 1676037725
transform 1 0 139104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1507
timestamp 1676037725
transform 1 0 139748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_1511
timestamp 1676037725
transform 1 0 140116 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1513
timestamp 1676037725
transform 1 0 140300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1536
timestamp 1676037725
transform 1 0 142416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_1540
timestamp 1676037725
transform 1 0 142784 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_1562
timestamp 1676037725
transform 1 0 144808 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1569
timestamp 1676037725
transform 1 0 145452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1592
timestamp 1676037725
transform 1 0 147568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_1596
timestamp 1676037725
transform 1 0 147936 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1599
timestamp 1676037725
transform 1 0 148212 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1622
timestamp 1676037725
transform 1 0 150328 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1625
timestamp 1676037725
transform 1 0 150604 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1648
timestamp 1676037725
transform 1 0 152720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1655
timestamp 1676037725
transform 1 0 153364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1662
timestamp 1676037725
transform 1 0 154008 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1669
timestamp 1676037725
transform 1 0 154652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1676
timestamp 1676037725
transform 1 0 155296 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1681
timestamp 1676037725
transform 1 0 155756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1706
timestamp 1676037725
transform 1 0 158056 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1714
timestamp 1676037725
transform 1 0 158792 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1722
timestamp 1676037725
transform 1 0 159528 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1734
timestamp 1676037725
transform 1 0 160632 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1737
timestamp 1676037725
transform 1 0 160908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1749
timestamp 1676037725
transform 1 0 162012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1761
timestamp 1676037725
transform 1 0 163116 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1773
timestamp 1676037725
transform 1 0 164220 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_1785
timestamp 1676037725
transform 1 0 165324 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_1791
timestamp 1676037725
transform 1 0 165876 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1793
timestamp 1676037725
transform 1 0 166060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_1805
timestamp 1676037725
transform 1 0 167164 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1816
timestamp 1676037725
transform 1 0 168176 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1828
timestamp 1676037725
transform 1 0 169280 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_1840
timestamp 1676037725
transform 1 0 170384 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1849
timestamp 1676037725
transform 1 0 171212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1861
timestamp 1676037725
transform 1 0 172316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1873
timestamp 1676037725
transform 1 0 173420 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1885
timestamp 1676037725
transform 1 0 174524 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_1897
timestamp 1676037725
transform 1 0 175628 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_1903
timestamp 1676037725
transform 1 0 176180 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1905
timestamp 1676037725
transform 1 0 176364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1917
timestamp 1676037725
transform 1 0 177468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1929
timestamp 1676037725
transform 1 0 178572 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1941
timestamp 1676037725
transform 1 0 179676 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_1953
timestamp 1676037725
transform 1 0 180780 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_1959
timestamp 1676037725
transform 1 0 181332 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1961
timestamp 1676037725
transform 1 0 181516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1973
timestamp 1676037725
transform 1 0 182620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1985
timestamp 1676037725
transform 1 0 183724 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1997
timestamp 1676037725
transform 1 0 184828 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_2009
timestamp 1676037725
transform 1 0 185932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2015
timestamp 1676037725
transform 1 0 186484 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2017
timestamp 1676037725
transform 1 0 186668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2029
timestamp 1676037725
transform 1 0 187772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2041
timestamp 1676037725
transform 1 0 188876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_2053
timestamp 1676037725
transform 1 0 189980 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_2061
timestamp 1676037725
transform 1 0 190716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2067
timestamp 1676037725
transform 1 0 191268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2071
timestamp 1676037725
transform 1 0 191636 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2073
timestamp 1676037725
transform 1 0 191820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2085
timestamp 1676037725
transform 1 0 192924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2097
timestamp 1676037725
transform 1 0 194028 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2109
timestamp 1676037725
transform 1 0 195132 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_2121
timestamp 1676037725
transform 1 0 196236 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2127
timestamp 1676037725
transform 1 0 196788 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2129
timestamp 1676037725
transform 1 0 196972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2141
timestamp 1676037725
transform 1 0 198076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2153
timestamp 1676037725
transform 1 0 199180 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2165
timestamp 1676037725
transform 1 0 200284 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_2177
timestamp 1676037725
transform 1 0 201388 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2183
timestamp 1676037725
transform 1 0 201940 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_2185
timestamp 1676037725
transform 1 0 202124 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_2193
timestamp 1676037725
transform 1 0 202860 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2199
timestamp 1676037725
transform 1 0 203412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2211
timestamp 1676037725
transform 1 0 204516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2223
timestamp 1676037725
transform 1 0 205620 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2235
timestamp 1676037725
transform 1 0 206724 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2239
timestamp 1676037725
transform 1 0 207092 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_2241
timestamp 1676037725
transform 1 0 207276 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_2253
timestamp 1676037725
transform 1 0 208380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_2257
timestamp 1676037725
transform 1 0 208748 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2280
timestamp 1676037725
transform 1 0 210864 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_2293
timestamp 1676037725
transform 1 0 212060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_2297
timestamp 1676037725
transform 1 0 212428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2320
timestamp 1676037725
transform 1 0 214544 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_2345
timestamp 1676037725
transform 1 0 216844 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2351
timestamp 1676037725
transform 1 0 217396 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_2353
timestamp 1676037725
transform 1 0 217580 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2380
timestamp 1676037725
transform 1 0 220064 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2390
timestamp 1676037725
transform 1 0 220984 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2403
timestamp 1676037725
transform 1 0 222180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2407
timestamp 1676037725
transform 1 0 222548 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_2409
timestamp 1676037725
transform 1 0 222732 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2415
timestamp 1676037725
transform 1 0 223284 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2437
timestamp 1676037725
transform 1 0 225308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2444
timestamp 1676037725
transform 1 0 225952 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2451
timestamp 1676037725
transform 1 0 226596 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2463
timestamp 1676037725
transform 1 0 227700 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2465
timestamp 1676037725
transform 1 0 227884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2477
timestamp 1676037725
transform 1 0 228988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2489
timestamp 1676037725
transform 1 0 230092 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2501
timestamp 1676037725
transform 1 0 231196 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_2513
timestamp 1676037725
transform 1 0 232300 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2519
timestamp 1676037725
transform 1 0 232852 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2521
timestamp 1676037725
transform 1 0 233036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2533
timestamp 1676037725
transform 1 0 234140 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2545
timestamp 1676037725
transform 1 0 235244 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2549
timestamp 1676037725
transform 1 0 235612 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2553
timestamp 1676037725
transform 1 0 235980 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_2565
timestamp 1676037725
transform 1 0 237084 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_2573
timestamp 1676037725
transform 1 0 237820 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2577
timestamp 1676037725
transform 1 0 238188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2589
timestamp 1676037725
transform 1 0 239292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2601
timestamp 1676037725
transform 1 0 240396 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2613
timestamp 1676037725
transform 1 0 241500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_2625
timestamp 1676037725
transform 1 0 242604 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2631
timestamp 1676037725
transform 1 0 243156 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_2633
timestamp 1676037725
transform 1 0 243340 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2639
timestamp 1676037725
transform 1 0 243892 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2646
timestamp 1676037725
transform 1 0 244536 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2671
timestamp 1676037725
transform 1 0 246836 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_2685
timestamp 1676037725
transform 1 0 248124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_2689
timestamp 1676037725
transform 1 0 248492 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2712
timestamp 1676037725
transform 1 0 250608 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_2737
timestamp 1676037725
transform 1 0 252908 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2743
timestamp 1676037725
transform 1 0 253460 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_2745
timestamp 1676037725
transform 1 0 253644 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2757
timestamp 1676037725
transform 1 0 254748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2782
timestamp 1676037725
transform 1 0 257048 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2796
timestamp 1676037725
transform 1 0 258336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_2801
timestamp 1676037725
transform 1 0 258796 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_2809
timestamp 1676037725
transform 1 0 259532 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2813
timestamp 1676037725
transform 1 0 259900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2822
timestamp 1676037725
transform 1 0 260728 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2830
timestamp 1676037725
transform 1 0 261464 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2838
timestamp 1676037725
transform 1 0 262200 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_2850
timestamp 1676037725
transform 1 0 263304 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2857
timestamp 1676037725
transform 1 0 263948 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_2869
timestamp 1676037725
transform 1 0 265052 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_2877
timestamp 1676037725
transform 1 0 265788 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2882
timestamp 1676037725
transform 1 0 266248 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2889
timestamp 1676037725
transform 1 0 266892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2896
timestamp 1676037725
transform 1 0 267536 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2903
timestamp 1676037725
transform 1 0 268180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_2910
timestamp 1676037725
transform 1 0 268824 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_2913
timestamp 1676037725
transform 1 0 269100 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_2925
timestamp 1676037725
transform 1 0 270204 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_2934
timestamp 1676037725
transform 1 0 271032 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_233
timestamp 1676037725
transform 1 0 22540 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_241
timestamp 1676037725
transform 1 0 23276 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_246
timestamp 1676037725
transform 1 0 23736 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1676037725
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1676037725
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1676037725
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1676037725
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1676037725
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1676037725
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1676037725
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1676037725
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_377
timestamp 1676037725
transform 1 0 35788 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_399
timestamp 1676037725
transform 1 0 37812 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_411
timestamp 1676037725
transform 1 0 38916 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1676037725
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_427
timestamp 1676037725
transform 1 0 40388 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_447
timestamp 1676037725
transform 1 0 42228 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_455
timestamp 1676037725
transform 1 0 42964 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_474
timestamp 1676037725
transform 1 0 44712 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_477
timestamp 1676037725
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_489
timestamp 1676037725
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_501
timestamp 1676037725
transform 1 0 47196 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_509
timestamp 1676037725
transform 1 0 47932 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_528
timestamp 1676037725
transform 1 0 49680 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_533
timestamp 1676037725
transform 1 0 50140 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_553
timestamp 1676037725
transform 1 0 51980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_565
timestamp 1676037725
transform 1 0 53084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_577
timestamp 1676037725
transform 1 0 54188 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_585
timestamp 1676037725
transform 1 0 54924 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_589
timestamp 1676037725
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_601
timestamp 1676037725
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_613
timestamp 1676037725
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_625
timestamp 1676037725
transform 1 0 58604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_637
timestamp 1676037725
transform 1 0 59708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_643
timestamp 1676037725
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_645
timestamp 1676037725
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_657
timestamp 1676037725
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_669
timestamp 1676037725
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_681
timestamp 1676037725
transform 1 0 63756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_693
timestamp 1676037725
transform 1 0 64860 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_699
timestamp 1676037725
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_701
timestamp 1676037725
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_713
timestamp 1676037725
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_725
timestamp 1676037725
transform 1 0 67804 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_733
timestamp 1676037725
transform 1 0 68540 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_738
timestamp 1676037725
transform 1 0 69000 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_750
timestamp 1676037725
transform 1 0 70104 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_757
timestamp 1676037725
transform 1 0 70748 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_769
timestamp 1676037725
transform 1 0 71852 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_781
timestamp 1676037725
transform 1 0 72956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_793
timestamp 1676037725
transform 1 0 74060 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_805
timestamp 1676037725
transform 1 0 75164 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_811
timestamp 1676037725
transform 1 0 75716 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_813
timestamp 1676037725
transform 1 0 75900 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_825
timestamp 1676037725
transform 1 0 77004 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_837
timestamp 1676037725
transform 1 0 78108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_849
timestamp 1676037725
transform 1 0 79212 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_861
timestamp 1676037725
transform 1 0 80316 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_867
timestamp 1676037725
transform 1 0 80868 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_869
timestamp 1676037725
transform 1 0 81052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_881
timestamp 1676037725
transform 1 0 82156 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_893
timestamp 1676037725
transform 1 0 83260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_905
timestamp 1676037725
transform 1 0 84364 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_917
timestamp 1676037725
transform 1 0 85468 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_923
timestamp 1676037725
transform 1 0 86020 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_925
timestamp 1676037725
transform 1 0 86204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_937
timestamp 1676037725
transform 1 0 87308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_949
timestamp 1676037725
transform 1 0 88412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_961
timestamp 1676037725
transform 1 0 89516 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_973
timestamp 1676037725
transform 1 0 90620 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_979
timestamp 1676037725
transform 1 0 91172 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_981
timestamp 1676037725
transform 1 0 91356 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_990
timestamp 1676037725
transform 1 0 92184 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_997
timestamp 1676037725
transform 1 0 92828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_1005
timestamp 1676037725
transform 1 0 93564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_1030
timestamp 1676037725
transform 1 0 95864 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_1037
timestamp 1676037725
transform 1 0 96508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1041
timestamp 1676037725
transform 1 0 96876 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_1047
timestamp 1676037725
transform 1 0 97428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_1061
timestamp 1676037725
transform 1 0 98716 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_1086
timestamp 1676037725
transform 1 0 101016 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1093
timestamp 1676037725
transform 1 0 101660 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_1100
timestamp 1676037725
transform 1 0 102304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1107
timestamp 1676037725
transform 1 0 102948 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1111
timestamp 1676037725
transform 1 0 103316 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_1134
timestamp 1676037725
transform 1 0 105432 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1138
timestamp 1676037725
transform 1 0 105800 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1146
timestamp 1676037725
transform 1 0 106536 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1149
timestamp 1676037725
transform 1 0 106812 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_1172
timestamp 1676037725
transform 1 0 108928 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1180
timestamp 1676037725
transform 1 0 109664 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1202
timestamp 1676037725
transform 1 0 111688 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1205
timestamp 1676037725
transform 1 0 111964 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_1228
timestamp 1676037725
transform 1 0 114080 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1236
timestamp 1676037725
transform 1 0 114816 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1258
timestamp 1676037725
transform 1 0 116840 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_1261
timestamp 1676037725
transform 1 0 117116 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1267
timestamp 1676037725
transform 1 0 117668 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_1289
timestamp 1676037725
transform 1 0 119692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1314
timestamp 1676037725
transform 1 0 121992 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1317
timestamp 1676037725
transform 1 0 122268 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1322
timestamp 1676037725
transform 1 0 122728 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1334
timestamp 1676037725
transform 1 0 123832 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1346
timestamp 1676037725
transform 1 0 124936 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1358
timestamp 1676037725
transform 1 0 126040 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1370
timestamp 1676037725
transform 1 0 127144 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1373
timestamp 1676037725
transform 1 0 127420 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1385
timestamp 1676037725
transform 1 0 128524 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1397
timestamp 1676037725
transform 1 0 129628 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1409
timestamp 1676037725
transform 1 0 130732 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_1421
timestamp 1676037725
transform 1 0 131836 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1427
timestamp 1676037725
transform 1 0 132388 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1429
timestamp 1676037725
transform 1 0 132572 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1441
timestamp 1676037725
transform 1 0 133676 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1453
timestamp 1676037725
transform 1 0 134780 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1465
timestamp 1676037725
transform 1 0 135884 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_1477
timestamp 1676037725
transform 1 0 136988 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1483
timestamp 1676037725
transform 1 0 137540 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_1485
timestamp 1676037725
transform 1 0 137724 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_1494
timestamp 1676037725
transform 1 0 138552 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_1501
timestamp 1676037725
transform 1 0 139196 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_1526
timestamp 1676037725
transform 1 0 141496 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_1537
timestamp 1676037725
transform 1 0 142508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1541
timestamp 1676037725
transform 1 0 142876 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_1564
timestamp 1676037725
transform 1 0 144992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_1589
timestamp 1676037725
transform 1 0 147292 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1595
timestamp 1676037725
transform 1 0 147844 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1597
timestamp 1676037725
transform 1 0 148028 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_1602
timestamp 1676037725
transform 1 0 148488 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1608
timestamp 1676037725
transform 1 0 149040 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_1616
timestamp 1676037725
transform 1 0 149776 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1620
timestamp 1676037725
transform 1 0 150144 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_1642
timestamp 1676037725
transform 1 0 152168 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_1649
timestamp 1676037725
transform 1 0 152812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1653
timestamp 1676037725
transform 1 0 153180 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_1676
timestamp 1676037725
transform 1 0 155296 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_1701
timestamp 1676037725
transform 1 0 157596 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1707
timestamp 1676037725
transform 1 0 158148 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1709
timestamp 1676037725
transform 1 0 158332 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_1714
timestamp 1676037725
transform 1 0 158792 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1721
timestamp 1676037725
transform 1 0 159436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1733
timestamp 1676037725
transform 1 0 160540 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1745
timestamp 1676037725
transform 1 0 161644 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_1757
timestamp 1676037725
transform 1 0 162748 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1763
timestamp 1676037725
transform 1 0 163300 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1765
timestamp 1676037725
transform 1 0 163484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1777
timestamp 1676037725
transform 1 0 164588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1789
timestamp 1676037725
transform 1 0 165692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_1801
timestamp 1676037725
transform 1 0 166796 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1809
timestamp 1676037725
transform 1 0 167532 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_1813
timestamp 1676037725
transform 1 0 167900 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1819
timestamp 1676037725
transform 1 0 168452 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1821
timestamp 1676037725
transform 1 0 168636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1833
timestamp 1676037725
transform 1 0 169740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1845
timestamp 1676037725
transform 1 0 170844 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1857
timestamp 1676037725
transform 1 0 171948 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_1869
timestamp 1676037725
transform 1 0 173052 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1875
timestamp 1676037725
transform 1 0 173604 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1877
timestamp 1676037725
transform 1 0 173788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1889
timestamp 1676037725
transform 1 0 174892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1901
timestamp 1676037725
transform 1 0 175996 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1913
timestamp 1676037725
transform 1 0 177100 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_1925
timestamp 1676037725
transform 1 0 178204 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1931
timestamp 1676037725
transform 1 0 178756 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1933
timestamp 1676037725
transform 1 0 178940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1945
timestamp 1676037725
transform 1 0 180044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1957
timestamp 1676037725
transform 1 0 181148 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1969
timestamp 1676037725
transform 1 0 182252 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_1981
timestamp 1676037725
transform 1 0 183356 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1987
timestamp 1676037725
transform 1 0 183908 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1989
timestamp 1676037725
transform 1 0 184092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2001
timestamp 1676037725
transform 1 0 185196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2013
timestamp 1676037725
transform 1 0 186300 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2025
timestamp 1676037725
transform 1 0 187404 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_2037
timestamp 1676037725
transform 1 0 188508 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_2043
timestamp 1676037725
transform 1 0 189060 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2045
timestamp 1676037725
transform 1 0 189244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2057
timestamp 1676037725
transform 1 0 190348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2069
timestamp 1676037725
transform 1 0 191452 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2081
timestamp 1676037725
transform 1 0 192556 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_2093
timestamp 1676037725
transform 1 0 193660 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_2099
timestamp 1676037725
transform 1 0 194212 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2101
timestamp 1676037725
transform 1 0 194396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2113
timestamp 1676037725
transform 1 0 195500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2125
timestamp 1676037725
transform 1 0 196604 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2137
timestamp 1676037725
transform 1 0 197708 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_2149
timestamp 1676037725
transform 1 0 198812 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_2155
timestamp 1676037725
transform 1 0 199364 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2157
timestamp 1676037725
transform 1 0 199548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2169
timestamp 1676037725
transform 1 0 200652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2181
timestamp 1676037725
transform 1 0 201756 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2193
timestamp 1676037725
transform 1 0 202860 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_2205
timestamp 1676037725
transform 1 0 203964 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_2211
timestamp 1676037725
transform 1 0 204516 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2213
timestamp 1676037725
transform 1 0 204700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2225
timestamp 1676037725
transform 1 0 205804 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_2237
timestamp 1676037725
transform 1 0 206908 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_2259
timestamp 1676037725
transform 1 0 208932 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_2267
timestamp 1676037725
transform 1 0 209668 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_2269
timestamp 1676037725
transform 1 0 209852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2281
timestamp 1676037725
transform 1 0 210956 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2294
timestamp 1676037725
transform 1 0 212152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2307
timestamp 1676037725
transform 1 0 213348 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2314
timestamp 1676037725
transform 1 0 213992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_2321
timestamp 1676037725
transform 1 0 214636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2325
timestamp 1676037725
transform 1 0 215004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_2329
timestamp 1676037725
transform 1 0 215372 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_2334
timestamp 1676037725
transform 1 0 215832 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2346
timestamp 1676037725
transform 1 0 216936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_2350
timestamp 1676037725
transform 1 0 217304 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_2372
timestamp 1676037725
transform 1 0 219328 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2381
timestamp 1676037725
transform 1 0 220156 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2386
timestamp 1676037725
transform 1 0 220616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_2390
timestamp 1676037725
transform 1 0 220984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2412
timestamp 1676037725
transform 1 0 223008 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2425
timestamp 1676037725
transform 1 0 224204 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2432
timestamp 1676037725
transform 1 0 224848 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2437
timestamp 1676037725
transform 1 0 225308 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2460
timestamp 1676037725
transform 1 0 227424 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2464
timestamp 1676037725
transform 1 0 227792 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2476
timestamp 1676037725
transform 1 0 228896 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2488
timestamp 1676037725
transform 1 0 230000 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2493
timestamp 1676037725
transform 1 0 230460 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2505
timestamp 1676037725
transform 1 0 231564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2517
timestamp 1676037725
transform 1 0 232668 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2529
timestamp 1676037725
transform 1 0 233772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_2541
timestamp 1676037725
transform 1 0 234876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_2547
timestamp 1676037725
transform 1 0 235428 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2549
timestamp 1676037725
transform 1 0 235612 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2561
timestamp 1676037725
transform 1 0 236716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2573
timestamp 1676037725
transform 1 0 237820 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2585
timestamp 1676037725
transform 1 0 238924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_2597
timestamp 1676037725
transform 1 0 240028 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_2603
timestamp 1676037725
transform 1 0 240580 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2605
timestamp 1676037725
transform 1 0 240764 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2617
timestamp 1676037725
transform 1 0 241868 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2629
timestamp 1676037725
transform 1 0 242972 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_2641
timestamp 1676037725
transform 1 0 244076 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2648
timestamp 1676037725
transform 1 0 244720 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2658
timestamp 1676037725
transform 1 0 245640 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_2661
timestamp 1676037725
transform 1 0 245916 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_2670
timestamp 1676037725
transform 1 0 246744 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2683
timestamp 1676037725
transform 1 0 247940 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2687
timestamp 1676037725
transform 1 0 248308 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_2710
timestamp 1676037725
transform 1 0 250424 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2717
timestamp 1676037725
transform 1 0 251068 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2729
timestamp 1676037725
transform 1 0 252172 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_2739
timestamp 1676037725
transform 1 0 253092 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2747
timestamp 1676037725
transform 1 0 253828 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2770
timestamp 1676037725
transform 1 0 255944 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2773
timestamp 1676037725
transform 1 0 256220 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2796
timestamp 1676037725
transform 1 0 258336 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2806
timestamp 1676037725
transform 1 0 259256 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2814
timestamp 1676037725
transform 1 0 259992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_2822
timestamp 1676037725
transform 1 0 260728 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2829
timestamp 1676037725
transform 1 0 261372 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2841
timestamp 1676037725
transform 1 0 262476 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2853
timestamp 1676037725
transform 1 0 263580 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2865
timestamp 1676037725
transform 1 0 264684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2877
timestamp 1676037725
transform 1 0 265788 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2882
timestamp 1676037725
transform 1 0 266248 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_2885
timestamp 1676037725
transform 1 0 266524 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2896
timestamp 1676037725
transform 1 0 267536 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2903
timestamp 1676037725
transform 1 0 268180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2910
timestamp 1676037725
transform 1 0 268824 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2917
timestamp 1676037725
transform 1 0 269468 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_2925
timestamp 1676037725
transform 1 0 270204 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2934
timestamp 1676037725
transform 1 0 271032 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1676037725
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1676037725
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1676037725
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1676037725
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1676037725
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1676037725
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1676037725
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_385
timestamp 1676037725
transform 1 0 36524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_390
timestamp 1676037725
transform 1 0 36984 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_413
timestamp 1676037725
transform 1 0 39100 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_417
timestamp 1676037725
transform 1 0 39468 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_421
timestamp 1676037725
transform 1 0 39836 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_433
timestamp 1676037725
transform 1 0 40940 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_439
timestamp 1676037725
transform 1 0 41492 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_446
timestamp 1676037725
transform 1 0 42136 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_457
timestamp 1676037725
transform 1 0 43148 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_487
timestamp 1676037725
transform 1 0 45908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_499
timestamp 1676037725
transform 1 0 47012 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_503
timestamp 1676037725
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_505
timestamp 1676037725
transform 1 0 47564 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_511
timestamp 1676037725
transform 1 0 48116 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_531
timestamp 1676037725
transform 1 0 49956 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_553
timestamp 1676037725
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_559
timestamp 1676037725
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_561
timestamp 1676037725
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_573
timestamp 1676037725
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_585
timestamp 1676037725
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_597
timestamp 1676037725
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_609
timestamp 1676037725
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_615
timestamp 1676037725
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_617
timestamp 1676037725
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_629
timestamp 1676037725
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_641
timestamp 1676037725
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_653
timestamp 1676037725
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_665
timestamp 1676037725
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_671
timestamp 1676037725
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_673
timestamp 1676037725
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_685
timestamp 1676037725
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_697
timestamp 1676037725
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_711
timestamp 1676037725
transform 1 0 66516 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_716
timestamp 1676037725
transform 1 0 66976 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_729
timestamp 1676037725
transform 1 0 68172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_741
timestamp 1676037725
transform 1 0 69276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_753
timestamp 1676037725
transform 1 0 70380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_765
timestamp 1676037725
transform 1 0 71484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_777
timestamp 1676037725
transform 1 0 72588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_783
timestamp 1676037725
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_785
timestamp 1676037725
transform 1 0 73324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_797
timestamp 1676037725
transform 1 0 74428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_809
timestamp 1676037725
transform 1 0 75532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_821
timestamp 1676037725
transform 1 0 76636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_833
timestamp 1676037725
transform 1 0 77740 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_839
timestamp 1676037725
transform 1 0 78292 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_841
timestamp 1676037725
transform 1 0 78476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_853
timestamp 1676037725
transform 1 0 79580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_865
timestamp 1676037725
transform 1 0 80684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_877
timestamp 1676037725
transform 1 0 81788 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_889
timestamp 1676037725
transform 1 0 82892 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_895
timestamp 1676037725
transform 1 0 83444 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_897
timestamp 1676037725
transform 1 0 83628 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_909
timestamp 1676037725
transform 1 0 84732 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_921
timestamp 1676037725
transform 1 0 85836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_933
timestamp 1676037725
transform 1 0 86940 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_945
timestamp 1676037725
transform 1 0 88044 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_951
timestamp 1676037725
transform 1 0 88596 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_953
timestamp 1676037725
transform 1 0 88780 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_965
timestamp 1676037725
transform 1 0 89884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_977
timestamp 1676037725
transform 1 0 90988 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_989
timestamp 1676037725
transform 1 0 92092 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_995
timestamp 1676037725
transform 1 0 92644 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_999
timestamp 1676037725
transform 1 0 93012 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1006
timestamp 1676037725
transform 1 0 93656 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_1009
timestamp 1676037725
transform 1 0 93932 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1015
timestamp 1676037725
transform 1 0 94484 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_1037
timestamp 1676037725
transform 1 0 96508 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1062
timestamp 1676037725
transform 1 0 98808 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1065
timestamp 1676037725
transform 1 0 99084 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_1088
timestamp 1676037725
transform 1 0 101200 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1096
timestamp 1676037725
transform 1 0 101936 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1118
timestamp 1676037725
transform 1 0 103960 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_1121
timestamp 1676037725
transform 1 0 104236 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1125
timestamp 1676037725
transform 1 0 104604 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_1133
timestamp 1676037725
transform 1 0 105340 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_1158
timestamp 1676037725
transform 1 0 107640 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1166
timestamp 1676037725
transform 1 0 108376 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1174
timestamp 1676037725
transform 1 0 109112 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1177
timestamp 1676037725
transform 1 0 109388 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_1182
timestamp 1676037725
transform 1 0 109848 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_1193
timestamp 1676037725
transform 1 0 110860 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_1222
timestamp 1676037725
transform 1 0 113528 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1226
timestamp 1676037725
transform 1 0 113896 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1230
timestamp 1676037725
transform 1 0 114264 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1233
timestamp 1676037725
transform 1 0 114540 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_1256
timestamp 1676037725
transform 1 0 116656 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_1281
timestamp 1676037725
transform 1 0 118956 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1287
timestamp 1676037725
transform 1 0 119508 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_1289
timestamp 1676037725
transform 1 0 119692 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_1304
timestamp 1676037725
transform 1 0 121072 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1329
timestamp 1676037725
transform 1 0 123372 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_1341
timestamp 1676037725
transform 1 0 124476 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1345
timestamp 1676037725
transform 1 0 124844 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1357
timestamp 1676037725
transform 1 0 125948 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1369
timestamp 1676037725
transform 1 0 127052 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1381
timestamp 1676037725
transform 1 0 128156 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_1393
timestamp 1676037725
transform 1 0 129260 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1399
timestamp 1676037725
transform 1 0 129812 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1401
timestamp 1676037725
transform 1 0 129996 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1413
timestamp 1676037725
transform 1 0 131100 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1425
timestamp 1676037725
transform 1 0 132204 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1437
timestamp 1676037725
transform 1 0 133308 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_1449
timestamp 1676037725
transform 1 0 134412 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1455
timestamp 1676037725
transform 1 0 134964 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1457
timestamp 1676037725
transform 1 0 135148 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1469
timestamp 1676037725
transform 1 0 136252 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_1481
timestamp 1676037725
transform 1 0 137356 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_1489
timestamp 1676037725
transform 1 0 138092 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_1499
timestamp 1676037725
transform 1 0 139012 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1510
timestamp 1676037725
transform 1 0 140024 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1513
timestamp 1676037725
transform 1 0 140300 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_1536
timestamp 1676037725
transform 1 0 142416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_1547
timestamp 1676037725
transform 1 0 143428 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_1558
timestamp 1676037725
transform 1 0 144440 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_1565
timestamp 1676037725
transform 1 0 145084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1569
timestamp 1676037725
transform 1 0 145452 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_1592
timestamp 1676037725
transform 1 0 147568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_1603
timestamp 1676037725
transform 1 0 148580 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_1614
timestamp 1676037725
transform 1 0 149592 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1618
timestamp 1676037725
transform 1 0 149960 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1622
timestamp 1676037725
transform 1 0 150328 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1625
timestamp 1676037725
transform 1 0 150604 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_1648
timestamp 1676037725
transform 1 0 152720 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1652
timestamp 1676037725
transform 1 0 153088 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_1674
timestamp 1676037725
transform 1 0 155112 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1681
timestamp 1676037725
transform 1 0 155756 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_1704
timestamp 1676037725
transform 1 0 157872 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_1729
timestamp 1676037725
transform 1 0 160172 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1735
timestamp 1676037725
transform 1 0 160724 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1737
timestamp 1676037725
transform 1 0 160908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1749
timestamp 1676037725
transform 1 0 162012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1761
timestamp 1676037725
transform 1 0 163116 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1773
timestamp 1676037725
transform 1 0 164220 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_1785
timestamp 1676037725
transform 1 0 165324 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1791
timestamp 1676037725
transform 1 0 165876 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1793
timestamp 1676037725
transform 1 0 166060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_1805
timestamp 1676037725
transform 1 0 167164 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1809
timestamp 1676037725
transform 1 0 167532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1818
timestamp 1676037725
transform 1 0 168360 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1830
timestamp 1676037725
transform 1 0 169464 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_1842
timestamp 1676037725
transform 1 0 170568 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1849
timestamp 1676037725
transform 1 0 171212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1861
timestamp 1676037725
transform 1 0 172316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1873
timestamp 1676037725
transform 1 0 173420 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1885
timestamp 1676037725
transform 1 0 174524 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_1897
timestamp 1676037725
transform 1 0 175628 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1903
timestamp 1676037725
transform 1 0 176180 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1905
timestamp 1676037725
transform 1 0 176364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1917
timestamp 1676037725
transform 1 0 177468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1929
timestamp 1676037725
transform 1 0 178572 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1941
timestamp 1676037725
transform 1 0 179676 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_1953
timestamp 1676037725
transform 1 0 180780 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1959
timestamp 1676037725
transform 1 0 181332 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1961
timestamp 1676037725
transform 1 0 181516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1973
timestamp 1676037725
transform 1 0 182620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1985
timestamp 1676037725
transform 1 0 183724 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1997
timestamp 1676037725
transform 1 0 184828 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_2009
timestamp 1676037725
transform 1 0 185932 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_2015
timestamp 1676037725
transform 1 0 186484 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2017
timestamp 1676037725
transform 1 0 186668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2029
timestamp 1676037725
transform 1 0 187772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2041
timestamp 1676037725
transform 1 0 188876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_2053
timestamp 1676037725
transform 1 0 189980 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2059
timestamp 1676037725
transform 1 0 190532 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_2071
timestamp 1676037725
transform 1 0 191636 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2073
timestamp 1676037725
transform 1 0 191820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2085
timestamp 1676037725
transform 1 0 192924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2097
timestamp 1676037725
transform 1 0 194028 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2109
timestamp 1676037725
transform 1 0 195132 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_2121
timestamp 1676037725
transform 1 0 196236 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_2127
timestamp 1676037725
transform 1 0 196788 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2129
timestamp 1676037725
transform 1 0 196972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2141
timestamp 1676037725
transform 1 0 198076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2153
timestamp 1676037725
transform 1 0 199180 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2165
timestamp 1676037725
transform 1 0 200284 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_2177
timestamp 1676037725
transform 1 0 201388 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_2183
timestamp 1676037725
transform 1 0 201940 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2185
timestamp 1676037725
transform 1 0 202124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2197
timestamp 1676037725
transform 1 0 203228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2209
timestamp 1676037725
transform 1 0 204332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_2221
timestamp 1676037725
transform 1 0 205436 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2228
timestamp 1676037725
transform 1 0 206080 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2238
timestamp 1676037725
transform 1 0 207000 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2241
timestamp 1676037725
transform 1 0 207276 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2264
timestamp 1676037725
transform 1 0 209392 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_2289
timestamp 1676037725
transform 1 0 211692 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_2295
timestamp 1676037725
transform 1 0 212244 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_2297
timestamp 1676037725
transform 1 0 212428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_2326
timestamp 1676037725
transform 1 0 215096 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2338
timestamp 1676037725
transform 1 0 216200 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2348
timestamp 1676037725
transform 1 0 217120 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2353
timestamp 1676037725
transform 1 0 217580 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2376
timestamp 1676037725
transform 1 0 219696 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_2401
timestamp 1676037725
transform 1 0 221996 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_2407
timestamp 1676037725
transform 1 0 222548 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2409
timestamp 1676037725
transform 1 0 222732 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2432
timestamp 1676037725
transform 1 0 224848 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_2457
timestamp 1676037725
transform 1 0 227148 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_2463
timestamp 1676037725
transform 1 0 227700 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2465
timestamp 1676037725
transform 1 0 227884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2477
timestamp 1676037725
transform 1 0 228988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2489
timestamp 1676037725
transform 1 0 230092 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2501
timestamp 1676037725
transform 1 0 231196 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_2513
timestamp 1676037725
transform 1 0 232300 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_2519
timestamp 1676037725
transform 1 0 232852 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2521
timestamp 1676037725
transform 1 0 233036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2533
timestamp 1676037725
transform 1 0 234140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2545
timestamp 1676037725
transform 1 0 235244 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2557
timestamp 1676037725
transform 1 0 236348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_2569
timestamp 1676037725
transform 1 0 237452 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_2575
timestamp 1676037725
transform 1 0 238004 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2577
timestamp 1676037725
transform 1 0 238188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2589
timestamp 1676037725
transform 1 0 239292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2601
timestamp 1676037725
transform 1 0 240396 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2613
timestamp 1676037725
transform 1 0 241500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_2625
timestamp 1676037725
transform 1 0 242604 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_2631
timestamp 1676037725
transform 1 0 243156 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_2633
timestamp 1676037725
transform 1 0 243340 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_2641
timestamp 1676037725
transform 1 0 244076 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2647
timestamp 1676037725
transform 1 0 244628 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2672
timestamp 1676037725
transform 1 0 246928 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2686
timestamp 1676037725
transform 1 0 248216 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2689
timestamp 1676037725
transform 1 0 248492 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2712
timestamp 1676037725
transform 1 0 250608 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_2726
timestamp 1676037725
transform 1 0 251896 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2734
timestamp 1676037725
transform 1 0 252632 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2742
timestamp 1676037725
transform 1 0 253368 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2745
timestamp 1676037725
transform 1 0 253644 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_2749
timestamp 1676037725
transform 1 0 254012 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2756
timestamp 1676037725
transform 1 0 254656 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2781
timestamp 1676037725
transform 1 0 256956 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2791
timestamp 1676037725
transform 1 0 257876 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2798
timestamp 1676037725
transform 1 0 258520 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2804
timestamp 1676037725
transform 1 0 259072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2808
timestamp 1676037725
transform 1 0 259440 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2831
timestamp 1676037725
transform 1 0 261556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2843
timestamp 1676037725
transform 1 0 262660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_2855
timestamp 1676037725
transform 1 0 263764 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_2857
timestamp 1676037725
transform 1 0 263948 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_2865
timestamp 1676037725
transform 1 0 264684 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2871
timestamp 1676037725
transform 1 0 265236 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2878
timestamp 1676037725
transform 1 0 265880 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2885
timestamp 1676037725
transform 1 0 266524 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2894
timestamp 1676037725
transform 1 0 267352 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2903
timestamp 1676037725
transform 1 0 268180 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2910
timestamp 1676037725
transform 1 0 268824 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2913
timestamp 1676037725
transform 1 0 269100 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2919
timestamp 1676037725
transform 1 0 269652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2927
timestamp 1676037725
transform 1 0 270388 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2934
timestamp 1676037725
transform 1 0 271032 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1676037725
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1676037725
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1676037725
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1676037725
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1676037725
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_369
timestamp 1676037725
transform 1 0 35052 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_372
timestamp 1676037725
transform 1 0 35328 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_392
timestamp 1676037725
transform 1 0 37168 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_404
timestamp 1676037725
transform 1 0 38272 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_416
timestamp 1676037725
transform 1 0 39376 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_435
timestamp 1676037725
transform 1 0 41124 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_455
timestamp 1676037725
transform 1 0 42964 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_467
timestamp 1676037725
transform 1 0 44068 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_475
timestamp 1676037725
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_477
timestamp 1676037725
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_489
timestamp 1676037725
transform 1 0 46092 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_493
timestamp 1676037725
transform 1 0 46460 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_512
timestamp 1676037725
transform 1 0 48208 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_524
timestamp 1676037725
transform 1 0 49312 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_533
timestamp 1676037725
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_545
timestamp 1676037725
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_557
timestamp 1676037725
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_569
timestamp 1676037725
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_581
timestamp 1676037725
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_587
timestamp 1676037725
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_589
timestamp 1676037725
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_601
timestamp 1676037725
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_613
timestamp 1676037725
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_625
timestamp 1676037725
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_637
timestamp 1676037725
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_643
timestamp 1676037725
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_645
timestamp 1676037725
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_657
timestamp 1676037725
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_669
timestamp 1676037725
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_681
timestamp 1676037725
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_693
timestamp 1676037725
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_699
timestamp 1676037725
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_701
timestamp 1676037725
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_713
timestamp 1676037725
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_725
timestamp 1676037725
transform 1 0 67804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_737
timestamp 1676037725
transform 1 0 68908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_749
timestamp 1676037725
transform 1 0 70012 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_755
timestamp 1676037725
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_757
timestamp 1676037725
transform 1 0 70748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_769
timestamp 1676037725
transform 1 0 71852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_781
timestamp 1676037725
transform 1 0 72956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_793
timestamp 1676037725
transform 1 0 74060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_805
timestamp 1676037725
transform 1 0 75164 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_811
timestamp 1676037725
transform 1 0 75716 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_813
timestamp 1676037725
transform 1 0 75900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_825
timestamp 1676037725
transform 1 0 77004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_837
timestamp 1676037725
transform 1 0 78108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_849
timestamp 1676037725
transform 1 0 79212 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_861
timestamp 1676037725
transform 1 0 80316 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_867
timestamp 1676037725
transform 1 0 80868 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_869
timestamp 1676037725
transform 1 0 81052 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_881
timestamp 1676037725
transform 1 0 82156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_893
timestamp 1676037725
transform 1 0 83260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_905
timestamp 1676037725
transform 1 0 84364 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_917
timestamp 1676037725
transform 1 0 85468 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_923
timestamp 1676037725
transform 1 0 86020 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_925
timestamp 1676037725
transform 1 0 86204 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_937
timestamp 1676037725
transform 1 0 87308 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_949
timestamp 1676037725
transform 1 0 88412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_961
timestamp 1676037725
transform 1 0 89516 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_973
timestamp 1676037725
transform 1 0 90620 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_979
timestamp 1676037725
transform 1 0 91172 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_981
timestamp 1676037725
transform 1 0 91356 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_1004
timestamp 1676037725
transform 1 0 93472 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1012
timestamp 1676037725
transform 1 0 94208 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1034
timestamp 1676037725
transform 1 0 96232 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1037
timestamp 1676037725
transform 1 0 96508 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1043
timestamp 1676037725
transform 1 0 97060 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1068
timestamp 1676037725
transform 1 0 99360 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1079
timestamp 1676037725
transform 1 0 100372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1090
timestamp 1676037725
transform 1 0 101384 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_1093
timestamp 1676037725
transform 1 0 101660 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1099
timestamp 1676037725
transform 1 0 102212 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1121
timestamp 1676037725
transform 1 0 104236 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1128
timestamp 1676037725
transform 1 0 104880 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1135
timestamp 1676037725
transform 1 0 105524 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1146
timestamp 1676037725
transform 1 0 106536 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1149
timestamp 1676037725
transform 1 0 106812 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1158
timestamp 1676037725
transform 1 0 107640 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1169
timestamp 1676037725
transform 1 0 108652 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1173
timestamp 1676037725
transform 1 0 109020 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1195
timestamp 1676037725
transform 1 0 111044 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1202
timestamp 1676037725
transform 1 0 111688 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1205
timestamp 1676037725
transform 1 0 111964 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1210
timestamp 1676037725
transform 1 0 112424 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1217
timestamp 1676037725
transform 1 0 113068 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1224
timestamp 1676037725
transform 1 0 113712 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1233
timestamp 1676037725
transform 1 0 114540 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1258
timestamp 1676037725
transform 1 0 116840 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1261
timestamp 1676037725
transform 1 0 117116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1274
timestamp 1676037725
transform 1 0 118312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1281
timestamp 1676037725
transform 1 0 118956 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_1289
timestamp 1676037725
transform 1 0 119692 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1302
timestamp 1676037725
transform 1 0 120888 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_1313
timestamp 1676037725
transform 1 0 121900 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1317
timestamp 1676037725
transform 1 0 122268 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1326
timestamp 1676037725
transform 1 0 123096 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1338
timestamp 1676037725
transform 1 0 124200 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1350
timestamp 1676037725
transform 1 0 125304 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_1362
timestamp 1676037725
transform 1 0 126408 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1370
timestamp 1676037725
transform 1 0 127144 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1373
timestamp 1676037725
transform 1 0 127420 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1385
timestamp 1676037725
transform 1 0 128524 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1397
timestamp 1676037725
transform 1 0 129628 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1409
timestamp 1676037725
transform 1 0 130732 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_1421
timestamp 1676037725
transform 1 0 131836 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1427
timestamp 1676037725
transform 1 0 132388 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1429
timestamp 1676037725
transform 1 0 132572 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1441
timestamp 1676037725
transform 1 0 133676 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1453
timestamp 1676037725
transform 1 0 134780 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1465
timestamp 1676037725
transform 1 0 135884 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_1477
timestamp 1676037725
transform 1 0 136988 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1483
timestamp 1676037725
transform 1 0 137540 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1485
timestamp 1676037725
transform 1 0 137724 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1489
timestamp 1676037725
transform 1 0 138092 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1511
timestamp 1676037725
transform 1 0 140116 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1536
timestamp 1676037725
transform 1 0 142416 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1541
timestamp 1676037725
transform 1 0 142876 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_1550
timestamp 1676037725
transform 1 0 143704 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_1579
timestamp 1676037725
transform 1 0 146372 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1585
timestamp 1676037725
transform 1 0 146924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_1590
timestamp 1676037725
transform 1 0 147384 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1597
timestamp 1676037725
transform 1 0 148028 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1602
timestamp 1676037725
transform 1 0 148488 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1606
timestamp 1676037725
transform 1 0 148856 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1628
timestamp 1676037725
transform 1 0 150880 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1639
timestamp 1676037725
transform 1 0 151892 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1650
timestamp 1676037725
transform 1 0 152904 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1653
timestamp 1676037725
transform 1 0 153180 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1676
timestamp 1676037725
transform 1 0 155296 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_1701
timestamp 1676037725
transform 1 0 157596 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1707
timestamp 1676037725
transform 1 0 158148 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1709
timestamp 1676037725
transform 1 0 158332 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1732
timestamp 1676037725
transform 1 0 160448 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1744
timestamp 1676037725
transform 1 0 161552 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_1756
timestamp 1676037725
transform 1 0 162656 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1765
timestamp 1676037725
transform 1 0 163484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_1777
timestamp 1676037725
transform 1 0 164588 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1785
timestamp 1676037725
transform 1 0 165324 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1789
timestamp 1676037725
transform 1 0 165692 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1793
timestamp 1676037725
transform 1 0 166060 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1816
timestamp 1676037725
transform 1 0 168176 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1821
timestamp 1676037725
transform 1 0 168636 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1827
timestamp 1676037725
transform 1 0 169188 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1839
timestamp 1676037725
transform 1 0 170292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1851
timestamp 1676037725
transform 1 0 171396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1863
timestamp 1676037725
transform 1 0 172500 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1875
timestamp 1676037725
transform 1 0 173604 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1877
timestamp 1676037725
transform 1 0 173788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1889
timestamp 1676037725
transform 1 0 174892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1901
timestamp 1676037725
transform 1 0 175996 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1913
timestamp 1676037725
transform 1 0 177100 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_1925
timestamp 1676037725
transform 1 0 178204 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1931
timestamp 1676037725
transform 1 0 178756 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1933
timestamp 1676037725
transform 1 0 178940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1945
timestamp 1676037725
transform 1 0 180044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1957
timestamp 1676037725
transform 1 0 181148 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1969
timestamp 1676037725
transform 1 0 182252 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_1981
timestamp 1676037725
transform 1 0 183356 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1987
timestamp 1676037725
transform 1 0 183908 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1989
timestamp 1676037725
transform 1 0 184092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2001
timestamp 1676037725
transform 1 0 185196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2013
timestamp 1676037725
transform 1 0 186300 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2025
timestamp 1676037725
transform 1 0 187404 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_2037
timestamp 1676037725
transform 1 0 188508 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2043
timestamp 1676037725
transform 1 0 189060 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2045
timestamp 1676037725
transform 1 0 189244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2057
timestamp 1676037725
transform 1 0 190348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2069
timestamp 1676037725
transform 1 0 191452 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2081
timestamp 1676037725
transform 1 0 192556 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_2093
timestamp 1676037725
transform 1 0 193660 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2099
timestamp 1676037725
transform 1 0 194212 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2101
timestamp 1676037725
transform 1 0 194396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2113
timestamp 1676037725
transform 1 0 195500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2125
timestamp 1676037725
transform 1 0 196604 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2137
timestamp 1676037725
transform 1 0 197708 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_2149
timestamp 1676037725
transform 1 0 198812 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2155
timestamp 1676037725
transform 1 0 199364 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2157
timestamp 1676037725
transform 1 0 199548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2169
timestamp 1676037725
transform 1 0 200652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2181
timestamp 1676037725
transform 1 0 201756 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2193
timestamp 1676037725
transform 1 0 202860 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_2205
timestamp 1676037725
transform 1 0 203964 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2211
timestamp 1676037725
transform 1 0 204516 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_2213
timestamp 1676037725
transform 1 0 204700 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2221
timestamp 1676037725
transform 1 0 205436 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2228
timestamp 1676037725
transform 1 0 206080 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2253
timestamp 1676037725
transform 1 0 208380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2263
timestamp 1676037725
transform 1 0 209300 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2267
timestamp 1676037725
transform 1 0 209668 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2269
timestamp 1676037725
transform 1 0 209852 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_2277
timestamp 1676037725
transform 1 0 210588 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2285
timestamp 1676037725
transform 1 0 211324 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2295
timestamp 1676037725
transform 1 0 212244 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2299
timestamp 1676037725
transform 1 0 212612 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2322
timestamp 1676037725
transform 1 0 214728 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2325
timestamp 1676037725
transform 1 0 215004 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_2348
timestamp 1676037725
transform 1 0 217120 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2356
timestamp 1676037725
transform 1 0 217856 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2378
timestamp 1676037725
transform 1 0 219880 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2381
timestamp 1676037725
transform 1 0 220156 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2386
timestamp 1676037725
transform 1 0 220616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2390
timestamp 1676037725
transform 1 0 220984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2412
timestamp 1676037725
transform 1 0 223008 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2424
timestamp 1676037725
transform 1 0 224112 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2431
timestamp 1676037725
transform 1 0 224756 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2435
timestamp 1676037725
transform 1 0 225124 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2437
timestamp 1676037725
transform 1 0 225308 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2460
timestamp 1676037725
transform 1 0 227424 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2472
timestamp 1676037725
transform 1 0 228528 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_2484
timestamp 1676037725
transform 1 0 229632 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2493
timestamp 1676037725
transform 1 0 230460 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2505
timestamp 1676037725
transform 1 0 231564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2517
timestamp 1676037725
transform 1 0 232668 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2529
timestamp 1676037725
transform 1 0 233772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_2541
timestamp 1676037725
transform 1 0 234876 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2547
timestamp 1676037725
transform 1 0 235428 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2549
timestamp 1676037725
transform 1 0 235612 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2561
timestamp 1676037725
transform 1 0 236716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2573
timestamp 1676037725
transform 1 0 237820 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2585
timestamp 1676037725
transform 1 0 238924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_2597
timestamp 1676037725
transform 1 0 240028 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2603
timestamp 1676037725
transform 1 0 240580 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2605
timestamp 1676037725
transform 1 0 240764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2617
timestamp 1676037725
transform 1 0 241868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2629
timestamp 1676037725
transform 1 0 242972 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_2641
timestamp 1676037725
transform 1 0 244076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2647
timestamp 1676037725
transform 1 0 244628 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2651
timestamp 1676037725
transform 1 0 244996 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2658
timestamp 1676037725
transform 1 0 245640 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_2661
timestamp 1676037725
transform 1 0 245916 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2675
timestamp 1676037725
transform 1 0 247204 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2689
timestamp 1676037725
transform 1 0 248492 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2714
timestamp 1676037725
transform 1 0 250792 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2717
timestamp 1676037725
transform 1 0 251068 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_2725
timestamp 1676037725
transform 1 0 251804 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2738
timestamp 1676037725
transform 1 0 253000 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2763
timestamp 1676037725
transform 1 0 255300 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2770
timestamp 1676037725
transform 1 0 255944 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2773
timestamp 1676037725
transform 1 0 256220 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2796
timestamp 1676037725
transform 1 0 258336 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2806
timestamp 1676037725
transform 1 0 259256 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2813
timestamp 1676037725
transform 1 0 259900 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_2825
timestamp 1676037725
transform 1 0 261004 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2829
timestamp 1676037725
transform 1 0 261372 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2834
timestamp 1676037725
transform 1 0 261832 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2846
timestamp 1676037725
transform 1 0 262936 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2861
timestamp 1676037725
transform 1 0 264316 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2868
timestamp 1676037725
transform 1 0 264960 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2875
timestamp 1676037725
transform 1 0 265604 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2882
timestamp 1676037725
transform 1 0 266248 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_2885
timestamp 1676037725
transform 1 0 266524 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_2897
timestamp 1676037725
transform 1 0 267628 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2905
timestamp 1676037725
transform 1 0 268364 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2915
timestamp 1676037725
transform 1 0 269284 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2924
timestamp 1676037725
transform 1 0 270112 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2932
timestamp 1676037725
transform 1 0 270848 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1676037725
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1676037725
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1676037725
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1676037725
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1676037725
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_361
timestamp 1676037725
transform 1 0 34316 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_369
timestamp 1676037725
transform 1 0 35052 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_390
timestamp 1676037725
transform 1 0 36984 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1676037725
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_417
timestamp 1676037725
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_429
timestamp 1676037725
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_441
timestamp 1676037725
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 1676037725
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_461
timestamp 1676037725
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_473
timestamp 1676037725
transform 1 0 44620 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_481
timestamp 1676037725
transform 1 0 45356 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_502
timestamp 1676037725
transform 1 0 47288 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_505
timestamp 1676037725
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_517
timestamp 1676037725
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_529
timestamp 1676037725
transform 1 0 49772 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_535
timestamp 1676037725
transform 1 0 50324 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_538
timestamp 1676037725
transform 1 0 50600 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_558
timestamp 1676037725
transform 1 0 52440 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_561
timestamp 1676037725
transform 1 0 52716 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_567
timestamp 1676037725
transform 1 0 53268 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_571
timestamp 1676037725
transform 1 0 53636 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_583
timestamp 1676037725
transform 1 0 54740 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_595
timestamp 1676037725
transform 1 0 55844 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_607
timestamp 1676037725
transform 1 0 56948 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_615
timestamp 1676037725
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_617
timestamp 1676037725
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_629
timestamp 1676037725
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_641
timestamp 1676037725
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_653
timestamp 1676037725
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_665
timestamp 1676037725
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_671
timestamp 1676037725
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_673
timestamp 1676037725
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_685
timestamp 1676037725
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_697
timestamp 1676037725
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_709
timestamp 1676037725
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_721
timestamp 1676037725
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_727
timestamp 1676037725
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_729
timestamp 1676037725
transform 1 0 68172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_741
timestamp 1676037725
transform 1 0 69276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_753
timestamp 1676037725
transform 1 0 70380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_765
timestamp 1676037725
transform 1 0 71484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_777
timestamp 1676037725
transform 1 0 72588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_783
timestamp 1676037725
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_785
timestamp 1676037725
transform 1 0 73324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_797
timestamp 1676037725
transform 1 0 74428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_809
timestamp 1676037725
transform 1 0 75532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_821
timestamp 1676037725
transform 1 0 76636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_833
timestamp 1676037725
transform 1 0 77740 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_839
timestamp 1676037725
transform 1 0 78292 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_841
timestamp 1676037725
transform 1 0 78476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_853
timestamp 1676037725
transform 1 0 79580 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_865
timestamp 1676037725
transform 1 0 80684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_877
timestamp 1676037725
transform 1 0 81788 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_889
timestamp 1676037725
transform 1 0 82892 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_895
timestamp 1676037725
transform 1 0 83444 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_897
timestamp 1676037725
transform 1 0 83628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_909
timestamp 1676037725
transform 1 0 84732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_921
timestamp 1676037725
transform 1 0 85836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_933
timestamp 1676037725
transform 1 0 86940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_945
timestamp 1676037725
transform 1 0 88044 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_951
timestamp 1676037725
transform 1 0 88596 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_953
timestamp 1676037725
transform 1 0 88780 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_965
timestamp 1676037725
transform 1 0 89884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_977
timestamp 1676037725
transform 1 0 90988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_989
timestamp 1676037725
transform 1 0 92092 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1001
timestamp 1676037725
transform 1 0 93196 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1006
timestamp 1676037725
transform 1 0 93656 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1009
timestamp 1676037725
transform 1 0 93932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1034
timestamp 1676037725
transform 1 0 96232 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1059
timestamp 1676037725
transform 1 0 98532 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1063
timestamp 1676037725
transform 1 0 98900 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1065
timestamp 1676037725
transform 1 0 99084 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1074
timestamp 1676037725
transform 1 0 99912 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1085
timestamp 1676037725
transform 1 0 100924 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1096
timestamp 1676037725
transform 1 0 101936 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1105
timestamp 1676037725
transform 1 0 102764 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_1112
timestamp 1676037725
transform 1 0 103408 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_1121
timestamp 1676037725
transform 1 0 104236 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1130
timestamp 1676037725
transform 1 0 105064 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1134
timestamp 1676037725
transform 1 0 105432 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_1142
timestamp 1676037725
transform 1 0 106168 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1150
timestamp 1676037725
transform 1 0 106904 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_1161
timestamp 1676037725
transform 1 0 107916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1167
timestamp 1676037725
transform 1 0 108468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_1173
timestamp 1676037725
transform 1 0 109020 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1177
timestamp 1676037725
transform 1 0 109388 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1188
timestamp 1676037725
transform 1 0 110400 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1213
timestamp 1676037725
transform 1 0 112700 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1217
timestamp 1676037725
transform 1 0 113068 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1221
timestamp 1676037725
transform 1 0 113436 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1230
timestamp 1676037725
transform 1 0 114264 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1233
timestamp 1676037725
transform 1 0 114540 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_1240
timestamp 1676037725
transform 1 0 115184 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1246
timestamp 1676037725
transform 1 0 115736 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1255
timestamp 1676037725
transform 1 0 116564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_1280
timestamp 1676037725
transform 1 0 118864 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1289
timestamp 1676037725
transform 1 0 119692 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1295
timestamp 1676037725
transform 1 0 120244 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1306
timestamp 1676037725
transform 1 0 121256 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1313
timestamp 1676037725
transform 1 0 121900 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1320
timestamp 1676037725
transform 1 0 122544 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1332
timestamp 1676037725
transform 1 0 123648 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1345
timestamp 1676037725
transform 1 0 124844 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1357
timestamp 1676037725
transform 1 0 125948 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1369
timestamp 1676037725
transform 1 0 127052 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1381
timestamp 1676037725
transform 1 0 128156 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_1393
timestamp 1676037725
transform 1 0 129260 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1399
timestamp 1676037725
transform 1 0 129812 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1401
timestamp 1676037725
transform 1 0 129996 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1413
timestamp 1676037725
transform 1 0 131100 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1425
timestamp 1676037725
transform 1 0 132204 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1437
timestamp 1676037725
transform 1 0 133308 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_1449
timestamp 1676037725
transform 1 0 134412 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1455
timestamp 1676037725
transform 1 0 134964 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1457
timestamp 1676037725
transform 1 0 135148 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1469
timestamp 1676037725
transform 1 0 136252 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1481
timestamp 1676037725
transform 1 0 137356 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_1489
timestamp 1676037725
transform 1 0 138092 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1499
timestamp 1676037725
transform 1 0 139012 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1510
timestamp 1676037725
transform 1 0 140024 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1513
timestamp 1676037725
transform 1 0 140300 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_1525
timestamp 1676037725
transform 1 0 141404 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1540
timestamp 1676037725
transform 1 0 142784 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1551
timestamp 1676037725
transform 1 0 143796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1558
timestamp 1676037725
transform 1 0 144440 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_1565
timestamp 1676037725
transform 1 0 145084 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1569
timestamp 1676037725
transform 1 0 145452 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_1592
timestamp 1676037725
transform 1 0 147568 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1598
timestamp 1676037725
transform 1 0 148120 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_1606
timestamp 1676037725
transform 1 0 148856 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1614
timestamp 1676037725
transform 1 0 149592 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1622
timestamp 1676037725
transform 1 0 150328 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1625
timestamp 1676037725
transform 1 0 150604 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1648
timestamp 1676037725
transform 1 0 152720 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_1673
timestamp 1676037725
transform 1 0 155020 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1679
timestamp 1676037725
transform 1 0 155572 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1681
timestamp 1676037725
transform 1 0 155756 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1704
timestamp 1676037725
transform 1 0 157872 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1716
timestamp 1676037725
transform 1 0 158976 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_1728
timestamp 1676037725
transform 1 0 160080 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1737
timestamp 1676037725
transform 1 0 160908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1749
timestamp 1676037725
transform 1 0 162012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1761
timestamp 1676037725
transform 1 0 163116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1773
timestamp 1676037725
transform 1 0 164220 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_1785
timestamp 1676037725
transform 1 0 165324 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1791
timestamp 1676037725
transform 1 0 165876 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1793
timestamp 1676037725
transform 1 0 166060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_1805
timestamp 1676037725
transform 1 0 167164 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1813
timestamp 1676037725
transform 1 0 167900 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1836
timestamp 1676037725
transform 1 0 170016 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1849
timestamp 1676037725
transform 1 0 171212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1861
timestamp 1676037725
transform 1 0 172316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1873
timestamp 1676037725
transform 1 0 173420 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1885
timestamp 1676037725
transform 1 0 174524 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_1897
timestamp 1676037725
transform 1 0 175628 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1903
timestamp 1676037725
transform 1 0 176180 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1905
timestamp 1676037725
transform 1 0 176364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1917
timestamp 1676037725
transform 1 0 177468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1929
timestamp 1676037725
transform 1 0 178572 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1941
timestamp 1676037725
transform 1 0 179676 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_1953
timestamp 1676037725
transform 1 0 180780 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1959
timestamp 1676037725
transform 1 0 181332 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1961
timestamp 1676037725
transform 1 0 181516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1973
timestamp 1676037725
transform 1 0 182620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1985
timestamp 1676037725
transform 1 0 183724 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1997
timestamp 1676037725
transform 1 0 184828 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2009
timestamp 1676037725
transform 1 0 185932 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2015
timestamp 1676037725
transform 1 0 186484 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2017
timestamp 1676037725
transform 1 0 186668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2029
timestamp 1676037725
transform 1 0 187772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2041
timestamp 1676037725
transform 1 0 188876 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2053
timestamp 1676037725
transform 1 0 189980 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2065
timestamp 1676037725
transform 1 0 191084 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2071
timestamp 1676037725
transform 1 0 191636 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2073
timestamp 1676037725
transform 1 0 191820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2085
timestamp 1676037725
transform 1 0 192924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2097
timestamp 1676037725
transform 1 0 194028 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2109
timestamp 1676037725
transform 1 0 195132 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2121
timestamp 1676037725
transform 1 0 196236 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2127
timestamp 1676037725
transform 1 0 196788 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2129
timestamp 1676037725
transform 1 0 196972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2141
timestamp 1676037725
transform 1 0 198076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2153
timestamp 1676037725
transform 1 0 199180 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2165
timestamp 1676037725
transform 1 0 200284 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2177
timestamp 1676037725
transform 1 0 201388 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2183
timestamp 1676037725
transform 1 0 201940 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2185
timestamp 1676037725
transform 1 0 202124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2197
timestamp 1676037725
transform 1 0 203228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2209
timestamp 1676037725
transform 1 0 204332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_2221
timestamp 1676037725
transform 1 0 205436 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_2229
timestamp 1676037725
transform 1 0 206172 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2238
timestamp 1676037725
transform 1 0 207000 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2241
timestamp 1676037725
transform 1 0 207276 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2264
timestamp 1676037725
transform 1 0 209392 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2274
timestamp 1676037725
transform 1 0 210312 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_2286
timestamp 1676037725
transform 1 0 211416 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2294
timestamp 1676037725
transform 1 0 212152 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2297
timestamp 1676037725
transform 1 0 212428 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2303
timestamp 1676037725
transform 1 0 212980 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2306
timestamp 1676037725
transform 1 0 213256 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2329
timestamp 1676037725
transform 1 0 215372 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2342
timestamp 1676037725
transform 1 0 216568 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_2349
timestamp 1676037725
transform 1 0 217212 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_2353
timestamp 1676037725
transform 1 0 217580 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2377
timestamp 1676037725
transform 1 0 219788 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2402
timestamp 1676037725
transform 1 0 222088 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2409
timestamp 1676037725
transform 1 0 222732 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2432
timestamp 1676037725
transform 1 0 224848 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2457
timestamp 1676037725
transform 1 0 227148 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2463
timestamp 1676037725
transform 1 0 227700 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2465
timestamp 1676037725
transform 1 0 227884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2477
timestamp 1676037725
transform 1 0 228988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2489
timestamp 1676037725
transform 1 0 230092 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2501
timestamp 1676037725
transform 1 0 231196 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2513
timestamp 1676037725
transform 1 0 232300 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2519
timestamp 1676037725
transform 1 0 232852 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2521
timestamp 1676037725
transform 1 0 233036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2533
timestamp 1676037725
transform 1 0 234140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2545
timestamp 1676037725
transform 1 0 235244 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2557
timestamp 1676037725
transform 1 0 236348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2569
timestamp 1676037725
transform 1 0 237452 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2575
timestamp 1676037725
transform 1 0 238004 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2577
timestamp 1676037725
transform 1 0 238188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2589
timestamp 1676037725
transform 1 0 239292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2601
timestamp 1676037725
transform 1 0 240396 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2613
timestamp 1676037725
transform 1 0 241500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2625
timestamp 1676037725
transform 1 0 242604 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2631
timestamp 1676037725
transform 1 0 243156 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2633
timestamp 1676037725
transform 1 0 243340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2645
timestamp 1676037725
transform 1 0 244444 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2657
timestamp 1676037725
transform 1 0 245548 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2664
timestamp 1676037725
transform 1 0 246192 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2676
timestamp 1676037725
transform 1 0 247296 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2686
timestamp 1676037725
transform 1 0 248216 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2689
timestamp 1676037725
transform 1 0 248492 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2712
timestamp 1676037725
transform 1 0 250608 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2720
timestamp 1676037725
transform 1 0 251344 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2727
timestamp 1676037725
transform 1 0 251988 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2742
timestamp 1676037725
transform 1 0 253368 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2745
timestamp 1676037725
transform 1 0 253644 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2757
timestamp 1676037725
transform 1 0 254748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2782
timestamp 1676037725
transform 1 0 257048 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_2792
timestamp 1676037725
transform 1 0 257968 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_2801
timestamp 1676037725
transform 1 0 258796 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2809
timestamp 1676037725
transform 1 0 259532 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2820
timestamp 1676037725
transform 1 0 260544 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2833
timestamp 1676037725
transform 1 0 261740 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_2842
timestamp 1676037725
transform 1 0 262568 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2850
timestamp 1676037725
transform 1 0 263304 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2854
timestamp 1676037725
transform 1 0 263672 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2857
timestamp 1676037725
transform 1 0 263948 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2861
timestamp 1676037725
transform 1 0 264316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2865
timestamp 1676037725
transform 1 0 264684 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2872
timestamp 1676037725
transform 1 0 265328 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2880
timestamp 1676037725
transform 1 0 266064 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2889
timestamp 1676037725
transform 1 0 266892 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2893
timestamp 1676037725
transform 1 0 267260 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2899
timestamp 1676037725
transform 1 0 267812 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2908
timestamp 1676037725
transform 1 0 268640 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2913
timestamp 1676037725
transform 1 0 269100 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2920
timestamp 1676037725
transform 1 0 269744 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2929
timestamp 1676037725
transform 1 0 270572 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2935
timestamp 1676037725
transform 1 0 271124 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1676037725
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1676037725
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1676037725
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1676037725
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1676037725
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1676037725
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1676037725
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1676037725
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1676037725
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1676037725
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_401
timestamp 1676037725
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_413
timestamp 1676037725
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 1676037725
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 1676037725
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 1676037725
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_457
timestamp 1676037725
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_469
timestamp 1676037725
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_475
timestamp 1676037725
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_477
timestamp 1676037725
transform 1 0 44988 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_497
timestamp 1676037725
transform 1 0 46828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_507
timestamp 1676037725
transform 1 0 47748 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_515
timestamp 1676037725
transform 1 0 48484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_527
timestamp 1676037725
transform 1 0 49588 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_531
timestamp 1676037725
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_533
timestamp 1676037725
transform 1 0 50140 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_541
timestamp 1676037725
transform 1 0 50876 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_545
timestamp 1676037725
transform 1 0 51244 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_549
timestamp 1676037725
transform 1 0 51612 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_569
timestamp 1676037725
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_581
timestamp 1676037725
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_587
timestamp 1676037725
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_589
timestamp 1676037725
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_601
timestamp 1676037725
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_613
timestamp 1676037725
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_625
timestamp 1676037725
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_637
timestamp 1676037725
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_643
timestamp 1676037725
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_645
timestamp 1676037725
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_657
timestamp 1676037725
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_669
timestamp 1676037725
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_681
timestamp 1676037725
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_693
timestamp 1676037725
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_699
timestamp 1676037725
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_701
timestamp 1676037725
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_713
timestamp 1676037725
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_725
timestamp 1676037725
transform 1 0 67804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_737
timestamp 1676037725
transform 1 0 68908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_749
timestamp 1676037725
transform 1 0 70012 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_755
timestamp 1676037725
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_757
timestamp 1676037725
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_769
timestamp 1676037725
transform 1 0 71852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_781
timestamp 1676037725
transform 1 0 72956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_793
timestamp 1676037725
transform 1 0 74060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_805
timestamp 1676037725
transform 1 0 75164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_811
timestamp 1676037725
transform 1 0 75716 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_813
timestamp 1676037725
transform 1 0 75900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_825
timestamp 1676037725
transform 1 0 77004 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_837
timestamp 1676037725
transform 1 0 78108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_849
timestamp 1676037725
transform 1 0 79212 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_861
timestamp 1676037725
transform 1 0 80316 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_867
timestamp 1676037725
transform 1 0 80868 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_869
timestamp 1676037725
transform 1 0 81052 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_881
timestamp 1676037725
transform 1 0 82156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_893
timestamp 1676037725
transform 1 0 83260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_905
timestamp 1676037725
transform 1 0 84364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_917
timestamp 1676037725
transform 1 0 85468 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_923
timestamp 1676037725
transform 1 0 86020 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_925
timestamp 1676037725
transform 1 0 86204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_937
timestamp 1676037725
transform 1 0 87308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_949
timestamp 1676037725
transform 1 0 88412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_961
timestamp 1676037725
transform 1 0 89516 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_973
timestamp 1676037725
transform 1 0 90620 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_979
timestamp 1676037725
transform 1 0 91172 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_981
timestamp 1676037725
transform 1 0 91356 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_993
timestamp 1676037725
transform 1 0 92460 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_1005
timestamp 1676037725
transform 1 0 93564 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1013
timestamp 1676037725
transform 1 0 94300 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1018
timestamp 1676037725
transform 1 0 94760 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1025
timestamp 1676037725
transform 1 0 95404 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1034
timestamp 1676037725
transform 1 0 96232 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1037
timestamp 1676037725
transform 1 0 96508 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1044
timestamp 1676037725
transform 1 0 97152 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1069
timestamp 1676037725
transform 1 0 99452 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1080
timestamp 1676037725
transform 1 0 100464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1084
timestamp 1676037725
transform 1 0 100832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1090
timestamp 1676037725
transform 1 0 101384 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1093
timestamp 1676037725
transform 1 0 101660 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1100
timestamp 1676037725
transform 1 0 102304 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1108
timestamp 1676037725
transform 1 0 103040 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_1115
timestamp 1676037725
transform 1 0 103684 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1121
timestamp 1676037725
transform 1 0 104236 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1125
timestamp 1676037725
transform 1 0 104604 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1132
timestamp 1676037725
transform 1 0 105248 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1139
timestamp 1676037725
transform 1 0 105892 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1146
timestamp 1676037725
transform 1 0 106536 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_1149
timestamp 1676037725
transform 1 0 106812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1159
timestamp 1676037725
transform 1 0 107732 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1169
timestamp 1676037725
transform 1 0 108652 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1194
timestamp 1676037725
transform 1 0 110952 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1202
timestamp 1676037725
transform 1 0 111688 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1205
timestamp 1676037725
transform 1 0 111964 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_1213
timestamp 1676037725
transform 1 0 112700 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1226
timestamp 1676037725
transform 1 0 113896 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1235
timestamp 1676037725
transform 1 0 114724 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1248
timestamp 1676037725
transform 1 0 115920 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1252
timestamp 1676037725
transform 1 0 116288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1258
timestamp 1676037725
transform 1 0 116840 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1261
timestamp 1676037725
transform 1 0 117116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1284
timestamp 1676037725
transform 1 0 119232 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1296
timestamp 1676037725
transform 1 0 120336 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1300
timestamp 1676037725
transform 1 0 120704 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1304
timestamp 1676037725
transform 1 0 121072 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1314
timestamp 1676037725
transform 1 0 121992 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1317
timestamp 1676037725
transform 1 0 122268 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1329
timestamp 1676037725
transform 1 0 123372 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1341
timestamp 1676037725
transform 1 0 124476 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1353
timestamp 1676037725
transform 1 0 125580 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_1365
timestamp 1676037725
transform 1 0 126684 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1371
timestamp 1676037725
transform 1 0 127236 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1373
timestamp 1676037725
transform 1 0 127420 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1381
timestamp 1676037725
transform 1 0 128156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1393
timestamp 1676037725
transform 1 0 129260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1405
timestamp 1676037725
transform 1 0 130364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_1417
timestamp 1676037725
transform 1 0 131468 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_1425
timestamp 1676037725
transform 1 0 132204 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1429
timestamp 1676037725
transform 1 0 132572 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1437
timestamp 1676037725
transform 1 0 133308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1449
timestamp 1676037725
transform 1 0 134412 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_1461
timestamp 1676037725
transform 1 0 135516 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1471
timestamp 1676037725
transform 1 0 136436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1483
timestamp 1676037725
transform 1 0 137540 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1485
timestamp 1676037725
transform 1 0 137724 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1497
timestamp 1676037725
transform 1 0 138828 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1501
timestamp 1676037725
transform 1 0 139196 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1505
timestamp 1676037725
transform 1 0 139564 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1512
timestamp 1676037725
transform 1 0 140208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_1537
timestamp 1676037725
transform 1 0 142508 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1541
timestamp 1676037725
transform 1 0 142876 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_1546
timestamp 1676037725
transform 1 0 143336 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1565
timestamp 1676037725
transform 1 0 145084 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1575
timestamp 1676037725
transform 1 0 146004 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1579
timestamp 1676037725
transform 1 0 146372 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_1590
timestamp 1676037725
transform 1 0 147384 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1597
timestamp 1676037725
transform 1 0 148028 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1606
timestamp 1676037725
transform 1 0 148856 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1610
timestamp 1676037725
transform 1 0 149224 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1614
timestamp 1676037725
transform 1 0 149592 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1625
timestamp 1676037725
transform 1 0 150604 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1650
timestamp 1676037725
transform 1 0 152904 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_1653
timestamp 1676037725
transform 1 0 153180 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1680
timestamp 1676037725
transform 1 0 155664 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1684
timestamp 1676037725
transform 1 0 156032 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1704
timestamp 1676037725
transform 1 0 157872 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1709
timestamp 1676037725
transform 1 0 158332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1721
timestamp 1676037725
transform 1 0 159436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1733
timestamp 1676037725
transform 1 0 160540 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1745
timestamp 1676037725
transform 1 0 161644 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_1757
timestamp 1676037725
transform 1 0 162748 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1763
timestamp 1676037725
transform 1 0 163300 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1765
timestamp 1676037725
transform 1 0 163484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1777
timestamp 1676037725
transform 1 0 164588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1789
timestamp 1676037725
transform 1 0 165692 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1801
timestamp 1676037725
transform 1 0 166796 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1813
timestamp 1676037725
transform 1 0 167900 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1818
timestamp 1676037725
transform 1 0 168360 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1821
timestamp 1676037725
transform 1 0 168636 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1830
timestamp 1676037725
transform 1 0 169464 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1837
timestamp 1676037725
transform 1 0 170108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1849
timestamp 1676037725
transform 1 0 171212 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1861
timestamp 1676037725
transform 1 0 172316 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_1873
timestamp 1676037725
transform 1 0 173420 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1877
timestamp 1676037725
transform 1 0 173788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1889
timestamp 1676037725
transform 1 0 174892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1901
timestamp 1676037725
transform 1 0 175996 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1913
timestamp 1676037725
transform 1 0 177100 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_1925
timestamp 1676037725
transform 1 0 178204 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1931
timestamp 1676037725
transform 1 0 178756 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1933
timestamp 1676037725
transform 1 0 178940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1945
timestamp 1676037725
transform 1 0 180044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1957
timestamp 1676037725
transform 1 0 181148 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1969
timestamp 1676037725
transform 1 0 182252 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_1981
timestamp 1676037725
transform 1 0 183356 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1987
timestamp 1676037725
transform 1 0 183908 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1989
timestamp 1676037725
transform 1 0 184092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2001
timestamp 1676037725
transform 1 0 185196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2013
timestamp 1676037725
transform 1 0 186300 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2025
timestamp 1676037725
transform 1 0 187404 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_2037
timestamp 1676037725
transform 1 0 188508 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2042
timestamp 1676037725
transform 1 0 188968 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2045
timestamp 1676037725
transform 1 0 189244 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2055
timestamp 1676037725
transform 1 0 190164 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2059
timestamp 1676037725
transform 1 0 190532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2071
timestamp 1676037725
transform 1 0 191636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2083
timestamp 1676037725
transform 1 0 192740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2095
timestamp 1676037725
transform 1 0 193844 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2099
timestamp 1676037725
transform 1 0 194212 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2101
timestamp 1676037725
transform 1 0 194396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2113
timestamp 1676037725
transform 1 0 195500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2125
timestamp 1676037725
transform 1 0 196604 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2137
timestamp 1676037725
transform 1 0 197708 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_2149
timestamp 1676037725
transform 1 0 198812 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2155
timestamp 1676037725
transform 1 0 199364 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2157
timestamp 1676037725
transform 1 0 199548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2169
timestamp 1676037725
transform 1 0 200652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2181
timestamp 1676037725
transform 1 0 201756 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2193
timestamp 1676037725
transform 1 0 202860 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_2205
timestamp 1676037725
transform 1 0 203964 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2211
timestamp 1676037725
transform 1 0 204516 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2213
timestamp 1676037725
transform 1 0 204700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2225
timestamp 1676037725
transform 1 0 205804 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2237
timestamp 1676037725
transform 1 0 206908 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_2262
timestamp 1676037725
transform 1 0 209208 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2269
timestamp 1676037725
transform 1 0 209852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2281
timestamp 1676037725
transform 1 0 210956 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_2293
timestamp 1676037725
transform 1 0 212060 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2299
timestamp 1676037725
transform 1 0 212612 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_2316
timestamp 1676037725
transform 1 0 214176 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2325
timestamp 1676037725
transform 1 0 215004 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_2330
timestamp 1676037725
transform 1 0 215464 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2338
timestamp 1676037725
transform 1 0 216200 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2342
timestamp 1676037725
transform 1 0 216568 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_2352
timestamp 1676037725
transform 1 0 217488 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2358
timestamp 1676037725
transform 1 0 218040 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2368
timestamp 1676037725
transform 1 0 218960 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2381
timestamp 1676037725
transform 1 0 220156 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_2404
timestamp 1676037725
transform 1 0 222272 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2412
timestamp 1676037725
transform 1 0 223008 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2434
timestamp 1676037725
transform 1 0 225032 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2437
timestamp 1676037725
transform 1 0 225308 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2443
timestamp 1676037725
transform 1 0 225860 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2455
timestamp 1676037725
transform 1 0 226964 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2467
timestamp 1676037725
transform 1 0 228068 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2479
timestamp 1676037725
transform 1 0 229172 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2491
timestamp 1676037725
transform 1 0 230276 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2493
timestamp 1676037725
transform 1 0 230460 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2505
timestamp 1676037725
transform 1 0 231564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2517
timestamp 1676037725
transform 1 0 232668 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2529
timestamp 1676037725
transform 1 0 233772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_2541
timestamp 1676037725
transform 1 0 234876 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2547
timestamp 1676037725
transform 1 0 235428 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2549
timestamp 1676037725
transform 1 0 235612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2561
timestamp 1676037725
transform 1 0 236716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2573
timestamp 1676037725
transform 1 0 237820 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2585
timestamp 1676037725
transform 1 0 238924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_2597
timestamp 1676037725
transform 1 0 240028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2603
timestamp 1676037725
transform 1 0 240580 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2605
timestamp 1676037725
transform 1 0 240764 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2617
timestamp 1676037725
transform 1 0 241868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2629
timestamp 1676037725
transform 1 0 242972 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2641
timestamp 1676037725
transform 1 0 244076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_2653
timestamp 1676037725
transform 1 0 245180 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2659
timestamp 1676037725
transform 1 0 245732 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2661
timestamp 1676037725
transform 1 0 245916 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2673
timestamp 1676037725
transform 1 0 247020 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2677
timestamp 1676037725
transform 1 0 247388 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2687
timestamp 1676037725
transform 1 0 248308 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2697
timestamp 1676037725
transform 1 0 249228 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2707
timestamp 1676037725
transform 1 0 250148 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2714
timestamp 1676037725
transform 1 0 250792 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2717
timestamp 1676037725
transform 1 0 251068 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2729
timestamp 1676037725
transform 1 0 252172 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2741
timestamp 1676037725
transform 1 0 253276 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2748
timestamp 1676037725
transform 1 0 253920 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2756
timestamp 1676037725
transform 1 0 254656 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2770
timestamp 1676037725
transform 1 0 255944 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2773
timestamp 1676037725
transform 1 0 256220 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2785
timestamp 1676037725
transform 1 0 257324 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2792
timestamp 1676037725
transform 1 0 257968 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2804
timestamp 1676037725
transform 1 0 259072 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2812
timestamp 1676037725
transform 1 0 259808 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2816
timestamp 1676037725
transform 1 0 260176 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2826
timestamp 1676037725
transform 1 0 261096 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2829
timestamp 1676037725
transform 1 0 261372 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2840
timestamp 1676037725
transform 1 0 262384 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2849
timestamp 1676037725
transform 1 0 263212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2853
timestamp 1676037725
transform 1 0 263580 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2863
timestamp 1676037725
transform 1 0 264500 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2872
timestamp 1676037725
transform 1 0 265328 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2879
timestamp 1676037725
transform 1 0 265972 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2883
timestamp 1676037725
transform 1 0 266340 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_2885
timestamp 1676037725
transform 1 0 266524 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_2897
timestamp 1676037725
transform 1 0 267628 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2903
timestamp 1676037725
transform 1 0 268180 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2913
timestamp 1676037725
transform 1 0 269100 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2922
timestamp 1676037725
transform 1 0 269928 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_2930
timestamp 1676037725
transform 1 0 270664 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1676037725
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1676037725
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1676037725
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1676037725
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 1676037725
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_405
timestamp 1676037725
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_417
timestamp 1676037725
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_429
timestamp 1676037725
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_441
timestamp 1676037725
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_447
timestamp 1676037725
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_461
timestamp 1676037725
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_473
timestamp 1676037725
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_485
timestamp 1676037725
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_497
timestamp 1676037725
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_503
timestamp 1676037725
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_505
timestamp 1676037725
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_517
timestamp 1676037725
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_529
timestamp 1676037725
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_541
timestamp 1676037725
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_553
timestamp 1676037725
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_559
timestamp 1676037725
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_561
timestamp 1676037725
transform 1 0 52716 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_569
timestamp 1676037725
transform 1 0 53452 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_573
timestamp 1676037725
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_585
timestamp 1676037725
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_597
timestamp 1676037725
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_609
timestamp 1676037725
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_615
timestamp 1676037725
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_617
timestamp 1676037725
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_629
timestamp 1676037725
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_641
timestamp 1676037725
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_653
timestamp 1676037725
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_665
timestamp 1676037725
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_671
timestamp 1676037725
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_673
timestamp 1676037725
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_685
timestamp 1676037725
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_697
timestamp 1676037725
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_709
timestamp 1676037725
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_721
timestamp 1676037725
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_727
timestamp 1676037725
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_729
timestamp 1676037725
transform 1 0 68172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_741
timestamp 1676037725
transform 1 0 69276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_753
timestamp 1676037725
transform 1 0 70380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_765
timestamp 1676037725
transform 1 0 71484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_777
timestamp 1676037725
transform 1 0 72588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_783
timestamp 1676037725
transform 1 0 73140 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_785
timestamp 1676037725
transform 1 0 73324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_797
timestamp 1676037725
transform 1 0 74428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_809
timestamp 1676037725
transform 1 0 75532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_821
timestamp 1676037725
transform 1 0 76636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_833
timestamp 1676037725
transform 1 0 77740 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_839
timestamp 1676037725
transform 1 0 78292 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_841
timestamp 1676037725
transform 1 0 78476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_853
timestamp 1676037725
transform 1 0 79580 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_865
timestamp 1676037725
transform 1 0 80684 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_877
timestamp 1676037725
transform 1 0 81788 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_889
timestamp 1676037725
transform 1 0 82892 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_895
timestamp 1676037725
transform 1 0 83444 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_897
timestamp 1676037725
transform 1 0 83628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_909
timestamp 1676037725
transform 1 0 84732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_921
timestamp 1676037725
transform 1 0 85836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_933
timestamp 1676037725
transform 1 0 86940 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_945
timestamp 1676037725
transform 1 0 88044 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_951
timestamp 1676037725
transform 1 0 88596 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_953
timestamp 1676037725
transform 1 0 88780 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_965
timestamp 1676037725
transform 1 0 89884 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_977
timestamp 1676037725
transform 1 0 90988 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_1006
timestamp 1676037725
transform 1 0 93656 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_1009
timestamp 1676037725
transform 1 0 93932 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1020
timestamp 1676037725
transform 1 0 94944 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1045
timestamp 1676037725
transform 1 0 97244 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1049
timestamp 1676037725
transform 1 0 97612 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1053
timestamp 1676037725
transform 1 0 97980 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_1062
timestamp 1676037725
transform 1 0 98808 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1065
timestamp 1676037725
transform 1 0 99084 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1076
timestamp 1676037725
transform 1 0 100096 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1083
timestamp 1676037725
transform 1 0 100740 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1092
timestamp 1676037725
transform 1 0 101568 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1101
timestamp 1676037725
transform 1 0 102396 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1109
timestamp 1676037725
transform 1 0 103132 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1116
timestamp 1676037725
transform 1 0 103776 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_1121
timestamp 1676037725
transform 1 0 104236 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_1126
timestamp 1676037725
transform 1 0 104696 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1137
timestamp 1676037725
transform 1 0 105708 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_1144
timestamp 1676037725
transform 1 0 106352 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1150
timestamp 1676037725
transform 1 0 106904 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1155
timestamp 1676037725
transform 1 0 107364 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1164
timestamp 1676037725
transform 1 0 108192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_1173
timestamp 1676037725
transform 1 0 109020 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_1177
timestamp 1676037725
transform 1 0 109388 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1200
timestamp 1676037725
transform 1 0 111504 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_1207
timestamp 1676037725
transform 1 0 112148 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1213
timestamp 1676037725
transform 1 0 112700 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1217
timestamp 1676037725
transform 1 0 113068 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1228
timestamp 1676037725
transform 1 0 114080 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1233
timestamp 1676037725
transform 1 0 114540 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1237
timestamp 1676037725
transform 1 0 114908 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_1259
timestamp 1676037725
transform 1 0 116932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1265
timestamp 1676037725
transform 1 0 117484 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1273
timestamp 1676037725
transform 1 0 118220 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1284
timestamp 1676037725
transform 1 0 119232 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1289
timestamp 1676037725
transform 1 0 119692 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1301
timestamp 1676037725
transform 1 0 120796 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1313
timestamp 1676037725
transform 1 0 121900 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1325
timestamp 1676037725
transform 1 0 123004 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_1337
timestamp 1676037725
transform 1 0 124108 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1343
timestamp 1676037725
transform 1 0 124660 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1345
timestamp 1676037725
transform 1 0 124844 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1357
timestamp 1676037725
transform 1 0 125948 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1369
timestamp 1676037725
transform 1 0 127052 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1381
timestamp 1676037725
transform 1 0 128156 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_1393
timestamp 1676037725
transform 1 0 129260 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1399
timestamp 1676037725
transform 1 0 129812 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1401
timestamp 1676037725
transform 1 0 129996 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1413
timestamp 1676037725
transform 1 0 131100 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1425
timestamp 1676037725
transform 1 0 132204 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1437
timestamp 1676037725
transform 1 0 133308 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_1449
timestamp 1676037725
transform 1 0 134412 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1455
timestamp 1676037725
transform 1 0 134964 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_1457
timestamp 1676037725
transform 1 0 135148 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1465
timestamp 1676037725
transform 1 0 135884 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1483
timestamp 1676037725
transform 1 0 137540 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1495
timestamp 1676037725
transform 1 0 138644 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1507
timestamp 1676037725
transform 1 0 139748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1511
timestamp 1676037725
transform 1 0 140116 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_1513
timestamp 1676037725
transform 1 0 140300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1521
timestamp 1676037725
transform 1 0 141036 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1529
timestamp 1676037725
transform 1 0 141772 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1537
timestamp 1676037725
transform 1 0 142508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1549
timestamp 1676037725
transform 1 0 143612 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_1561
timestamp 1676037725
transform 1 0 144716 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1567
timestamp 1676037725
transform 1 0 145268 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1569
timestamp 1676037725
transform 1 0 145452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1581
timestamp 1676037725
transform 1 0 146556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1593
timestamp 1676037725
transform 1 0 147660 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1605
timestamp 1676037725
transform 1 0 148764 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_1617
timestamp 1676037725
transform 1 0 149868 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_1622
timestamp 1676037725
transform 1 0 150328 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_1625
timestamp 1676037725
transform 1 0 150604 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1634
timestamp 1676037725
transform 1 0 151432 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1645
timestamp 1676037725
transform 1 0 152444 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1655
timestamp 1676037725
transform 1 0 153364 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1665
timestamp 1676037725
transform 1 0 154284 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_1672
timestamp 1676037725
transform 1 0 154928 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_1681
timestamp 1676037725
transform 1 0 155756 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1686
timestamp 1676037725
transform 1 0 156216 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1698
timestamp 1676037725
transform 1 0 157320 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1710
timestamp 1676037725
transform 1 0 158424 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1722
timestamp 1676037725
transform 1 0 159528 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_1734
timestamp 1676037725
transform 1 0 160632 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1737
timestamp 1676037725
transform 1 0 160908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1749
timestamp 1676037725
transform 1 0 162012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1761
timestamp 1676037725
transform 1 0 163116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1773
timestamp 1676037725
transform 1 0 164220 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_1785
timestamp 1676037725
transform 1 0 165324 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1791
timestamp 1676037725
transform 1 0 165876 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1793
timestamp 1676037725
transform 1 0 166060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1805
timestamp 1676037725
transform 1 0 167164 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1809
timestamp 1676037725
transform 1 0 167532 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_1812
timestamp 1676037725
transform 1 0 167808 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_1816
timestamp 1676037725
transform 1 0 168176 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1826
timestamp 1676037725
transform 1 0 169096 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1836
timestamp 1676037725
transform 1 0 170016 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1849
timestamp 1676037725
transform 1 0 171212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1861
timestamp 1676037725
transform 1 0 172316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1873
timestamp 1676037725
transform 1 0 173420 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1885
timestamp 1676037725
transform 1 0 174524 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_1897
timestamp 1676037725
transform 1 0 175628 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1903
timestamp 1676037725
transform 1 0 176180 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1905
timestamp 1676037725
transform 1 0 176364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1917
timestamp 1676037725
transform 1 0 177468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1929
timestamp 1676037725
transform 1 0 178572 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1941
timestamp 1676037725
transform 1 0 179676 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_1953
timestamp 1676037725
transform 1 0 180780 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1959
timestamp 1676037725
transform 1 0 181332 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1961
timestamp 1676037725
transform 1 0 181516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1973
timestamp 1676037725
transform 1 0 182620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1985
timestamp 1676037725
transform 1 0 183724 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1997
timestamp 1676037725
transform 1 0 184828 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_2009
timestamp 1676037725
transform 1 0 185932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2015
timestamp 1676037725
transform 1 0 186484 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2017
timestamp 1676037725
transform 1 0 186668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_2029
timestamp 1676037725
transform 1 0 187772 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_2037
timestamp 1676037725
transform 1 0 188508 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2042
timestamp 1676037725
transform 1 0 188968 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2051
timestamp 1676037725
transform 1 0 189796 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2055
timestamp 1676037725
transform 1 0 190164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2067
timestamp 1676037725
transform 1 0 191268 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2071
timestamp 1676037725
transform 1 0 191636 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2073
timestamp 1676037725
transform 1 0 191820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2085
timestamp 1676037725
transform 1 0 192924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2097
timestamp 1676037725
transform 1 0 194028 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2109
timestamp 1676037725
transform 1 0 195132 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_2121
timestamp 1676037725
transform 1 0 196236 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2127
timestamp 1676037725
transform 1 0 196788 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2129
timestamp 1676037725
transform 1 0 196972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2141
timestamp 1676037725
transform 1 0 198076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2153
timestamp 1676037725
transform 1 0 199180 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2165
timestamp 1676037725
transform 1 0 200284 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_2177
timestamp 1676037725
transform 1 0 201388 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2183
timestamp 1676037725
transform 1 0 201940 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2185
timestamp 1676037725
transform 1 0 202124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2197
timestamp 1676037725
transform 1 0 203228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2209
timestamp 1676037725
transform 1 0 204332 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2221
timestamp 1676037725
transform 1 0 205436 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_2233
timestamp 1676037725
transform 1 0 206540 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2239
timestamp 1676037725
transform 1 0 207092 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_2241
timestamp 1676037725
transform 1 0 207276 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2249
timestamp 1676037725
transform 1 0 208012 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2272
timestamp 1676037725
transform 1 0 210128 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2284
timestamp 1676037725
transform 1 0 211232 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2297
timestamp 1676037725
transform 1 0 212428 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2301
timestamp 1676037725
transform 1 0 212796 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2314
timestamp 1676037725
transform 1 0 213992 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_2326
timestamp 1676037725
transform 1 0 215096 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2332
timestamp 1676037725
transform 1 0 215648 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2335
timestamp 1676037725
transform 1 0 215924 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2345
timestamp 1676037725
transform 1 0 216844 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_2349
timestamp 1676037725
transform 1 0 217212 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2353
timestamp 1676037725
transform 1 0 217580 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2361
timestamp 1676037725
transform 1 0 218316 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2365
timestamp 1676037725
transform 1 0 218684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_2387
timestamp 1676037725
transform 1 0 220708 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2395
timestamp 1676037725
transform 1 0 221444 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_2402
timestamp 1676037725
transform 1 0 222088 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2430
timestamp 1676037725
transform 1 0 224664 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2434
timestamp 1676037725
transform 1 0 225032 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_2457
timestamp 1676037725
transform 1 0 227148 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2463
timestamp 1676037725
transform 1 0 227700 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2465
timestamp 1676037725
transform 1 0 227884 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2477
timestamp 1676037725
transform 1 0 228988 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2489
timestamp 1676037725
transform 1 0 230092 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2501
timestamp 1676037725
transform 1 0 231196 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_2513
timestamp 1676037725
transform 1 0 232300 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2519
timestamp 1676037725
transform 1 0 232852 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2521
timestamp 1676037725
transform 1 0 233036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2533
timestamp 1676037725
transform 1 0 234140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2545
timestamp 1676037725
transform 1 0 235244 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2557
timestamp 1676037725
transform 1 0 236348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_2569
timestamp 1676037725
transform 1 0 237452 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2575
timestamp 1676037725
transform 1 0 238004 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2577
timestamp 1676037725
transform 1 0 238188 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2589
timestamp 1676037725
transform 1 0 239292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2601
timestamp 1676037725
transform 1 0 240396 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2613
timestamp 1676037725
transform 1 0 241500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_2625
timestamp 1676037725
transform 1 0 242604 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2631
timestamp 1676037725
transform 1 0 243156 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2633
timestamp 1676037725
transform 1 0 243340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2645
timestamp 1676037725
transform 1 0 244444 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2657
timestamp 1676037725
transform 1 0 245548 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2669
timestamp 1676037725
transform 1 0 246652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2681
timestamp 1676037725
transform 1 0 247756 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2686
timestamp 1676037725
transform 1 0 248216 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2689
timestamp 1676037725
transform 1 0 248492 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2699
timestamp 1676037725
transform 1 0 249412 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2706
timestamp 1676037725
transform 1 0 250056 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2713
timestamp 1676037725
transform 1 0 250700 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_2725
timestamp 1676037725
transform 1 0 251804 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2733
timestamp 1676037725
transform 1 0 252540 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2740
timestamp 1676037725
transform 1 0 253184 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_2745
timestamp 1676037725
transform 1 0 253644 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_2753
timestamp 1676037725
transform 1 0 254380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2759
timestamp 1676037725
transform 1 0 254932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2769
timestamp 1676037725
transform 1 0 255852 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2779
timestamp 1676037725
transform 1 0 256772 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2786
timestamp 1676037725
transform 1 0 257416 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2798
timestamp 1676037725
transform 1 0 258520 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2801
timestamp 1676037725
transform 1 0 258796 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2818
timestamp 1676037725
transform 1 0 260360 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2827
timestamp 1676037725
transform 1 0 261188 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2840
timestamp 1676037725
transform 1 0 262384 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2844
timestamp 1676037725
transform 1 0 262752 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2854
timestamp 1676037725
transform 1 0 263672 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2857
timestamp 1676037725
transform 1 0 263948 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2868
timestamp 1676037725
transform 1 0 264960 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2881
timestamp 1676037725
transform 1 0 266156 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2894
timestamp 1676037725
transform 1 0 267352 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2907
timestamp 1676037725
transform 1 0 268548 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2911
timestamp 1676037725
transform 1 0 268916 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2913
timestamp 1676037725
transform 1 0 269100 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2924
timestamp 1676037725
transform 1 0 270112 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_2933
timestamp 1676037725
transform 1 0 270940 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1676037725
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1676037725
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1676037725
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1676037725
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1676037725
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1676037725
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1676037725
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1676037725
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 1676037725
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1676037725
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1676037725
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_401
timestamp 1676037725
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_413
timestamp 1676037725
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_419
timestamp 1676037725
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_433
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_445
timestamp 1676037725
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_457
timestamp 1676037725
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_469
timestamp 1676037725
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_475
timestamp 1676037725
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_477
timestamp 1676037725
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_489
timestamp 1676037725
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_501
timestamp 1676037725
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_513
timestamp 1676037725
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_525
timestamp 1676037725
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_531
timestamp 1676037725
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_533
timestamp 1676037725
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_545
timestamp 1676037725
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_557
timestamp 1676037725
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_569
timestamp 1676037725
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_581
timestamp 1676037725
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_587
timestamp 1676037725
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_589
timestamp 1676037725
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_601
timestamp 1676037725
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_613
timestamp 1676037725
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_625
timestamp 1676037725
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_637
timestamp 1676037725
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_643
timestamp 1676037725
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_645
timestamp 1676037725
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_657
timestamp 1676037725
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_669
timestamp 1676037725
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_681
timestamp 1676037725
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_693
timestamp 1676037725
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_699
timestamp 1676037725
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_701
timestamp 1676037725
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_713
timestamp 1676037725
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_725
timestamp 1676037725
transform 1 0 67804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_737
timestamp 1676037725
transform 1 0 68908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_749
timestamp 1676037725
transform 1 0 70012 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_755
timestamp 1676037725
transform 1 0 70564 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_757
timestamp 1676037725
transform 1 0 70748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_769
timestamp 1676037725
transform 1 0 71852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_781
timestamp 1676037725
transform 1 0 72956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_793
timestamp 1676037725
transform 1 0 74060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_805
timestamp 1676037725
transform 1 0 75164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_811
timestamp 1676037725
transform 1 0 75716 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_813
timestamp 1676037725
transform 1 0 75900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_825
timestamp 1676037725
transform 1 0 77004 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_837
timestamp 1676037725
transform 1 0 78108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_849
timestamp 1676037725
transform 1 0 79212 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_861
timestamp 1676037725
transform 1 0 80316 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_867
timestamp 1676037725
transform 1 0 80868 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_869
timestamp 1676037725
transform 1 0 81052 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_881
timestamp 1676037725
transform 1 0 82156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_893
timestamp 1676037725
transform 1 0 83260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_905
timestamp 1676037725
transform 1 0 84364 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_917
timestamp 1676037725
transform 1 0 85468 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_923
timestamp 1676037725
transform 1 0 86020 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_925
timestamp 1676037725
transform 1 0 86204 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_937
timestamp 1676037725
transform 1 0 87308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_949
timestamp 1676037725
transform 1 0 88412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_961
timestamp 1676037725
transform 1 0 89516 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_973
timestamp 1676037725
transform 1 0 90620 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_979
timestamp 1676037725
transform 1 0 91172 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_981
timestamp 1676037725
transform 1 0 91356 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_993
timestamp 1676037725
transform 1 0 92460 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1005
timestamp 1676037725
transform 1 0 93564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1017
timestamp 1676037725
transform 1 0 94668 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_1029
timestamp 1676037725
transform 1 0 95772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_1034
timestamp 1676037725
transform 1 0 96232 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_1037
timestamp 1676037725
transform 1 0 96508 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_1042
timestamp 1676037725
transform 1 0 96968 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1046
timestamp 1676037725
transform 1 0 97336 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_1052
timestamp 1676037725
transform 1 0 97888 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_1061
timestamp 1676037725
transform 1 0 98716 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_1069
timestamp 1676037725
transform 1 0 99452 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_1074
timestamp 1676037725
transform 1 0 99912 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_1082
timestamp 1676037725
transform 1 0 100648 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1086
timestamp 1676037725
transform 1 0 101016 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_1090
timestamp 1676037725
transform 1 0 101384 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_1093
timestamp 1676037725
transform 1 0 101660 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_1098
timestamp 1676037725
transform 1 0 102120 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1105
timestamp 1676037725
transform 1 0 102764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1117
timestamp 1676037725
transform 1 0 103868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1129
timestamp 1676037725
transform 1 0 104972 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1141
timestamp 1676037725
transform 1 0 106076 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_1145
timestamp 1676037725
transform 1 0 106444 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_1149
timestamp 1676037725
transform 1 0 106812 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1153
timestamp 1676037725
transform 1 0 107180 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_1157
timestamp 1676037725
transform 1 0 107548 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_1164
timestamp 1676037725
transform 1 0 108192 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_1173
timestamp 1676037725
transform 1 0 109020 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_1181
timestamp 1676037725
transform 1 0 109756 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1185
timestamp 1676037725
transform 1 0 110124 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_1191
timestamp 1676037725
transform 1 0 110676 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_1198
timestamp 1676037725
transform 1 0 111320 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_1205
timestamp 1676037725
transform 1 0 111964 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_1210
timestamp 1676037725
transform 1 0 112424 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_1217
timestamp 1676037725
transform 1 0 113068 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1223
timestamp 1676037725
transform 1 0 113620 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_1245
timestamp 1676037725
transform 1 0 115644 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_1257
timestamp 1676037725
transform 1 0 116748 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_1261
timestamp 1676037725
transform 1 0 117116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_1269
timestamp 1676037725
transform 1 0 117852 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1277
timestamp 1676037725
transform 1 0 118588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1289
timestamp 1676037725
transform 1 0 119692 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1301
timestamp 1676037725
transform 1 0 120796 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_1313
timestamp 1676037725
transform 1 0 121900 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1317
timestamp 1676037725
transform 1 0 122268 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1329
timestamp 1676037725
transform 1 0 123372 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1341
timestamp 1676037725
transform 1 0 124476 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1353
timestamp 1676037725
transform 1 0 125580 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_1365
timestamp 1676037725
transform 1 0 126684 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1371
timestamp 1676037725
transform 1 0 127236 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1373
timestamp 1676037725
transform 1 0 127420 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1385
timestamp 1676037725
transform 1 0 128524 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1397
timestamp 1676037725
transform 1 0 129628 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1409
timestamp 1676037725
transform 1 0 130732 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_1421
timestamp 1676037725
transform 1 0 131836 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1427
timestamp 1676037725
transform 1 0 132388 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1429
timestamp 1676037725
transform 1 0 132572 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1441
timestamp 1676037725
transform 1 0 133676 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1453
timestamp 1676037725
transform 1 0 134780 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1465
timestamp 1676037725
transform 1 0 135884 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_1477
timestamp 1676037725
transform 1 0 136988 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1483
timestamp 1676037725
transform 1 0 137540 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1485
timestamp 1676037725
transform 1 0 137724 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1497
timestamp 1676037725
transform 1 0 138828 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1509
timestamp 1676037725
transform 1 0 139932 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1521
timestamp 1676037725
transform 1 0 141036 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_1533
timestamp 1676037725
transform 1 0 142140 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1539
timestamp 1676037725
transform 1 0 142692 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1541
timestamp 1676037725
transform 1 0 142876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1553
timestamp 1676037725
transform 1 0 143980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1565
timestamp 1676037725
transform 1 0 145084 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1577
timestamp 1676037725
transform 1 0 146188 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_1589
timestamp 1676037725
transform 1 0 147292 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1595
timestamp 1676037725
transform 1 0 147844 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1597
timestamp 1676037725
transform 1 0 148028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1609
timestamp 1676037725
transform 1 0 149132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_1621
timestamp 1676037725
transform 1 0 150236 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_1636
timestamp 1676037725
transform 1 0 151616 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_1640
timestamp 1676037725
transform 1 0 151984 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_1648
timestamp 1676037725
transform 1 0 152720 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_1653
timestamp 1676037725
transform 1 0 153180 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1658
timestamp 1676037725
transform 1 0 153640 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1670
timestamp 1676037725
transform 1 0 154744 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1682
timestamp 1676037725
transform 1 0 155848 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1694
timestamp 1676037725
transform 1 0 156952 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_1706
timestamp 1676037725
transform 1 0 158056 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1709
timestamp 1676037725
transform 1 0 158332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1721
timestamp 1676037725
transform 1 0 159436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1733
timestamp 1676037725
transform 1 0 160540 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1745
timestamp 1676037725
transform 1 0 161644 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_1757
timestamp 1676037725
transform 1 0 162748 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1763
timestamp 1676037725
transform 1 0 163300 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1765
timestamp 1676037725
transform 1 0 163484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1777
timestamp 1676037725
transform 1 0 164588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1789
timestamp 1676037725
transform 1 0 165692 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1801
timestamp 1676037725
transform 1 0 166796 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_1813
timestamp 1676037725
transform 1 0 167900 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1819
timestamp 1676037725
transform 1 0 168452 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1821
timestamp 1676037725
transform 1 0 168636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1833
timestamp 1676037725
transform 1 0 169740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1845
timestamp 1676037725
transform 1 0 170844 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1857
timestamp 1676037725
transform 1 0 171948 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_1869
timestamp 1676037725
transform 1 0 173052 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1875
timestamp 1676037725
transform 1 0 173604 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1877
timestamp 1676037725
transform 1 0 173788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1889
timestamp 1676037725
transform 1 0 174892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1901
timestamp 1676037725
transform 1 0 175996 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1913
timestamp 1676037725
transform 1 0 177100 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_1925
timestamp 1676037725
transform 1 0 178204 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1931
timestamp 1676037725
transform 1 0 178756 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1933
timestamp 1676037725
transform 1 0 178940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1945
timestamp 1676037725
transform 1 0 180044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1957
timestamp 1676037725
transform 1 0 181148 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1969
timestamp 1676037725
transform 1 0 182252 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_1981
timestamp 1676037725
transform 1 0 183356 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1987
timestamp 1676037725
transform 1 0 183908 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1989
timestamp 1676037725
transform 1 0 184092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2001
timestamp 1676037725
transform 1 0 185196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2013
timestamp 1676037725
transform 1 0 186300 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2025
timestamp 1676037725
transform 1 0 187404 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_2037
timestamp 1676037725
transform 1 0 188508 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_2043
timestamp 1676037725
transform 1 0 189060 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_2045
timestamp 1676037725
transform 1 0 189244 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2053
timestamp 1676037725
transform 1 0 189980 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2058
timestamp 1676037725
transform 1 0 190440 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2070
timestamp 1676037725
transform 1 0 191544 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2082
timestamp 1676037725
transform 1 0 192648 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_2094
timestamp 1676037725
transform 1 0 193752 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2101
timestamp 1676037725
transform 1 0 194396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2113
timestamp 1676037725
transform 1 0 195500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2125
timestamp 1676037725
transform 1 0 196604 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2137
timestamp 1676037725
transform 1 0 197708 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_2149
timestamp 1676037725
transform 1 0 198812 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_2155
timestamp 1676037725
transform 1 0 199364 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2157
timestamp 1676037725
transform 1 0 199548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2169
timestamp 1676037725
transform 1 0 200652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2181
timestamp 1676037725
transform 1 0 201756 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2193
timestamp 1676037725
transform 1 0 202860 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_2205
timestamp 1676037725
transform 1 0 203964 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_2211
timestamp 1676037725
transform 1 0 204516 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2213
timestamp 1676037725
transform 1 0 204700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2225
timestamp 1676037725
transform 1 0 205804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2237
timestamp 1676037725
transform 1 0 206908 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2249
timestamp 1676037725
transform 1 0 208012 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_2261
timestamp 1676037725
transform 1 0 209116 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_2267
timestamp 1676037725
transform 1 0 209668 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2269
timestamp 1676037725
transform 1 0 209852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2281
timestamp 1676037725
transform 1 0 210956 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_2293
timestamp 1676037725
transform 1 0 212060 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2301
timestamp 1676037725
transform 1 0 212796 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_2315
timestamp 1676037725
transform 1 0 214084 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_2323
timestamp 1676037725
transform 1 0 214820 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_2325
timestamp 1676037725
transform 1 0 215004 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2333
timestamp 1676037725
transform 1 0 215740 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2337
timestamp 1676037725
transform 1 0 216108 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_2346
timestamp 1676037725
transform 1 0 216936 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2353
timestamp 1676037725
transform 1 0 217580 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2365
timestamp 1676037725
transform 1 0 218684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_2377
timestamp 1676037725
transform 1 0 219788 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2381
timestamp 1676037725
transform 1 0 220156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2393
timestamp 1676037725
transform 1 0 221260 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_2405
timestamp 1676037725
transform 1 0 222364 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2413
timestamp 1676037725
transform 1 0 223100 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_2419
timestamp 1676037725
transform 1 0 223652 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_2429
timestamp 1676037725
transform 1 0 224572 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_2435
timestamp 1676037725
transform 1 0 225124 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2437
timestamp 1676037725
transform 1 0 225308 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_2445
timestamp 1676037725
transform 1 0 226044 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2460
timestamp 1676037725
transform 1 0 227424 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2472
timestamp 1676037725
transform 1 0 228528 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_2484
timestamp 1676037725
transform 1 0 229632 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2493
timestamp 1676037725
transform 1 0 230460 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2505
timestamp 1676037725
transform 1 0 231564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2517
timestamp 1676037725
transform 1 0 232668 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2529
timestamp 1676037725
transform 1 0 233772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_2541
timestamp 1676037725
transform 1 0 234876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_2547
timestamp 1676037725
transform 1 0 235428 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2549
timestamp 1676037725
transform 1 0 235612 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2561
timestamp 1676037725
transform 1 0 236716 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_2573
timestamp 1676037725
transform 1 0 237820 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2589
timestamp 1676037725
transform 1 0 239292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_2601
timestamp 1676037725
transform 1 0 240396 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2605
timestamp 1676037725
transform 1 0 240764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2617
timestamp 1676037725
transform 1 0 241868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2629
timestamp 1676037725
transform 1 0 242972 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2641
timestamp 1676037725
transform 1 0 244076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_2653
timestamp 1676037725
transform 1 0 245180 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_2659
timestamp 1676037725
transform 1 0 245732 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2661
timestamp 1676037725
transform 1 0 245916 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2673
timestamp 1676037725
transform 1 0 247020 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_2685
timestamp 1676037725
transform 1 0 248124 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_2692
timestamp 1676037725
transform 1 0 248768 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2699
timestamp 1676037725
transform 1 0 249412 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_2711
timestamp 1676037725
transform 1 0 250516 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_2715
timestamp 1676037725
transform 1 0 250884 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2717
timestamp 1676037725
transform 1 0 251068 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2725
timestamp 1676037725
transform 1 0 251804 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_2737
timestamp 1676037725
transform 1 0 252908 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2748
timestamp 1676037725
transform 1 0 253920 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_2760
timestamp 1676037725
transform 1 0 255024 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2770
timestamp 1676037725
transform 1 0 255944 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2773
timestamp 1676037725
transform 1 0 256220 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2778
timestamp 1676037725
transform 1 0 256680 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2790
timestamp 1676037725
transform 1 0 257784 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2802
timestamp 1676037725
transform 1 0 258888 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_2814
timestamp 1676037725
transform 1 0 259992 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2822
timestamp 1676037725
transform 1 0 260728 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2826
timestamp 1676037725
transform 1 0 261096 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_2829
timestamp 1676037725
transform 1 0 261372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2836
timestamp 1676037725
transform 1 0 262016 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2841
timestamp 1676037725
transform 1 0 262476 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2845
timestamp 1676037725
transform 1 0 262844 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2850
timestamp 1676037725
transform 1 0 263304 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_2857
timestamp 1676037725
transform 1 0 263948 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_2870
timestamp 1676037725
transform 1 0 265144 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2882
timestamp 1676037725
transform 1 0 266248 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2885
timestamp 1676037725
transform 1 0 266524 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_2892
timestamp 1676037725
transform 1 0 267168 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_2909
timestamp 1676037725
transform 1 0 268732 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2934
timestamp 1676037725
transform 1 0 271032 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1676037725
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1676037725
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1676037725
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1676037725
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1676037725
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1676037725
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1676037725
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1676037725
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1676037725
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1676037725
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1676037725
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1676037725
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 1676037725
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 1676037725
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 1676037725
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1676037725
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_405
timestamp 1676037725
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_417
timestamp 1676037725
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_429
timestamp 1676037725
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_441
timestamp 1676037725
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_447
timestamp 1676037725
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_461
timestamp 1676037725
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_473
timestamp 1676037725
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_485
timestamp 1676037725
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_497
timestamp 1676037725
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_503
timestamp 1676037725
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_505
timestamp 1676037725
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_517
timestamp 1676037725
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_529
timestamp 1676037725
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_541
timestamp 1676037725
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_553
timestamp 1676037725
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_559
timestamp 1676037725
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_561
timestamp 1676037725
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_573
timestamp 1676037725
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_585
timestamp 1676037725
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_597
timestamp 1676037725
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_609
timestamp 1676037725
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_615
timestamp 1676037725
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_617
timestamp 1676037725
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_629
timestamp 1676037725
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_641
timestamp 1676037725
transform 1 0 60076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_653
timestamp 1676037725
transform 1 0 61180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_665
timestamp 1676037725
transform 1 0 62284 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_671
timestamp 1676037725
transform 1 0 62836 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_673
timestamp 1676037725
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_685
timestamp 1676037725
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_697
timestamp 1676037725
transform 1 0 65228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_709
timestamp 1676037725
transform 1 0 66332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_721
timestamp 1676037725
transform 1 0 67436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_727
timestamp 1676037725
transform 1 0 67988 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_729
timestamp 1676037725
transform 1 0 68172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_741
timestamp 1676037725
transform 1 0 69276 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_753
timestamp 1676037725
transform 1 0 70380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_765
timestamp 1676037725
transform 1 0 71484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_777
timestamp 1676037725
transform 1 0 72588 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_783
timestamp 1676037725
transform 1 0 73140 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_785
timestamp 1676037725
transform 1 0 73324 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_797
timestamp 1676037725
transform 1 0 74428 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_809
timestamp 1676037725
transform 1 0 75532 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_817
timestamp 1676037725
transform 1 0 76268 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_821
timestamp 1676037725
transform 1 0 76636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_833
timestamp 1676037725
transform 1 0 77740 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_839
timestamp 1676037725
transform 1 0 78292 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_841
timestamp 1676037725
transform 1 0 78476 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_847
timestamp 1676037725
transform 1 0 79028 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_859
timestamp 1676037725
transform 1 0 80132 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_871
timestamp 1676037725
transform 1 0 81236 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_883
timestamp 1676037725
transform 1 0 82340 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_895
timestamp 1676037725
transform 1 0 83444 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_897
timestamp 1676037725
transform 1 0 83628 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_909
timestamp 1676037725
transform 1 0 84732 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_921
timestamp 1676037725
transform 1 0 85836 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_933
timestamp 1676037725
transform 1 0 86940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_945
timestamp 1676037725
transform 1 0 88044 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_951
timestamp 1676037725
transform 1 0 88596 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_953
timestamp 1676037725
transform 1 0 88780 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_965
timestamp 1676037725
transform 1 0 89884 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_977
timestamp 1676037725
transform 1 0 90988 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_989
timestamp 1676037725
transform 1 0 92092 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1001
timestamp 1676037725
transform 1 0 93196 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1007
timestamp 1676037725
transform 1 0 93748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_1009
timestamp 1676037725
transform 1 0 93932 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1017
timestamp 1676037725
transform 1 0 94668 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1039
timestamp 1676037725
transform 1 0 96692 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1045
timestamp 1676037725
transform 1 0 97244 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1051
timestamp 1676037725
transform 1 0 97796 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1057
timestamp 1676037725
transform 1 0 98348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_1061
timestamp 1676037725
transform 1 0 98716 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_1065
timestamp 1676037725
transform 1 0 99084 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_1070
timestamp 1676037725
transform 1 0 99544 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1077
timestamp 1676037725
transform 1 0 100188 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1092
timestamp 1676037725
transform 1 0 101568 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1104
timestamp 1676037725
transform 1 0 102672 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_1116
timestamp 1676037725
transform 1 0 103776 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1121
timestamp 1676037725
transform 1 0 104236 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1133
timestamp 1676037725
transform 1 0 105340 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_1145
timestamp 1676037725
transform 1 0 106444 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1149
timestamp 1676037725
transform 1 0 106812 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_1153
timestamp 1676037725
transform 1 0 107180 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_1161
timestamp 1676037725
transform 1 0 107916 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_1167
timestamp 1676037725
transform 1 0 108468 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_1174
timestamp 1676037725
transform 1 0 109112 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_1177
timestamp 1676037725
transform 1 0 109388 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_1182
timestamp 1676037725
transform 1 0 109848 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_1193
timestamp 1676037725
transform 1 0 110860 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_1198
timestamp 1676037725
transform 1 0 111320 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_1202
timestamp 1676037725
transform 1 0 111688 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1225
timestamp 1676037725
transform 1 0 113804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1231
timestamp 1676037725
transform 1 0 114356 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_1233
timestamp 1676037725
transform 1 0 114540 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1237
timestamp 1676037725
transform 1 0 114908 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_1247
timestamp 1676037725
transform 1 0 115828 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1257
timestamp 1676037725
transform 1 0 116748 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_1267
timestamp 1676037725
transform 1 0 117668 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1274
timestamp 1676037725
transform 1 0 118312 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_1286
timestamp 1676037725
transform 1 0 119416 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_1289
timestamp 1676037725
transform 1 0 119692 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1294
timestamp 1676037725
transform 1 0 120152 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1306
timestamp 1676037725
transform 1 0 121256 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1318
timestamp 1676037725
transform 1 0 122360 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1330
timestamp 1676037725
transform 1 0 123464 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_1342
timestamp 1676037725
transform 1 0 124568 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1345
timestamp 1676037725
transform 1 0 124844 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1357
timestamp 1676037725
transform 1 0 125948 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1369
timestamp 1676037725
transform 1 0 127052 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1381
timestamp 1676037725
transform 1 0 128156 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1393
timestamp 1676037725
transform 1 0 129260 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1399
timestamp 1676037725
transform 1 0 129812 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1401
timestamp 1676037725
transform 1 0 129996 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1413
timestamp 1676037725
transform 1 0 131100 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1425
timestamp 1676037725
transform 1 0 132204 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1437
timestamp 1676037725
transform 1 0 133308 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1449
timestamp 1676037725
transform 1 0 134412 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1455
timestamp 1676037725
transform 1 0 134964 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1457
timestamp 1676037725
transform 1 0 135148 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1469
timestamp 1676037725
transform 1 0 136252 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1481
timestamp 1676037725
transform 1 0 137356 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1493
timestamp 1676037725
transform 1 0 138460 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1505
timestamp 1676037725
transform 1 0 139564 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1511
timestamp 1676037725
transform 1 0 140116 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1513
timestamp 1676037725
transform 1 0 140300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1525
timestamp 1676037725
transform 1 0 141404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1537
timestamp 1676037725
transform 1 0 142508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1549
timestamp 1676037725
transform 1 0 143612 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1561
timestamp 1676037725
transform 1 0 144716 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1567
timestamp 1676037725
transform 1 0 145268 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1569
timestamp 1676037725
transform 1 0 145452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1581
timestamp 1676037725
transform 1 0 146556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1593
timestamp 1676037725
transform 1 0 147660 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1605
timestamp 1676037725
transform 1 0 148764 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1617
timestamp 1676037725
transform 1 0 149868 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1623
timestamp 1676037725
transform 1 0 150420 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1625
timestamp 1676037725
transform 1 0 150604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1637
timestamp 1676037725
transform 1 0 151708 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_1644
timestamp 1676037725
transform 1 0 152352 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1652
timestamp 1676037725
transform 1 0 153088 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1664
timestamp 1676037725
transform 1 0 154192 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_1676
timestamp 1676037725
transform 1 0 155296 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1681
timestamp 1676037725
transform 1 0 155756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1693
timestamp 1676037725
transform 1 0 156860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1705
timestamp 1676037725
transform 1 0 157964 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1717
timestamp 1676037725
transform 1 0 159068 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1729
timestamp 1676037725
transform 1 0 160172 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1735
timestamp 1676037725
transform 1 0 160724 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1737
timestamp 1676037725
transform 1 0 160908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_1749
timestamp 1676037725
transform 1 0 162012 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_1755
timestamp 1676037725
transform 1 0 162564 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1763
timestamp 1676037725
transform 1 0 163300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1775
timestamp 1676037725
transform 1 0 164404 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_1787
timestamp 1676037725
transform 1 0 165508 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1791
timestamp 1676037725
transform 1 0 165876 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1793
timestamp 1676037725
transform 1 0 166060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1799
timestamp 1676037725
transform 1 0 166612 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1804
timestamp 1676037725
transform 1 0 167072 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_1816
timestamp 1676037725
transform 1 0 168176 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1823
timestamp 1676037725
transform 1 0 168820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1835
timestamp 1676037725
transform 1 0 169924 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1847
timestamp 1676037725
transform 1 0 171028 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1849
timestamp 1676037725
transform 1 0 171212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1861
timestamp 1676037725
transform 1 0 172316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1873
timestamp 1676037725
transform 1 0 173420 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1885
timestamp 1676037725
transform 1 0 174524 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1897
timestamp 1676037725
transform 1 0 175628 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1903
timestamp 1676037725
transform 1 0 176180 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1905
timestamp 1676037725
transform 1 0 176364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1917
timestamp 1676037725
transform 1 0 177468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1929
timestamp 1676037725
transform 1 0 178572 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1941
timestamp 1676037725
transform 1 0 179676 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1953
timestamp 1676037725
transform 1 0 180780 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1959
timestamp 1676037725
transform 1 0 181332 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1961
timestamp 1676037725
transform 1 0 181516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1973
timestamp 1676037725
transform 1 0 182620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1985
timestamp 1676037725
transform 1 0 183724 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1997
timestamp 1676037725
transform 1 0 184828 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_2009
timestamp 1676037725
transform 1 0 185932 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2015
timestamp 1676037725
transform 1 0 186484 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2017
timestamp 1676037725
transform 1 0 186668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2029
timestamp 1676037725
transform 1 0 187772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2041
timestamp 1676037725
transform 1 0 188876 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2053
timestamp 1676037725
transform 1 0 189980 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_2065
timestamp 1676037725
transform 1 0 191084 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2071
timestamp 1676037725
transform 1 0 191636 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2073
timestamp 1676037725
transform 1 0 191820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2085
timestamp 1676037725
transform 1 0 192924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2097
timestamp 1676037725
transform 1 0 194028 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2109
timestamp 1676037725
transform 1 0 195132 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_2121
timestamp 1676037725
transform 1 0 196236 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2127
timestamp 1676037725
transform 1 0 196788 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2129
timestamp 1676037725
transform 1 0 196972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2141
timestamp 1676037725
transform 1 0 198076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2153
timestamp 1676037725
transform 1 0 199180 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2165
timestamp 1676037725
transform 1 0 200284 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_2177
timestamp 1676037725
transform 1 0 201388 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2183
timestamp 1676037725
transform 1 0 201940 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2185
timestamp 1676037725
transform 1 0 202124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2197
timestamp 1676037725
transform 1 0 203228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2209
timestamp 1676037725
transform 1 0 204332 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2221
timestamp 1676037725
transform 1 0 205436 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_2233
timestamp 1676037725
transform 1 0 206540 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2239
timestamp 1676037725
transform 1 0 207092 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2241
timestamp 1676037725
transform 1 0 207276 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2253
timestamp 1676037725
transform 1 0 208380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2265
timestamp 1676037725
transform 1 0 209484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2277
timestamp 1676037725
transform 1 0 210588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_2289
timestamp 1676037725
transform 1 0 211692 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2295
timestamp 1676037725
transform 1 0 212244 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_2297
timestamp 1676037725
transform 1 0 212428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2305
timestamp 1676037725
transform 1 0 213164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2318
timestamp 1676037725
transform 1 0 214360 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2330
timestamp 1676037725
transform 1 0 215464 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_2342
timestamp 1676037725
transform 1 0 216568 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_2350
timestamp 1676037725
transform 1 0 217304 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_2353
timestamp 1676037725
transform 1 0 217580 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2361
timestamp 1676037725
transform 1 0 218316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2366
timestamp 1676037725
transform 1 0 218776 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2378
timestamp 1676037725
transform 1 0 219880 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2390
timestamp 1676037725
transform 1 0 220984 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2394
timestamp 1676037725
transform 1 0 221352 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_2398
timestamp 1676037725
transform 1 0 221720 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_2406
timestamp 1676037725
transform 1 0 222456 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_2409
timestamp 1676037725
transform 1 0 222732 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_2417
timestamp 1676037725
transform 1 0 223468 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2423
timestamp 1676037725
transform 1 0 224020 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2439
timestamp 1676037725
transform 1 0 225492 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2452
timestamp 1676037725
transform 1 0 226688 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2465
timestamp 1676037725
transform 1 0 227884 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2477
timestamp 1676037725
transform 1 0 228988 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2489
timestamp 1676037725
transform 1 0 230092 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2501
timestamp 1676037725
transform 1 0 231196 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_2513
timestamp 1676037725
transform 1 0 232300 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2519
timestamp 1676037725
transform 1 0 232852 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2521
timestamp 1676037725
transform 1 0 233036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2533
timestamp 1676037725
transform 1 0 234140 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2545
timestamp 1676037725
transform 1 0 235244 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2557
timestamp 1676037725
transform 1 0 236348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_2569
timestamp 1676037725
transform 1 0 237452 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2575
timestamp 1676037725
transform 1 0 238004 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2577
timestamp 1676037725
transform 1 0 238188 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2589
timestamp 1676037725
transform 1 0 239292 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2601
timestamp 1676037725
transform 1 0 240396 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2613
timestamp 1676037725
transform 1 0 241500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_2625
timestamp 1676037725
transform 1 0 242604 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2631
timestamp 1676037725
transform 1 0 243156 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2633
timestamp 1676037725
transform 1 0 243340 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2645
timestamp 1676037725
transform 1 0 244444 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2657
timestamp 1676037725
transform 1 0 245548 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2669
timestamp 1676037725
transform 1 0 246652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_2681
timestamp 1676037725
transform 1 0 247756 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2687
timestamp 1676037725
transform 1 0 248308 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2689
timestamp 1676037725
transform 1 0 248492 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2701
timestamp 1676037725
transform 1 0 249596 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2710
timestamp 1676037725
transform 1 0 250424 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2720
timestamp 1676037725
transform 1 0 251344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2730
timestamp 1676037725
transform 1 0 252264 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2734
timestamp 1676037725
transform 1 0 252632 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2740
timestamp 1676037725
transform 1 0 253184 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2745
timestamp 1676037725
transform 1 0 253644 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2757
timestamp 1676037725
transform 1 0 254748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2769
timestamp 1676037725
transform 1 0 255852 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2781
timestamp 1676037725
transform 1 0 256956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_2793
timestamp 1676037725
transform 1 0 258060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2799
timestamp 1676037725
transform 1 0 258612 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2801
timestamp 1676037725
transform 1 0 258796 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_2813
timestamp 1676037725
transform 1 0 259900 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_2819
timestamp 1676037725
transform 1 0 260452 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_2824
timestamp 1676037725
transform 1 0 260912 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_2828
timestamp 1676037725
transform 1 0 261280 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2833
timestamp 1676037725
transform 1 0 261740 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2840
timestamp 1676037725
transform 1 0 262384 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2847
timestamp 1676037725
transform 1 0 263028 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_2854
timestamp 1676037725
transform 1 0 263672 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_2857
timestamp 1676037725
transform 1 0 263948 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_2863
timestamp 1676037725
transform 1 0 264500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2875
timestamp 1676037725
transform 1 0 265604 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_2883
timestamp 1676037725
transform 1 0 266340 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2896
timestamp 1676037725
transform 1 0 267536 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_2905
timestamp 1676037725
transform 1 0 268364 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2911
timestamp 1676037725
transform 1 0 268916 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2913
timestamp 1676037725
transform 1 0 269100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2917
timestamp 1676037725
transform 1 0 269468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2927
timestamp 1676037725
transform 1 0 270388 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_2934
timestamp 1676037725
transform 1 0 271032 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1676037725
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1676037725
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_221
timestamp 1676037725
transform 1 0 21436 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_228
timestamp 1676037725
transform 1 0 22080 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_234
timestamp 1676037725
transform 1 0 22632 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_239
timestamp 1676037725
transform 1 0 23092 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_247
timestamp 1676037725
transform 1 0 23828 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1676037725
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_259
timestamp 1676037725
transform 1 0 24932 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_264
timestamp 1676037725
transform 1 0 25392 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_276
timestamp 1676037725
transform 1 0 26496 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_288
timestamp 1676037725
transform 1 0 27600 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_300
timestamp 1676037725
transform 1 0 28704 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1676037725
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1676037725
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_348
timestamp 1676037725
transform 1 0 33120 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_360
timestamp 1676037725
transform 1 0 34224 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 1676037725
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_389
timestamp 1676037725
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_401
timestamp 1676037725
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_413
timestamp 1676037725
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_419
timestamp 1676037725
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_433
timestamp 1676037725
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_445
timestamp 1676037725
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_457
timestamp 1676037725
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_469
timestamp 1676037725
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_475
timestamp 1676037725
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_477
timestamp 1676037725
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_489
timestamp 1676037725
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_501
timestamp 1676037725
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_513
timestamp 1676037725
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_525
timestamp 1676037725
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_531
timestamp 1676037725
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_533
timestamp 1676037725
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_545
timestamp 1676037725
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_557
timestamp 1676037725
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_569
timestamp 1676037725
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_581
timestamp 1676037725
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_587
timestamp 1676037725
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_589
timestamp 1676037725
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_601
timestamp 1676037725
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_613
timestamp 1676037725
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_625
timestamp 1676037725
transform 1 0 58604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_637
timestamp 1676037725
transform 1 0 59708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_643
timestamp 1676037725
transform 1 0 60260 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_645
timestamp 1676037725
transform 1 0 60444 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_657
timestamp 1676037725
transform 1 0 61548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_669
timestamp 1676037725
transform 1 0 62652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_681
timestamp 1676037725
transform 1 0 63756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_693
timestamp 1676037725
transform 1 0 64860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_699
timestamp 1676037725
transform 1 0 65412 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_701
timestamp 1676037725
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_713
timestamp 1676037725
transform 1 0 66700 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_720
timestamp 1676037725
transform 1 0 67344 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_727
timestamp 1676037725
transform 1 0 67988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_739
timestamp 1676037725
transform 1 0 69092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_751
timestamp 1676037725
transform 1 0 70196 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_755
timestamp 1676037725
transform 1 0 70564 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_757
timestamp 1676037725
transform 1 0 70748 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_769
timestamp 1676037725
transform 1 0 71852 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_781
timestamp 1676037725
transform 1 0 72956 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_793
timestamp 1676037725
transform 1 0 74060 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_805
timestamp 1676037725
transform 1 0 75164 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_811
timestamp 1676037725
transform 1 0 75716 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_813
timestamp 1676037725
transform 1 0 75900 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_825
timestamp 1676037725
transform 1 0 77004 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_837
timestamp 1676037725
transform 1 0 78108 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_849
timestamp 1676037725
transform 1 0 79212 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_861
timestamp 1676037725
transform 1 0 80316 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_867
timestamp 1676037725
transform 1 0 80868 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_869
timestamp 1676037725
transform 1 0 81052 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_881
timestamp 1676037725
transform 1 0 82156 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_893
timestamp 1676037725
transform 1 0 83260 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_905
timestamp 1676037725
transform 1 0 84364 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_917
timestamp 1676037725
transform 1 0 85468 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_923
timestamp 1676037725
transform 1 0 86020 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_925
timestamp 1676037725
transform 1 0 86204 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_937
timestamp 1676037725
transform 1 0 87308 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_949
timestamp 1676037725
transform 1 0 88412 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_965
timestamp 1676037725
transform 1 0 89884 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_977
timestamp 1676037725
transform 1 0 90988 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_981
timestamp 1676037725
transform 1 0 91356 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_993
timestamp 1676037725
transform 1 0 92460 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1005
timestamp 1676037725
transform 1 0 93564 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1017
timestamp 1676037725
transform 1 0 94668 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1029
timestamp 1676037725
transform 1 0 95772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1035
timestamp 1676037725
transform 1 0 96324 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1037
timestamp 1676037725
transform 1 0 96508 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_1049
timestamp 1676037725
transform 1 0 97612 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1054
timestamp 1676037725
transform 1 0 98072 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1066
timestamp 1676037725
transform 1 0 99176 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_1078
timestamp 1676037725
transform 1 0 100280 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1085
timestamp 1676037725
transform 1 0 100924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1091
timestamp 1676037725
transform 1 0 101476 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1093
timestamp 1676037725
transform 1 0 101660 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1105
timestamp 1676037725
transform 1 0 102764 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1117
timestamp 1676037725
transform 1 0 103868 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1129
timestamp 1676037725
transform 1 0 104972 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1141
timestamp 1676037725
transform 1 0 106076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1147
timestamp 1676037725
transform 1 0 106628 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1149
timestamp 1676037725
transform 1 0 106812 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1161
timestamp 1676037725
transform 1 0 107916 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1173
timestamp 1676037725
transform 1 0 109020 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_1177
timestamp 1676037725
transform 1 0 109388 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1181
timestamp 1676037725
transform 1 0 109756 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1185
timestamp 1676037725
transform 1 0 110124 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1197
timestamp 1676037725
transform 1 0 111228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1203
timestamp 1676037725
transform 1 0 111780 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1205
timestamp 1676037725
transform 1 0 111964 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1217
timestamp 1676037725
transform 1 0 113068 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_1229
timestamp 1676037725
transform 1 0 114172 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_1245
timestamp 1676037725
transform 1 0 115644 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1249
timestamp 1676037725
transform 1 0 116012 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1253
timestamp 1676037725
transform 1 0 116380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1259
timestamp 1676037725
transform 1 0 116932 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1261
timestamp 1676037725
transform 1 0 117116 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1273
timestamp 1676037725
transform 1 0 118220 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1285
timestamp 1676037725
transform 1 0 119324 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1297
timestamp 1676037725
transform 1 0 120428 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1309
timestamp 1676037725
transform 1 0 121532 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1315
timestamp 1676037725
transform 1 0 122084 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1317
timestamp 1676037725
transform 1 0 122268 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1329
timestamp 1676037725
transform 1 0 123372 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1341
timestamp 1676037725
transform 1 0 124476 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1353
timestamp 1676037725
transform 1 0 125580 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1365
timestamp 1676037725
transform 1 0 126684 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1371
timestamp 1676037725
transform 1 0 127236 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1373
timestamp 1676037725
transform 1 0 127420 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1385
timestamp 1676037725
transform 1 0 128524 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1395
timestamp 1676037725
transform 1 0 129444 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1407
timestamp 1676037725
transform 1 0 130548 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_1419
timestamp 1676037725
transform 1 0 131652 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1427
timestamp 1676037725
transform 1 0 132388 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_1429
timestamp 1676037725
transform 1 0 132572 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1435
timestamp 1676037725
transform 1 0 133124 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1450
timestamp 1676037725
transform 1 0 134504 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1462
timestamp 1676037725
transform 1 0 135608 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_1474
timestamp 1676037725
transform 1 0 136712 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_1482
timestamp 1676037725
transform 1 0 137448 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1485
timestamp 1676037725
transform 1 0 137724 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1497
timestamp 1676037725
transform 1 0 138828 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1509
timestamp 1676037725
transform 1 0 139932 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1521
timestamp 1676037725
transform 1 0 141036 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1533
timestamp 1676037725
transform 1 0 142140 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1539
timestamp 1676037725
transform 1 0 142692 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1541
timestamp 1676037725
transform 1 0 142876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1553
timestamp 1676037725
transform 1 0 143980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1565
timestamp 1676037725
transform 1 0 145084 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1577
timestamp 1676037725
transform 1 0 146188 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1589
timestamp 1676037725
transform 1 0 147292 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1595
timestamp 1676037725
transform 1 0 147844 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1597
timestamp 1676037725
transform 1 0 148028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1609
timestamp 1676037725
transform 1 0 149132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1621
timestamp 1676037725
transform 1 0 150236 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1633
timestamp 1676037725
transform 1 0 151340 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1645
timestamp 1676037725
transform 1 0 152444 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1651
timestamp 1676037725
transform 1 0 152996 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1653
timestamp 1676037725
transform 1 0 153180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1665
timestamp 1676037725
transform 1 0 154284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1677
timestamp 1676037725
transform 1 0 155388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1689
timestamp 1676037725
transform 1 0 156492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_1699
timestamp 1676037725
transform 1 0 157412 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1707
timestamp 1676037725
transform 1 0 158148 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_1709
timestamp 1676037725
transform 1 0 158332 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_1715
timestamp 1676037725
transform 1 0 158884 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_1723
timestamp 1676037725
transform 1 0 159620 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_1731
timestamp 1676037725
transform 1 0 160356 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_1739
timestamp 1676037725
transform 1 0 161092 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_1747
timestamp 1676037725
transform 1 0 161828 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_1755
timestamp 1676037725
transform 1 0 162564 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1763
timestamp 1676037725
transform 1 0 163300 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_1765
timestamp 1676037725
transform 1 0 163484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_1771
timestamp 1676037725
transform 1 0 164036 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_1779
timestamp 1676037725
transform 1 0 164772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_1787
timestamp 1676037725
transform 1 0 165508 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_1795
timestamp 1676037725
transform 1 0 166244 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_1803
timestamp 1676037725
transform 1 0 166980 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1811
timestamp 1676037725
transform 1 0 167716 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_1817
timestamp 1676037725
transform 1 0 168268 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_1821
timestamp 1676037725
transform 1 0 168636 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1828
timestamp 1676037725
transform 1 0 169280 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1840
timestamp 1676037725
transform 1 0 170384 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1852
timestamp 1676037725
transform 1 0 171488 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1864
timestamp 1676037725
transform 1 0 172592 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1877
timestamp 1676037725
transform 1 0 173788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1889
timestamp 1676037725
transform 1 0 174892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1901
timestamp 1676037725
transform 1 0 175996 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1913
timestamp 1676037725
transform 1 0 177100 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1925
timestamp 1676037725
transform 1 0 178204 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1931
timestamp 1676037725
transform 1 0 178756 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1933
timestamp 1676037725
transform 1 0 178940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1945
timestamp 1676037725
transform 1 0 180044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1957
timestamp 1676037725
transform 1 0 181148 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1969
timestamp 1676037725
transform 1 0 182252 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1981
timestamp 1676037725
transform 1 0 183356 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1987
timestamp 1676037725
transform 1 0 183908 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1989
timestamp 1676037725
transform 1 0 184092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2001
timestamp 1676037725
transform 1 0 185196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2013
timestamp 1676037725
transform 1 0 186300 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2025
timestamp 1676037725
transform 1 0 187404 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_2037
timestamp 1676037725
transform 1 0 188508 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2043
timestamp 1676037725
transform 1 0 189060 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2045
timestamp 1676037725
transform 1 0 189244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2057
timestamp 1676037725
transform 1 0 190348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2069
timestamp 1676037725
transform 1 0 191452 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2081
timestamp 1676037725
transform 1 0 192556 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_2093
timestamp 1676037725
transform 1 0 193660 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2099
timestamp 1676037725
transform 1 0 194212 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2101
timestamp 1676037725
transform 1 0 194396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2113
timestamp 1676037725
transform 1 0 195500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2125
timestamp 1676037725
transform 1 0 196604 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2137
timestamp 1676037725
transform 1 0 197708 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_2149
timestamp 1676037725
transform 1 0 198812 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2155
timestamp 1676037725
transform 1 0 199364 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2157
timestamp 1676037725
transform 1 0 199548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2169
timestamp 1676037725
transform 1 0 200652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2181
timestamp 1676037725
transform 1 0 201756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2193
timestamp 1676037725
transform 1 0 202860 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2197
timestamp 1676037725
transform 1 0 203228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_2209
timestamp 1676037725
transform 1 0 204332 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2213
timestamp 1676037725
transform 1 0 204700 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2225
timestamp 1676037725
transform 1 0 205804 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2237
timestamp 1676037725
transform 1 0 206908 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2249
timestamp 1676037725
transform 1 0 208012 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_2261
timestamp 1676037725
transform 1 0 209116 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2267
timestamp 1676037725
transform 1 0 209668 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2269
timestamp 1676037725
transform 1 0 209852 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2281
timestamp 1676037725
transform 1 0 210956 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2293
timestamp 1676037725
transform 1 0 212060 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2305
timestamp 1676037725
transform 1 0 213164 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_2317
timestamp 1676037725
transform 1 0 214268 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2323
timestamp 1676037725
transform 1 0 214820 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2325
timestamp 1676037725
transform 1 0 215004 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2337
timestamp 1676037725
transform 1 0 216108 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2349
timestamp 1676037725
transform 1 0 217212 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2361
timestamp 1676037725
transform 1 0 218316 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_2373
timestamp 1676037725
transform 1 0 219420 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2379
timestamp 1676037725
transform 1 0 219972 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2381
timestamp 1676037725
transform 1 0 220156 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2393
timestamp 1676037725
transform 1 0 221260 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2405
timestamp 1676037725
transform 1 0 222364 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_2417
timestamp 1676037725
transform 1 0 223468 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2425
timestamp 1676037725
transform 1 0 224204 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2432
timestamp 1676037725
transform 1 0 224848 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_2437
timestamp 1676037725
transform 1 0 225308 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2443
timestamp 1676037725
transform 1 0 225860 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2455
timestamp 1676037725
transform 1 0 226964 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2467
timestamp 1676037725
transform 1 0 228068 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2479
timestamp 1676037725
transform 1 0 229172 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2491
timestamp 1676037725
transform 1 0 230276 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2493
timestamp 1676037725
transform 1 0 230460 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2505
timestamp 1676037725
transform 1 0 231564 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2517
timestamp 1676037725
transform 1 0 232668 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_2529
timestamp 1676037725
transform 1 0 233772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_2537
timestamp 1676037725
transform 1 0 234508 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2543
timestamp 1676037725
transform 1 0 235060 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2547
timestamp 1676037725
transform 1 0 235428 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_2549
timestamp 1676037725
transform 1 0 235612 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2554
timestamp 1676037725
transform 1 0 236072 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2566
timestamp 1676037725
transform 1 0 237176 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2578
timestamp 1676037725
transform 1 0 238280 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2590
timestamp 1676037725
transform 1 0 239384 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_2602
timestamp 1676037725
transform 1 0 240488 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2605
timestamp 1676037725
transform 1 0 240764 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2617
timestamp 1676037725
transform 1 0 241868 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2629
timestamp 1676037725
transform 1 0 242972 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2641
timestamp 1676037725
transform 1 0 244076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_2653
timestamp 1676037725
transform 1 0 245180 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2659
timestamp 1676037725
transform 1 0 245732 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2661
timestamp 1676037725
transform 1 0 245916 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2673
timestamp 1676037725
transform 1 0 247020 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2685
timestamp 1676037725
transform 1 0 248124 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2697
timestamp 1676037725
transform 1 0 249228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_2709
timestamp 1676037725
transform 1 0 250332 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2715
timestamp 1676037725
transform 1 0 250884 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2717
timestamp 1676037725
transform 1 0 251068 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2729
timestamp 1676037725
transform 1 0 252172 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2741
timestamp 1676037725
transform 1 0 253276 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2753
timestamp 1676037725
transform 1 0 254380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_2765
timestamp 1676037725
transform 1 0 255484 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2771
timestamp 1676037725
transform 1 0 256036 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2773
timestamp 1676037725
transform 1 0 256220 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2785
timestamp 1676037725
transform 1 0 257324 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_2797
timestamp 1676037725
transform 1 0 258428 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_2805
timestamp 1676037725
transform 1 0 259164 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_2810
timestamp 1676037725
transform 1 0 259624 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_2814
timestamp 1676037725
transform 1 0 259992 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2819
timestamp 1676037725
transform 1 0 260452 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_2826
timestamp 1676037725
transform 1 0 261096 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_2829
timestamp 1676037725
transform 1 0 261372 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2835
timestamp 1676037725
transform 1 0 261924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2843
timestamp 1676037725
transform 1 0 262660 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2847
timestamp 1676037725
transform 1 0 263028 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2852
timestamp 1676037725
transform 1 0 263488 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2856
timestamp 1676037725
transform 1 0 263856 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2862
timestamp 1676037725
transform 1 0 264408 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2870
timestamp 1676037725
transform 1 0 265144 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2879
timestamp 1676037725
transform 1 0 265972 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2883
timestamp 1676037725
transform 1 0 266340 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_2885
timestamp 1676037725
transform 1 0 266524 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2896
timestamp 1676037725
transform 1 0 267536 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2905
timestamp 1676037725
transform 1 0 268364 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2915
timestamp 1676037725
transform 1 0 269284 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2927
timestamp 1676037725
transform 1 0 270388 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_2934
timestamp 1676037725
transform 1 0 271032 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 1676037725
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_217
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_222
timestamp 1676037725
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_232
timestamp 1676037725
transform 1 0 22448 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_239
timestamp 1676037725
transform 1 0 23092 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_243
timestamp 1676037725
transform 1 0 23460 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_250
timestamp 1676037725
transform 1 0 24104 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_254
timestamp 1676037725
transform 1 0 24472 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_261
timestamp 1676037725
transform 1 0 25116 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_267
timestamp 1676037725
transform 1 0 25668 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_270
timestamp 1676037725
transform 1 0 25944 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_277
timestamp 1676037725
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_288
timestamp 1676037725
transform 1 0 27600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_296
timestamp 1676037725
transform 1 0 28336 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_304
timestamp 1676037725
transform 1 0 29072 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_313
timestamp 1676037725
transform 1 0 29900 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_321
timestamp 1676037725
transform 1 0 30636 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_327
timestamp 1676037725
transform 1 0 31188 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 1676037725
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_343
timestamp 1676037725
transform 1 0 32660 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_349
timestamp 1676037725
transform 1 0 33212 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_357
timestamp 1676037725
transform 1 0 33948 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_369
timestamp 1676037725
transform 1 0 35052 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_381
timestamp 1676037725
transform 1 0 36156 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_389
timestamp 1676037725
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_405
timestamp 1676037725
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_417
timestamp 1676037725
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_429
timestamp 1676037725
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_441
timestamp 1676037725
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_447
timestamp 1676037725
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_461
timestamp 1676037725
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_473
timestamp 1676037725
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_485
timestamp 1676037725
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_497
timestamp 1676037725
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_503
timestamp 1676037725
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_505
timestamp 1676037725
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_517
timestamp 1676037725
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_529
timestamp 1676037725
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_541
timestamp 1676037725
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_553
timestamp 1676037725
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_559
timestamp 1676037725
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_561
timestamp 1676037725
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_573
timestamp 1676037725
transform 1 0 53820 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_579
timestamp 1676037725
transform 1 0 54372 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_585
timestamp 1676037725
transform 1 0 54924 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_596
timestamp 1676037725
transform 1 0 55936 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_602
timestamp 1676037725
transform 1 0 56488 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_605
timestamp 1676037725
transform 1 0 56764 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_612
timestamp 1676037725
transform 1 0 57408 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_617
timestamp 1676037725
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_629
timestamp 1676037725
transform 1 0 58972 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_637
timestamp 1676037725
transform 1 0 59708 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_645
timestamp 1676037725
transform 1 0 60444 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_653
timestamp 1676037725
transform 1 0 61180 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_657
timestamp 1676037725
transform 1 0 61548 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_660
timestamp 1676037725
transform 1 0 61824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_669
timestamp 1676037725
transform 1 0 62652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_673
timestamp 1676037725
transform 1 0 63020 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_685
timestamp 1676037725
transform 1 0 64124 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_693
timestamp 1676037725
transform 1 0 64860 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_697
timestamp 1676037725
transform 1 0 65228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_702
timestamp 1676037725
transform 1 0 65688 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_710
timestamp 1676037725
transform 1 0 66424 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_726
timestamp 1676037725
transform 1 0 67896 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_729
timestamp 1676037725
transform 1 0 68172 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_741
timestamp 1676037725
transform 1 0 69276 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_753
timestamp 1676037725
transform 1 0 70380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_765
timestamp 1676037725
transform 1 0 71484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_777
timestamp 1676037725
transform 1 0 72588 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_783
timestamp 1676037725
transform 1 0 73140 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_785
timestamp 1676037725
transform 1 0 73324 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_793
timestamp 1676037725
transform 1 0 74060 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_805
timestamp 1676037725
transform 1 0 75164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_817
timestamp 1676037725
transform 1 0 76268 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_829
timestamp 1676037725
transform 1 0 77372 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_837
timestamp 1676037725
transform 1 0 78108 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_841
timestamp 1676037725
transform 1 0 78476 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_853
timestamp 1676037725
transform 1 0 79580 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_865
timestamp 1676037725
transform 1 0 80684 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_877
timestamp 1676037725
transform 1 0 81788 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_889
timestamp 1676037725
transform 1 0 82892 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_895
timestamp 1676037725
transform 1 0 83444 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_897
timestamp 1676037725
transform 1 0 83628 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_909
timestamp 1676037725
transform 1 0 84732 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_921
timestamp 1676037725
transform 1 0 85836 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_933
timestamp 1676037725
transform 1 0 86940 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_945
timestamp 1676037725
transform 1 0 88044 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_951
timestamp 1676037725
transform 1 0 88596 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_957
timestamp 1676037725
transform 1 0 89148 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_961
timestamp 1676037725
transform 1 0 89516 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_968
timestamp 1676037725
transform 1 0 90160 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_972
timestamp 1676037725
transform 1 0 90528 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_977
timestamp 1676037725
transform 1 0 90988 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_981
timestamp 1676037725
transform 1 0 91356 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_988
timestamp 1676037725
transform 1 0 92000 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_996
timestamp 1676037725
transform 1 0 92736 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1004
timestamp 1676037725
transform 1 0 93472 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1009
timestamp 1676037725
transform 1 0 93932 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1013
timestamp 1676037725
transform 1 0 94300 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1018
timestamp 1676037725
transform 1 0 94760 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1023
timestamp 1676037725
transform 1 0 95220 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1027
timestamp 1676037725
transform 1 0 95588 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_1034
timestamp 1676037725
transform 1 0 96232 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1042
timestamp 1676037725
transform 1 0 96968 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1050
timestamp 1676037725
transform 1 0 97704 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1058
timestamp 1676037725
transform 1 0 98440 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1065
timestamp 1676037725
transform 1 0 99084 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1075
timestamp 1676037725
transform 1 0 100004 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1081
timestamp 1676037725
transform 1 0 100556 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1092
timestamp 1676037725
transform 1 0 101568 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1099
timestamp 1676037725
transform 1 0 102212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_1111
timestamp 1676037725
transform 1 0 103316 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1119
timestamp 1676037725
transform 1 0 104052 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1121
timestamp 1676037725
transform 1 0 104236 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1133
timestamp 1676037725
transform 1 0 105340 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1145
timestamp 1676037725
transform 1 0 106444 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1157
timestamp 1676037725
transform 1 0 107548 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1169
timestamp 1676037725
transform 1 0 108652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1175
timestamp 1676037725
transform 1 0 109204 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1177
timestamp 1676037725
transform 1 0 109388 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1189
timestamp 1676037725
transform 1 0 110492 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1201
timestamp 1676037725
transform 1 0 111596 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1213
timestamp 1676037725
transform 1 0 112700 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1225
timestamp 1676037725
transform 1 0 113804 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1231
timestamp 1676037725
transform 1 0 114356 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1233
timestamp 1676037725
transform 1 0 114540 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1245
timestamp 1676037725
transform 1 0 115644 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1257
timestamp 1676037725
transform 1 0 116748 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1269
timestamp 1676037725
transform 1 0 117852 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1281
timestamp 1676037725
transform 1 0 118956 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1287
timestamp 1676037725
transform 1 0 119508 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1289
timestamp 1676037725
transform 1 0 119692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1301
timestamp 1676037725
transform 1 0 120796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1305
timestamp 1676037725
transform 1 0 121164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1311
timestamp 1676037725
transform 1 0 121716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1315
timestamp 1676037725
transform 1 0 122084 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1320
timestamp 1676037725
transform 1 0 122544 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1324
timestamp 1676037725
transform 1 0 122912 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1329
timestamp 1676037725
transform 1 0 123372 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1333
timestamp 1676037725
transform 1 0 123740 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1338
timestamp 1676037725
transform 1 0 124200 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1345
timestamp 1676037725
transform 1 0 124844 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_1355
timestamp 1676037725
transform 1 0 125764 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_1363
timestamp 1676037725
transform 1 0 126500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1370
timestamp 1676037725
transform 1 0 127144 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1378
timestamp 1676037725
transform 1 0 127880 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1384
timestamp 1676037725
transform 1 0 128432 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1388
timestamp 1676037725
transform 1 0 128800 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1395
timestamp 1676037725
transform 1 0 129444 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1399
timestamp 1676037725
transform 1 0 129812 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1401
timestamp 1676037725
transform 1 0 129996 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1408
timestamp 1676037725
transform 1 0 130640 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_1412
timestamp 1676037725
transform 1 0 131008 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1420
timestamp 1676037725
transform 1 0 131744 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1426
timestamp 1676037725
transform 1 0 132296 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_1435
timestamp 1676037725
transform 1 0 133124 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_1443
timestamp 1676037725
transform 1 0 133860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1451
timestamp 1676037725
transform 1 0 134596 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1455
timestamp 1676037725
transform 1 0 134964 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1457
timestamp 1676037725
transform 1 0 135148 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1469
timestamp 1676037725
transform 1 0 136252 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1481
timestamp 1676037725
transform 1 0 137356 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1493
timestamp 1676037725
transform 1 0 138460 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1505
timestamp 1676037725
transform 1 0 139564 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1511
timestamp 1676037725
transform 1 0 140116 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1513
timestamp 1676037725
transform 1 0 140300 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1525
timestamp 1676037725
transform 1 0 141404 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1537
timestamp 1676037725
transform 1 0 142508 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1549
timestamp 1676037725
transform 1 0 143612 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1561
timestamp 1676037725
transform 1 0 144716 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1567
timestamp 1676037725
transform 1 0 145268 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1569
timestamp 1676037725
transform 1 0 145452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1581
timestamp 1676037725
transform 1 0 146556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1593
timestamp 1676037725
transform 1 0 147660 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1605
timestamp 1676037725
transform 1 0 148764 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1617
timestamp 1676037725
transform 1 0 149868 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1623
timestamp 1676037725
transform 1 0 150420 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1625
timestamp 1676037725
transform 1 0 150604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1637
timestamp 1676037725
transform 1 0 151708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1649
timestamp 1676037725
transform 1 0 152812 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1661
timestamp 1676037725
transform 1 0 153916 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1673
timestamp 1676037725
transform 1 0 155020 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1679
timestamp 1676037725
transform 1 0 155572 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1681
timestamp 1676037725
transform 1 0 155756 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1687
timestamp 1676037725
transform 1 0 156308 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1696
timestamp 1676037725
transform 1 0 157136 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1702
timestamp 1676037725
transform 1 0 157688 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1708
timestamp 1676037725
transform 1 0 158240 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1712
timestamp 1676037725
transform 1 0 158608 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1723
timestamp 1676037725
transform 1 0 159620 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1732
timestamp 1676037725
transform 1 0 160448 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1737
timestamp 1676037725
transform 1 0 160908 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1743
timestamp 1676037725
transform 1 0 161460 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1747
timestamp 1676037725
transform 1 0 161828 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1758
timestamp 1676037725
transform 1 0 162840 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1764
timestamp 1676037725
transform 1 0 163392 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1775
timestamp 1676037725
transform 1 0 164404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1779
timestamp 1676037725
transform 1 0 164772 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1790
timestamp 1676037725
transform 1 0 165784 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1793
timestamp 1676037725
transform 1 0 166060 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1800
timestamp 1676037725
transform 1 0 166704 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1804
timestamp 1676037725
transform 1 0 167072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1815
timestamp 1676037725
transform 1 0 168084 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1831
timestamp 1676037725
transform 1 0 169556 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_1838
timestamp 1676037725
transform 1 0 170200 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1846
timestamp 1676037725
transform 1 0 170936 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1849
timestamp 1676037725
transform 1 0 171212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1861
timestamp 1676037725
transform 1 0 172316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1873
timestamp 1676037725
transform 1 0 173420 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1885
timestamp 1676037725
transform 1 0 174524 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1897
timestamp 1676037725
transform 1 0 175628 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1903
timestamp 1676037725
transform 1 0 176180 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1905
timestamp 1676037725
transform 1 0 176364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1917
timestamp 1676037725
transform 1 0 177468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1929
timestamp 1676037725
transform 1 0 178572 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1941
timestamp 1676037725
transform 1 0 179676 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1953
timestamp 1676037725
transform 1 0 180780 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1959
timestamp 1676037725
transform 1 0 181332 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1961
timestamp 1676037725
transform 1 0 181516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1973
timestamp 1676037725
transform 1 0 182620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1985
timestamp 1676037725
transform 1 0 183724 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1997
timestamp 1676037725
transform 1 0 184828 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_2009
timestamp 1676037725
transform 1 0 185932 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2015
timestamp 1676037725
transform 1 0 186484 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_2017
timestamp 1676037725
transform 1 0 186668 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2030
timestamp 1676037725
transform 1 0 187864 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2042
timestamp 1676037725
transform 1 0 188968 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_2054
timestamp 1676037725
transform 1 0 190072 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2061
timestamp 1676037725
transform 1 0 190716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_2069
timestamp 1676037725
transform 1 0 191452 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2073
timestamp 1676037725
transform 1 0 191820 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2077
timestamp 1676037725
transform 1 0 192188 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2083
timestamp 1676037725
transform 1 0 192740 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2091
timestamp 1676037725
transform 1 0 193476 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_2099
timestamp 1676037725
transform 1 0 194212 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_2107
timestamp 1676037725
transform 1 0 194948 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2115
timestamp 1676037725
transform 1 0 195684 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2123
timestamp 1676037725
transform 1 0 196420 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2127
timestamp 1676037725
transform 1 0 196788 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2129
timestamp 1676037725
transform 1 0 196972 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_2136
timestamp 1676037725
transform 1 0 197616 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2147
timestamp 1676037725
transform 1 0 198628 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2155
timestamp 1676037725
transform 1 0 199364 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2163
timestamp 1676037725
transform 1 0 200100 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2167
timestamp 1676037725
transform 1 0 200468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2172
timestamp 1676037725
transform 1 0 200928 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2180
timestamp 1676037725
transform 1 0 201664 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2185
timestamp 1676037725
transform 1 0 202124 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2192
timestamp 1676037725
transform 1 0 202768 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2201
timestamp 1676037725
transform 1 0 203596 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2213
timestamp 1676037725
transform 1 0 204700 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2225
timestamp 1676037725
transform 1 0 205804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_2237
timestamp 1676037725
transform 1 0 206908 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2241
timestamp 1676037725
transform 1 0 207276 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2253
timestamp 1676037725
transform 1 0 208380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2265
timestamp 1676037725
transform 1 0 209484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2277
timestamp 1676037725
transform 1 0 210588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_2289
timestamp 1676037725
transform 1 0 211692 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2295
timestamp 1676037725
transform 1 0 212244 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2297
timestamp 1676037725
transform 1 0 212428 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2309
timestamp 1676037725
transform 1 0 213532 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2321
timestamp 1676037725
transform 1 0 214636 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2333
timestamp 1676037725
transform 1 0 215740 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_2345
timestamp 1676037725
transform 1 0 216844 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2351
timestamp 1676037725
transform 1 0 217396 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2353
timestamp 1676037725
transform 1 0 217580 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2365
timestamp 1676037725
transform 1 0 218684 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2377
timestamp 1676037725
transform 1 0 219788 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2389
timestamp 1676037725
transform 1 0 220892 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_2401
timestamp 1676037725
transform 1 0 221996 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2407
timestamp 1676037725
transform 1 0 222548 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_2409
timestamp 1676037725
transform 1 0 222732 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2417
timestamp 1676037725
transform 1 0 223468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_2422
timestamp 1676037725
transform 1 0 223928 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2432
timestamp 1676037725
transform 1 0 224848 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2436
timestamp 1676037725
transform 1 0 225216 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2441
timestamp 1676037725
transform 1 0 225676 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2449
timestamp 1676037725
transform 1 0 226412 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_2457
timestamp 1676037725
transform 1 0 227148 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2463
timestamp 1676037725
transform 1 0 227700 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2465
timestamp 1676037725
transform 1 0 227884 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2472
timestamp 1676037725
transform 1 0 228528 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2476
timestamp 1676037725
transform 1 0 228896 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_2481
timestamp 1676037725
transform 1 0 229356 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2492
timestamp 1676037725
transform 1 0 230368 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2500
timestamp 1676037725
transform 1 0 231104 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_2508
timestamp 1676037725
transform 1 0 231840 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2518
timestamp 1676037725
transform 1 0 232760 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2521
timestamp 1676037725
transform 1 0 233036 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2530
timestamp 1676037725
transform 1 0 233864 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2538
timestamp 1676037725
transform 1 0 234600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2542
timestamp 1676037725
transform 1 0 234968 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_2548
timestamp 1676037725
transform 1 0 235520 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2558
timestamp 1676037725
transform 1 0 236440 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_2570
timestamp 1676037725
transform 1 0 237544 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2577
timestamp 1676037725
transform 1 0 238188 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2589
timestamp 1676037725
transform 1 0 239292 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2601
timestamp 1676037725
transform 1 0 240396 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2613
timestamp 1676037725
transform 1 0 241500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_2625
timestamp 1676037725
transform 1 0 242604 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2631
timestamp 1676037725
transform 1 0 243156 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2633
timestamp 1676037725
transform 1 0 243340 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2645
timestamp 1676037725
transform 1 0 244444 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2657
timestamp 1676037725
transform 1 0 245548 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2669
timestamp 1676037725
transform 1 0 246652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_2681
timestamp 1676037725
transform 1 0 247756 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2687
timestamp 1676037725
transform 1 0 248308 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2689
timestamp 1676037725
transform 1 0 248492 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2701
timestamp 1676037725
transform 1 0 249596 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2713
timestamp 1676037725
transform 1 0 250700 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2725
timestamp 1676037725
transform 1 0 251804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_2737
timestamp 1676037725
transform 1 0 252908 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2743
timestamp 1676037725
transform 1 0 253460 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2745
timestamp 1676037725
transform 1 0 253644 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2757
timestamp 1676037725
transform 1 0 254748 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_2769
timestamp 1676037725
transform 1 0 255852 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2777
timestamp 1676037725
transform 1 0 256588 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2788
timestamp 1676037725
transform 1 0 257600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2792
timestamp 1676037725
transform 1 0 257968 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_2797
timestamp 1676037725
transform 1 0 258428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2801
timestamp 1676037725
transform 1 0 258796 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2807
timestamp 1676037725
transform 1 0 259348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2815
timestamp 1676037725
transform 1 0 260084 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2821
timestamp 1676037725
transform 1 0 260636 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2825
timestamp 1676037725
transform 1 0 261004 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2833
timestamp 1676037725
transform 1 0 261740 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2841
timestamp 1676037725
transform 1 0 262476 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2851
timestamp 1676037725
transform 1 0 263396 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2855
timestamp 1676037725
transform 1 0 263764 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2857
timestamp 1676037725
transform 1 0 263948 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2865
timestamp 1676037725
transform 1 0 264684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2869
timestamp 1676037725
transform 1 0 265052 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2873
timestamp 1676037725
transform 1 0 265420 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2881
timestamp 1676037725
transform 1 0 266156 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2890
timestamp 1676037725
transform 1 0 266984 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2894
timestamp 1676037725
transform 1 0 267352 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2900
timestamp 1676037725
transform 1 0 267904 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2910
timestamp 1676037725
transform 1 0 268824 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_2913
timestamp 1676037725
transform 1 0 269100 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2923
timestamp 1676037725
transform 1 0 270020 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2932
timestamp 1676037725
transform 1 0 270848 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_8
timestamp 1676037725
transform 1 0 1840 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_20
timestamp 1676037725
transform 1 0 2944 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_25
timestamp 1676037725
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_81
timestamp 1676037725
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_137
timestamp 1676037725
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 1676037725
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 1676037725
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1676037725
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_205
timestamp 1676037725
transform 1 0 19964 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_212
timestamp 1676037725
transform 1 0 20608 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_225
timestamp 1676037725
transform 1 0 21804 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_232
timestamp 1676037725
transform 1 0 22448 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_242
timestamp 1676037725
transform 1 0 23368 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_250
timestamp 1676037725
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_261
timestamp 1676037725
transform 1 0 25116 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_275
timestamp 1676037725
transform 1 0 26404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_279
timestamp 1676037725
transform 1 0 26772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_286
timestamp 1676037725
transform 1 0 27416 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_295
timestamp 1676037725
transform 1 0 28244 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_304
timestamp 1676037725
transform 1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_313
timestamp 1676037725
transform 1 0 29900 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_319
timestamp 1676037725
transform 1 0 30452 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_327
timestamp 1676037725
transform 1 0 31188 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_331
timestamp 1676037725
transform 1 0 31556 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_338
timestamp 1676037725
transform 1 0 32200 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_344
timestamp 1676037725
transform 1 0 32752 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_349
timestamp 1676037725
transform 1 0 33212 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_361
timestamp 1676037725
transform 1 0 34316 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_371
timestamp 1676037725
transform 1 0 35236 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_383
timestamp 1676037725
transform 1 0 36340 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_395
timestamp 1676037725
transform 1 0 37444 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_407
timestamp 1676037725
transform 1 0 38548 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_419
timestamp 1676037725
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_421
timestamp 1676037725
transform 1 0 39836 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_427
timestamp 1676037725
transform 1 0 40388 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_439
timestamp 1676037725
transform 1 0 41492 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_451
timestamp 1676037725
transform 1 0 42596 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_463
timestamp 1676037725
transform 1 0 43700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_475
timestamp 1676037725
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_477
timestamp 1676037725
transform 1 0 44988 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_483
timestamp 1676037725
transform 1 0 45540 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_495
timestamp 1676037725
transform 1 0 46644 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_507
timestamp 1676037725
transform 1 0 47748 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_519
timestamp 1676037725
transform 1 0 48852 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_531
timestamp 1676037725
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_533
timestamp 1676037725
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_545
timestamp 1676037725
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_557
timestamp 1676037725
transform 1 0 52348 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_569
timestamp 1676037725
transform 1 0 53452 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_575
timestamp 1676037725
transform 1 0 54004 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_579
timestamp 1676037725
transform 1 0 54372 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_586
timestamp 1676037725
transform 1 0 55016 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_589
timestamp 1676037725
transform 1 0 55292 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_595
timestamp 1676037725
transform 1 0 55844 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_604
timestamp 1676037725
transform 1 0 56672 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_611
timestamp 1676037725
transform 1 0 57316 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_615
timestamp 1676037725
transform 1 0 57684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_622
timestamp 1676037725
transform 1 0 58328 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_626
timestamp 1676037725
transform 1 0 58696 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_633
timestamp 1676037725
transform 1 0 59340 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_642
timestamp 1676037725
transform 1 0 60168 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_645
timestamp 1676037725
transform 1 0 60444 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_652
timestamp 1676037725
transform 1 0 61088 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_658
timestamp 1676037725
transform 1 0 61640 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_665
timestamp 1676037725
transform 1 0 62284 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_671
timestamp 1676037725
transform 1 0 62836 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_680
timestamp 1676037725
transform 1 0 63664 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_689
timestamp 1676037725
transform 1 0 64492 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_698
timestamp 1676037725
transform 1 0 65320 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_701
timestamp 1676037725
transform 1 0 65596 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_705
timestamp 1676037725
transform 1 0 65964 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_711
timestamp 1676037725
transform 1 0 66516 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_715
timestamp 1676037725
transform 1 0 66884 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_720
timestamp 1676037725
transform 1 0 67344 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_732
timestamp 1676037725
transform 1 0 68448 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_744
timestamp 1676037725
transform 1 0 69552 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_750
timestamp 1676037725
transform 1 0 70104 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_757
timestamp 1676037725
transform 1 0 70748 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_769
timestamp 1676037725
transform 1 0 71852 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_781
timestamp 1676037725
transform 1 0 72956 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_785
timestamp 1676037725
transform 1 0 73324 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_796
timestamp 1676037725
transform 1 0 74336 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_810
timestamp 1676037725
transform 1 0 75624 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_813
timestamp 1676037725
transform 1 0 75900 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_825
timestamp 1676037725
transform 1 0 77004 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_837
timestamp 1676037725
transform 1 0 78108 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_853
timestamp 1676037725
transform 1 0 79580 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_865
timestamp 1676037725
transform 1 0 80684 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_869
timestamp 1676037725
transform 1 0 81052 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_881
timestamp 1676037725
transform 1 0 82156 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_889
timestamp 1676037725
transform 1 0 82892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_901
timestamp 1676037725
transform 1 0 83996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_913
timestamp 1676037725
transform 1 0 85100 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_921
timestamp 1676037725
transform 1 0 85836 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_925
timestamp 1676037725
transform 1 0 86204 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_937
timestamp 1676037725
transform 1 0 87308 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_945
timestamp 1676037725
transform 1 0 88044 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_951
timestamp 1676037725
transform 1 0 88596 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_960
timestamp 1676037725
transform 1 0 89424 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_969
timestamp 1676037725
transform 1 0 90252 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_978
timestamp 1676037725
transform 1 0 91080 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_981
timestamp 1676037725
transform 1 0 91356 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_987
timestamp 1676037725
transform 1 0 91908 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_996
timestamp 1676037725
transform 1 0 92736 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1000
timestamp 1676037725
transform 1 0 93104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1007
timestamp 1676037725
transform 1 0 93748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1016
timestamp 1676037725
transform 1 0 94576 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1025
timestamp 1676037725
transform 1 0 95404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1029
timestamp 1676037725
transform 1 0 95772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_1033
timestamp 1676037725
transform 1 0 96140 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1037
timestamp 1676037725
transform 1 0 96508 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1046
timestamp 1676037725
transform 1 0 97336 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1055
timestamp 1676037725
transform 1 0 98164 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1064
timestamp 1676037725
transform 1 0 98992 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1071
timestamp 1676037725
transform 1 0 99636 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1075
timestamp 1676037725
transform 1 0 100004 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1082
timestamp 1676037725
transform 1 0 100648 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1090
timestamp 1676037725
transform 1 0 101384 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1093
timestamp 1676037725
transform 1 0 101660 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1105
timestamp 1676037725
transform 1 0 102764 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1117
timestamp 1676037725
transform 1 0 103868 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1129
timestamp 1676037725
transform 1 0 104972 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_1141
timestamp 1676037725
transform 1 0 106076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_1147
timestamp 1676037725
transform 1 0 106628 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1149
timestamp 1676037725
transform 1 0 106812 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1154
timestamp 1676037725
transform 1 0 107272 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1166
timestamp 1676037725
transform 1 0 108376 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1178
timestamp 1676037725
transform 1 0 109480 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1190
timestamp 1676037725
transform 1 0 110584 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1202
timestamp 1676037725
transform 1 0 111688 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1205
timestamp 1676037725
transform 1 0 111964 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1210
timestamp 1676037725
transform 1 0 112424 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1222
timestamp 1676037725
transform 1 0 113528 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1234
timestamp 1676037725
transform 1 0 114632 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1246
timestamp 1676037725
transform 1 0 115736 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1258
timestamp 1676037725
transform 1 0 116840 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1261
timestamp 1676037725
transform 1 0 117116 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1266
timestamp 1676037725
transform 1 0 117576 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1278
timestamp 1676037725
transform 1 0 118680 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_1290
timestamp 1676037725
transform 1 0 119784 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_1298
timestamp 1676037725
transform 1 0 120520 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1305
timestamp 1676037725
transform 1 0 121164 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1314
timestamp 1676037725
transform 1 0 121992 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_1317
timestamp 1676037725
transform 1 0 122268 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1325
timestamp 1676037725
transform 1 0 123004 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1334
timestamp 1676037725
transform 1 0 123832 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1341
timestamp 1676037725
transform 1 0 124476 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1345
timestamp 1676037725
transform 1 0 124844 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1352
timestamp 1676037725
transform 1 0 125488 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1361
timestamp 1676037725
transform 1 0 126316 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1370
timestamp 1676037725
transform 1 0 127144 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1373
timestamp 1676037725
transform 1 0 127420 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1380
timestamp 1676037725
transform 1 0 128064 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_1384
timestamp 1676037725
transform 1 0 128432 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_1395
timestamp 1676037725
transform 1 0 129444 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1408
timestamp 1676037725
transform 1 0 130640 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1417
timestamp 1676037725
transform 1 0 131468 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1426
timestamp 1676037725
transform 1 0 132296 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_1429
timestamp 1676037725
transform 1 0 132572 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1435
timestamp 1676037725
transform 1 0 133124 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1439
timestamp 1676037725
transform 1 0 133492 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1446
timestamp 1676037725
transform 1 0 134136 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1454
timestamp 1676037725
transform 1 0 134872 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1466
timestamp 1676037725
transform 1 0 135976 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_1478
timestamp 1676037725
transform 1 0 137080 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1485
timestamp 1676037725
transform 1 0 137724 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_1497
timestamp 1676037725
transform 1 0 138828 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1508
timestamp 1676037725
transform 1 0 139840 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1520
timestamp 1676037725
transform 1 0 140944 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_1532
timestamp 1676037725
transform 1 0 142048 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1541
timestamp 1676037725
transform 1 0 142876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_1553
timestamp 1676037725
transform 1 0 143980 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1564
timestamp 1676037725
transform 1 0 144992 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1576
timestamp 1676037725
transform 1 0 146096 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_1588
timestamp 1676037725
transform 1 0 147200 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1597
timestamp 1676037725
transform 1 0 148028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_1609
timestamp 1676037725
transform 1 0 149132 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1620
timestamp 1676037725
transform 1 0 150144 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1632
timestamp 1676037725
transform 1 0 151248 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_1644
timestamp 1676037725
transform 1 0 152352 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1653
timestamp 1676037725
transform 1 0 153180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_1665
timestamp 1676037725
transform 1 0 154284 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_1676
timestamp 1676037725
transform 1 0 155296 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_1684
timestamp 1676037725
transform 1 0 156032 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1690
timestamp 1676037725
transform 1 0 156584 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_1699
timestamp 1676037725
transform 1 0 157412 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_1707
timestamp 1676037725
transform 1 0 158148 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1709
timestamp 1676037725
transform 1 0 158332 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1720
timestamp 1676037725
transform 1 0 159344 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1724
timestamp 1676037725
transform 1 0 159712 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_1728
timestamp 1676037725
transform 1 0 160080 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1741
timestamp 1676037725
transform 1 0 161276 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1745
timestamp 1676037725
transform 1 0 161644 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1756
timestamp 1676037725
transform 1 0 162656 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1762
timestamp 1676037725
transform 1 0 163208 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1765
timestamp 1676037725
transform 1 0 163484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1776
timestamp 1676037725
transform 1 0 164496 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1789
timestamp 1676037725
transform 1 0 165692 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1802
timestamp 1676037725
transform 1 0 166888 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1815
timestamp 1676037725
transform 1 0 168084 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_1819
timestamp 1676037725
transform 1 0 168452 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1821
timestamp 1676037725
transform 1 0 168636 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1832
timestamp 1676037725
transform 1 0 169648 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1840
timestamp 1676037725
transform 1 0 170384 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1852
timestamp 1676037725
transform 1 0 171488 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1864
timestamp 1676037725
transform 1 0 172592 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1877
timestamp 1676037725
transform 1 0 173788 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_1883
timestamp 1676037725
transform 1 0 174340 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_1891
timestamp 1676037725
transform 1 0 175076 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1896
timestamp 1676037725
transform 1 0 175536 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1912
timestamp 1676037725
transform 1 0 177008 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1920
timestamp 1676037725
transform 1 0 177744 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1933
timestamp 1676037725
transform 1 0 178940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_1945
timestamp 1676037725
transform 1 0 180044 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1952
timestamp 1676037725
transform 1 0 180688 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1968
timestamp 1676037725
transform 1 0 182160 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_1980
timestamp 1676037725
transform 1 0 183264 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1989
timestamp 1676037725
transform 1 0 184092 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2001
timestamp 1676037725
transform 1 0 185196 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2015
timestamp 1676037725
transform 1 0 186484 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2029
timestamp 1676037725
transform 1 0 187772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_2041
timestamp 1676037725
transform 1 0 188876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2045
timestamp 1676037725
transform 1 0 189244 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2057
timestamp 1676037725
transform 1 0 190348 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2066
timestamp 1676037725
transform 1 0 191176 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2075
timestamp 1676037725
transform 1 0 192004 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2084
timestamp 1676037725
transform 1 0 192832 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2093
timestamp 1676037725
transform 1 0 193660 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_2099
timestamp 1676037725
transform 1 0 194212 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2101
timestamp 1676037725
transform 1 0 194396 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2108
timestamp 1676037725
transform 1 0 195040 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2117
timestamp 1676037725
transform 1 0 195868 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_2126
timestamp 1676037725
transform 1 0 196696 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2134
timestamp 1676037725
transform 1 0 197432 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2146
timestamp 1676037725
transform 1 0 198536 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2154
timestamp 1676037725
transform 1 0 199272 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2157
timestamp 1676037725
transform 1 0 199548 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2164
timestamp 1676037725
transform 1 0 200192 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2173
timestamp 1676037725
transform 1 0 201020 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2182
timestamp 1676037725
transform 1 0 201848 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2191
timestamp 1676037725
transform 1 0 202676 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2200
timestamp 1676037725
transform 1 0 203504 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2208
timestamp 1676037725
transform 1 0 204240 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2213
timestamp 1676037725
transform 1 0 204700 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2225
timestamp 1676037725
transform 1 0 205804 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2237
timestamp 1676037725
transform 1 0 206908 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2249
timestamp 1676037725
transform 1 0 208012 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2261
timestamp 1676037725
transform 1 0 209116 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_2267
timestamp 1676037725
transform 1 0 209668 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2269
timestamp 1676037725
transform 1 0 209852 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2281
timestamp 1676037725
transform 1 0 210956 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2290
timestamp 1676037725
transform 1 0 211784 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2302
timestamp 1676037725
transform 1 0 212888 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_2314
timestamp 1676037725
transform 1 0 213992 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2322
timestamp 1676037725
transform 1 0 214728 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2325
timestamp 1676037725
transform 1 0 215004 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2337
timestamp 1676037725
transform 1 0 216108 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2346
timestamp 1676037725
transform 1 0 216936 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2358
timestamp 1676037725
transform 1 0 218040 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_2370
timestamp 1676037725
transform 1 0 219144 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2378
timestamp 1676037725
transform 1 0 219880 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2381
timestamp 1676037725
transform 1 0 220156 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2393
timestamp 1676037725
transform 1 0 221260 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2402
timestamp 1676037725
transform 1 0 222088 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2414
timestamp 1676037725
transform 1 0 223192 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2421
timestamp 1676037725
transform 1 0 223836 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2430
timestamp 1676037725
transform 1 0 224664 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2437
timestamp 1676037725
transform 1 0 225308 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2444
timestamp 1676037725
transform 1 0 225952 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2453
timestamp 1676037725
transform 1 0 226780 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2462
timestamp 1676037725
transform 1 0 227608 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2471
timestamp 1676037725
transform 1 0 228436 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2480
timestamp 1676037725
transform 1 0 229264 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_2489
timestamp 1676037725
transform 1 0 230092 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2493
timestamp 1676037725
transform 1 0 230460 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2505
timestamp 1676037725
transform 1 0 231564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2514
timestamp 1676037725
transform 1 0 232392 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2523
timestamp 1676037725
transform 1 0 233220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2532
timestamp 1676037725
transform 1 0 234048 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2541
timestamp 1676037725
transform 1 0 234876 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_2547
timestamp 1676037725
transform 1 0 235428 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2549
timestamp 1676037725
transform 1 0 235612 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2556
timestamp 1676037725
transform 1 0 236256 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2564
timestamp 1676037725
transform 1 0 236992 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2576
timestamp 1676037725
transform 1 0 238096 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2588
timestamp 1676037725
transform 1 0 239200 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2600
timestamp 1676037725
transform 1 0 240304 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2605
timestamp 1676037725
transform 1 0 240764 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_2609
timestamp 1676037725
transform 1 0 241132 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2620
timestamp 1676037725
transform 1 0 242144 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2632
timestamp 1676037725
transform 1 0 243248 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2644
timestamp 1676037725
transform 1 0 244352 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2654
timestamp 1676037725
transform 1 0 245272 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2661
timestamp 1676037725
transform 1 0 245916 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2667
timestamp 1676037725
transform 1 0 246468 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_2673
timestamp 1676037725
transform 1 0 247020 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2684
timestamp 1676037725
transform 1 0 248032 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2694
timestamp 1676037725
transform 1 0 248952 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2710
timestamp 1676037725
transform 1 0 250424 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2717
timestamp 1676037725
transform 1 0 251068 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2723
timestamp 1676037725
transform 1 0 251620 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_2729
timestamp 1676037725
transform 1 0 252172 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2740
timestamp 1676037725
transform 1 0 253184 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2756
timestamp 1676037725
transform 1 0 254656 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2770
timestamp 1676037725
transform 1 0 255944 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2773
timestamp 1676037725
transform 1 0 256220 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2785
timestamp 1676037725
transform 1 0 257324 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2799
timestamp 1676037725
transform 1 0 258612 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2808
timestamp 1676037725
transform 1 0 259440 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2817
timestamp 1676037725
transform 1 0 260268 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2826
timestamp 1676037725
transform 1 0 261096 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2829
timestamp 1676037725
transform 1 0 261372 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2837
timestamp 1676037725
transform 1 0 262108 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2847
timestamp 1676037725
transform 1 0 263028 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2856
timestamp 1676037725
transform 1 0 263856 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2870
timestamp 1676037725
transform 1 0 265144 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2878
timestamp 1676037725
transform 1 0 265880 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2882
timestamp 1676037725
transform 1 0 266248 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2885
timestamp 1676037725
transform 1 0 266524 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2893
timestamp 1676037725
transform 1 0 267260 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2903
timestamp 1676037725
transform 1 0 268180 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2913
timestamp 1676037725
transform 1 0 269100 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2917
timestamp 1676037725
transform 1 0 269468 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2925
timestamp 1676037725
transform 1 0 270204 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_2933
timestamp 1676037725
transform 1 0 270940 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_9
timestamp 1676037725
transform 1 0 1932 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_17
timestamp 1676037725
transform 1 0 2668 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_21
timestamp 1676037725
transform 1 0 3036 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_26
timestamp 1676037725
transform 1 0 3496 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_29
timestamp 1676037725
transform 1 0 3772 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_33
timestamp 1676037725
transform 1 0 4140 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_38
timestamp 1676037725
transform 1 0 4600 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_46
timestamp 1676037725
transform 1 0 5336 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 1676037725
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_65
timestamp 1676037725
transform 1 0 7084 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_73
timestamp 1676037725
transform 1 0 7820 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_77
timestamp 1676037725
transform 1 0 8188 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_82
timestamp 1676037725
transform 1 0 8648 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_85
timestamp 1676037725
transform 1 0 8924 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_89
timestamp 1676037725
transform 1 0 9292 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_94
timestamp 1676037725
transform 1 0 9752 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_102
timestamp 1676037725
transform 1 0 10488 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_110
timestamp 1676037725
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_121
timestamp 1676037725
transform 1 0 12236 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_129
timestamp 1676037725
transform 1 0 12972 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_133
timestamp 1676037725
transform 1 0 13340 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_138
timestamp 1676037725
transform 1 0 13800 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_141
timestamp 1676037725
transform 1 0 14076 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_145
timestamp 1676037725
transform 1 0 14444 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_150
timestamp 1676037725
transform 1 0 14904 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_158
timestamp 1676037725
transform 1 0 15640 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_166
timestamp 1676037725
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_177
timestamp 1676037725
transform 1 0 17388 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_185
timestamp 1676037725
transform 1 0 18124 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_193
timestamp 1676037725
transform 1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_197
timestamp 1676037725
transform 1 0 19228 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_209
timestamp 1676037725
transform 1 0 20332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_221
timestamp 1676037725
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_236
timestamp 1676037725
transform 1 0 22816 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_240
timestamp 1676037725
transform 1 0 23184 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_246
timestamp 1676037725
transform 1 0 23736 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_253
timestamp 1676037725
transform 1 0 24380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_259
timestamp 1676037725
transform 1 0 24932 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_263
timestamp 1676037725
transform 1 0 25300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_270
timestamp 1676037725
transform 1 0 25944 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_278
timestamp 1676037725
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_287
timestamp 1676037725
transform 1 0 27508 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_299
timestamp 1676037725
transform 1 0 28612 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_306
timestamp 1676037725
transform 1 0 29256 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_309
timestamp 1676037725
transform 1 0 29532 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_315
timestamp 1676037725
transform 1 0 30084 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_320
timestamp 1676037725
transform 1 0 30544 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_332
timestamp 1676037725
transform 1 0 31648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_343
timestamp 1676037725
transform 1 0 32660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_355
timestamp 1676037725
transform 1 0 33764 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_363
timestamp 1676037725
transform 1 0 34500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_365
timestamp 1676037725
transform 1 0 34684 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_376
timestamp 1676037725
transform 1 0 35696 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_383
timestamp 1676037725
transform 1 0 36340 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_390
timestamp 1676037725
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_399
timestamp 1676037725
transform 1 0 37812 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_403
timestamp 1676037725
transform 1 0 38180 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_407
timestamp 1676037725
transform 1 0 38548 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_411
timestamp 1676037725
transform 1 0 38916 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_418
timestamp 1676037725
transform 1 0 39560 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_421
timestamp 1676037725
transform 1 0 39836 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_432
timestamp 1676037725
transform 1 0 40848 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_439
timestamp 1676037725
transform 1 0 41492 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_446
timestamp 1676037725
transform 1 0 42136 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_455
timestamp 1676037725
transform 1 0 42964 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_459
timestamp 1676037725
transform 1 0 43332 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_463
timestamp 1676037725
transform 1 0 43700 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_467
timestamp 1676037725
transform 1 0 44068 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_474
timestamp 1676037725
transform 1 0 44712 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_477
timestamp 1676037725
transform 1 0 44988 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_488
timestamp 1676037725
transform 1 0 46000 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_495
timestamp 1676037725
transform 1 0 46644 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_502
timestamp 1676037725
transform 1 0 47288 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_505
timestamp 1676037725
transform 1 0 47564 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_511
timestamp 1676037725
transform 1 0 48116 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_515
timestamp 1676037725
transform 1 0 48484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_519
timestamp 1676037725
transform 1 0 48852 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_523
timestamp 1676037725
transform 1 0 49220 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_530
timestamp 1676037725
transform 1 0 49864 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_533
timestamp 1676037725
transform 1 0 50140 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_539
timestamp 1676037725
transform 1 0 50692 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_543
timestamp 1676037725
transform 1 0 51060 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_547
timestamp 1676037725
transform 1 0 51428 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_551
timestamp 1676037725
transform 1 0 51796 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_555
timestamp 1676037725
transform 1 0 52164 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_559
timestamp 1676037725
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_561
timestamp 1676037725
transform 1 0 52716 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_566
timestamp 1676037725
transform 1 0 53176 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_583
timestamp 1676037725
transform 1 0 54740 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_587
timestamp 1676037725
transform 1 0 55108 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_589
timestamp 1676037725
transform 1 0 55292 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_595
timestamp 1676037725
transform 1 0 55844 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_599
timestamp 1676037725
transform 1 0 56212 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_604
timestamp 1676037725
transform 1 0 56672 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_608
timestamp 1676037725
transform 1 0 57040 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_613
timestamp 1676037725
transform 1 0 57500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_617
timestamp 1676037725
transform 1 0 57868 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_623
timestamp 1676037725
transform 1 0 58420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_635
timestamp 1676037725
transform 1 0 59524 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_643
timestamp 1676037725
transform 1 0 60260 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_645
timestamp 1676037725
transform 1 0 60444 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_651
timestamp 1676037725
transform 1 0 60996 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_656
timestamp 1676037725
transform 1 0 61456 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_661
timestamp 1676037725
transform 1 0 61916 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_669
timestamp 1676037725
transform 1 0 62652 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_673
timestamp 1676037725
transform 1 0 63020 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_679
timestamp 1676037725
transform 1 0 63572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_691
timestamp 1676037725
transform 1 0 64676 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_699
timestamp 1676037725
transform 1 0 65412 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_701
timestamp 1676037725
transform 1 0 65596 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_713
timestamp 1676037725
transform 1 0 66700 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_725
timestamp 1676037725
transform 1 0 67804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_729
timestamp 1676037725
transform 1 0 68172 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_740
timestamp 1676037725
transform 1 0 69184 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_754
timestamp 1676037725
transform 1 0 70472 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_757
timestamp 1676037725
transform 1 0 70748 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_766
timestamp 1676037725
transform 1 0 71576 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_782
timestamp 1676037725
transform 1 0 73048 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_785
timestamp 1676037725
transform 1 0 73324 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_797
timestamp 1676037725
transform 1 0 74428 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_810
timestamp 1676037725
transform 1 0 75624 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_813
timestamp 1676037725
transform 1 0 75900 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_825
timestamp 1676037725
transform 1 0 77004 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_838
timestamp 1676037725
transform 1 0 78200 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_841
timestamp 1676037725
transform 1 0 78476 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_847
timestamp 1676037725
transform 1 0 79028 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_852
timestamp 1676037725
transform 1 0 79488 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_866
timestamp 1676037725
transform 1 0 80776 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_869
timestamp 1676037725
transform 1 0 81052 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_885
timestamp 1676037725
transform 1 0 82524 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_889
timestamp 1676037725
transform 1 0 82892 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_894
timestamp 1676037725
transform 1 0 83352 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_897
timestamp 1676037725
transform 1 0 83628 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_903
timestamp 1676037725
transform 1 0 84180 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_911
timestamp 1676037725
transform 1 0 84916 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_919
timestamp 1676037725
transform 1 0 85652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_923
timestamp 1676037725
transform 1 0 86020 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_925
timestamp 1676037725
transform 1 0 86204 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_941
timestamp 1676037725
transform 1 0 87676 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_949
timestamp 1676037725
transform 1 0 88412 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_953
timestamp 1676037725
transform 1 0 88780 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_962
timestamp 1676037725
transform 1 0 89608 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_972
timestamp 1676037725
transform 1 0 90528 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_981
timestamp 1676037725
transform 1 0 91356 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_987
timestamp 1676037725
transform 1 0 91908 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_993
timestamp 1676037725
transform 1 0 92460 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_998
timestamp 1676037725
transform 1 0 92920 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1006
timestamp 1676037725
transform 1 0 93656 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1009
timestamp 1676037725
transform 1 0 93932 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1021
timestamp 1676037725
transform 1 0 95036 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1029
timestamp 1676037725
transform 1 0 95772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1034
timestamp 1676037725
transform 1 0 96232 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1037
timestamp 1676037725
transform 1 0 96508 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_1043
timestamp 1676037725
transform 1 0 97060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1055
timestamp 1676037725
transform 1 0 98164 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1063
timestamp 1676037725
transform 1 0 98900 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1065
timestamp 1676037725
transform 1 0 99084 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_1071
timestamp 1676037725
transform 1 0 99636 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1077
timestamp 1676037725
transform 1 0 100188 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1082
timestamp 1676037725
transform 1 0 100648 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1090
timestamp 1676037725
transform 1 0 101384 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_1093
timestamp 1676037725
transform 1 0 101660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_1105
timestamp 1676037725
transform 1 0 102764 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1111
timestamp 1676037725
transform 1 0 103316 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1118
timestamp 1676037725
transform 1 0 103960 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1121
timestamp 1676037725
transform 1 0 104236 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1125
timestamp 1676037725
transform 1 0 104604 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1129
timestamp 1676037725
transform 1 0 104972 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1133
timestamp 1676037725
transform 1 0 105340 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1137
timestamp 1676037725
transform 1 0 105708 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1141
timestamp 1676037725
transform 1 0 106076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_1145
timestamp 1676037725
transform 1 0 106444 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1149
timestamp 1676037725
transform 1 0 106812 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1160
timestamp 1676037725
transform 1 0 107824 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1167
timestamp 1676037725
transform 1 0 108468 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1174
timestamp 1676037725
transform 1 0 109112 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1177
timestamp 1676037725
transform 1 0 109388 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1181
timestamp 1676037725
transform 1 0 109756 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1185
timestamp 1676037725
transform 1 0 110124 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1189
timestamp 1676037725
transform 1 0 110492 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1193
timestamp 1676037725
transform 1 0 110860 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1197
timestamp 1676037725
transform 1 0 111228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_1201
timestamp 1676037725
transform 1 0 111596 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1205
timestamp 1676037725
transform 1 0 111964 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1216
timestamp 1676037725
transform 1 0 112976 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1223
timestamp 1676037725
transform 1 0 113620 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1230
timestamp 1676037725
transform 1 0 114264 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1233
timestamp 1676037725
transform 1 0 114540 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1237
timestamp 1676037725
transform 1 0 114908 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1241
timestamp 1676037725
transform 1 0 115276 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1245
timestamp 1676037725
transform 1 0 115644 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1249
timestamp 1676037725
transform 1 0 116012 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1253
timestamp 1676037725
transform 1 0 116380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_1257
timestamp 1676037725
transform 1 0 116748 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1261
timestamp 1676037725
transform 1 0 117116 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1272
timestamp 1676037725
transform 1 0 118128 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1279
timestamp 1676037725
transform 1 0 118772 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1286
timestamp 1676037725
transform 1 0 119416 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1289
timestamp 1676037725
transform 1 0 119692 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1293
timestamp 1676037725
transform 1 0 120060 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1297
timestamp 1676037725
transform 1 0 120428 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1301
timestamp 1676037725
transform 1 0 120796 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1305
timestamp 1676037725
transform 1 0 121164 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_1313
timestamp 1676037725
transform 1 0 121900 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_1317
timestamp 1676037725
transform 1 0 122268 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_1329
timestamp 1676037725
transform 1 0 123372 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_1341
timestamp 1676037725
transform 1 0 124476 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1345
timestamp 1676037725
transform 1 0 124844 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1351
timestamp 1676037725
transform 1 0 125396 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1363
timestamp 1676037725
transform 1 0 126500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1371
timestamp 1676037725
transform 1 0 127236 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1373
timestamp 1676037725
transform 1 0 127420 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1377
timestamp 1676037725
transform 1 0 127788 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1380
timestamp 1676037725
transform 1 0 128064 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_1387
timestamp 1676037725
transform 1 0 128708 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1393
timestamp 1676037725
transform 1 0 129260 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1398
timestamp 1676037725
transform 1 0 129720 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_1401
timestamp 1676037725
transform 1 0 129996 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1411
timestamp 1676037725
transform 1 0 130916 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1419
timestamp 1676037725
transform 1 0 131652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1427
timestamp 1676037725
transform 1 0 132388 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_1429
timestamp 1676037725
transform 1 0 132572 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1435
timestamp 1676037725
transform 1 0 133124 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1440
timestamp 1676037725
transform 1 0 133584 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1448
timestamp 1676037725
transform 1 0 134320 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_1457
timestamp 1676037725
transform 1 0 135148 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_1469
timestamp 1676037725
transform 1 0 136252 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_1481
timestamp 1676037725
transform 1 0 137356 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1485
timestamp 1676037725
transform 1 0 137724 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1490
timestamp 1676037725
transform 1 0 138184 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1497
timestamp 1676037725
transform 1 0 138828 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1504
timestamp 1676037725
transform 1 0 139472 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1513
timestamp 1676037725
transform 1 0 140300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1518
timestamp 1676037725
transform 1 0 140760 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1525
timestamp 1676037725
transform 1 0 141404 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1532
timestamp 1676037725
transform 1 0 142048 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1541
timestamp 1676037725
transform 1 0 142876 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1546
timestamp 1676037725
transform 1 0 143336 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1553
timestamp 1676037725
transform 1 0 143980 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1560
timestamp 1676037725
transform 1 0 144624 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1569
timestamp 1676037725
transform 1 0 145452 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1574
timestamp 1676037725
transform 1 0 145912 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1581
timestamp 1676037725
transform 1 0 146556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1588
timestamp 1676037725
transform 1 0 147200 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1597
timestamp 1676037725
transform 1 0 148028 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1602
timestamp 1676037725
transform 1 0 148488 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1609
timestamp 1676037725
transform 1 0 149132 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1616
timestamp 1676037725
transform 1 0 149776 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1625
timestamp 1676037725
transform 1 0 150604 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1630
timestamp 1676037725
transform 1 0 151064 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1637
timestamp 1676037725
transform 1 0 151708 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1644
timestamp 1676037725
transform 1 0 152352 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1653
timestamp 1676037725
transform 1 0 153180 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1658
timestamp 1676037725
transform 1 0 153640 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1665
timestamp 1676037725
transform 1 0 154284 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1672
timestamp 1676037725
transform 1 0 154928 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1681
timestamp 1676037725
transform 1 0 155756 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1693
timestamp 1676037725
transform 1 0 156860 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_1702
timestamp 1676037725
transform 1 0 157688 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1709
timestamp 1676037725
transform 1 0 158332 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1713
timestamp 1676037725
transform 1 0 158700 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1719
timestamp 1676037725
transform 1 0 159252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1732
timestamp 1676037725
transform 1 0 160448 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1737
timestamp 1676037725
transform 1 0 160908 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1744
timestamp 1676037725
transform 1 0 161552 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1753
timestamp 1676037725
transform 1 0 162380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1762
timestamp 1676037725
transform 1 0 163208 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1765
timestamp 1676037725
transform 1 0 163484 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1772
timestamp 1676037725
transform 1 0 164128 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1781
timestamp 1676037725
transform 1 0 164956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1790
timestamp 1676037725
transform 1 0 165784 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1793
timestamp 1676037725
transform 1 0 166060 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1802
timestamp 1676037725
transform 1 0 166888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1811
timestamp 1676037725
transform 1 0 167716 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1819
timestamp 1676037725
transform 1 0 168452 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1821
timestamp 1676037725
transform 1 0 168636 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1827
timestamp 1676037725
transform 1 0 169188 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_1835
timestamp 1676037725
transform 1 0 169924 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1847
timestamp 1676037725
transform 1 0 171028 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_1849
timestamp 1676037725
transform 1 0 171212 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1855
timestamp 1676037725
transform 1 0 171764 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1859
timestamp 1676037725
transform 1 0 172132 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_1870
timestamp 1676037725
transform 1 0 173144 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1877
timestamp 1676037725
transform 1 0 173788 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1889
timestamp 1676037725
transform 1 0 174892 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_1897
timestamp 1676037725
transform 1 0 175628 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1903
timestamp 1676037725
transform 1 0 176180 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1905
timestamp 1676037725
transform 1 0 176364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1911
timestamp 1676037725
transform 1 0 176916 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1919
timestamp 1676037725
transform 1 0 177652 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1930
timestamp 1676037725
transform 1 0 178664 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1933
timestamp 1676037725
transform 1 0 178940 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1945
timestamp 1676037725
transform 1 0 180044 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_1953
timestamp 1676037725
transform 1 0 180780 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1959
timestamp 1676037725
transform 1 0 181332 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1961
timestamp 1676037725
transform 1 0 181516 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1967
timestamp 1676037725
transform 1 0 182068 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1971
timestamp 1676037725
transform 1 0 182436 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_1982
timestamp 1676037725
transform 1 0 183448 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1989
timestamp 1676037725
transform 1 0 184092 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2001
timestamp 1676037725
transform 1 0 185196 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_2013
timestamp 1676037725
transform 1 0 186300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2017
timestamp 1676037725
transform 1 0 186668 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_2029
timestamp 1676037725
transform 1 0 187772 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2035
timestamp 1676037725
transform 1 0 188324 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2039
timestamp 1676037725
transform 1 0 188692 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2043
timestamp 1676037725
transform 1 0 189060 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2045
timestamp 1676037725
transform 1 0 189244 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2057
timestamp 1676037725
transform 1 0 190348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_2065
timestamp 1676037725
transform 1 0 191084 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2071
timestamp 1676037725
transform 1 0 191636 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2073
timestamp 1676037725
transform 1 0 191820 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2079
timestamp 1676037725
transform 1 0 192372 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2087
timestamp 1676037725
transform 1 0 193108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2099
timestamp 1676037725
transform 1 0 194212 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2101
timestamp 1676037725
transform 1 0 194396 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2107
timestamp 1676037725
transform 1 0 194948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_2115
timestamp 1676037725
transform 1 0 195684 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2121
timestamp 1676037725
transform 1 0 196236 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2126
timestamp 1676037725
transform 1 0 196696 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2129
timestamp 1676037725
transform 1 0 196972 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2133
timestamp 1676037725
transform 1 0 197340 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2139
timestamp 1676037725
transform 1 0 197892 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2147
timestamp 1676037725
transform 1 0 198628 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2155
timestamp 1676037725
transform 1 0 199364 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2157
timestamp 1676037725
transform 1 0 199548 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2169
timestamp 1676037725
transform 1 0 200652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_2181
timestamp 1676037725
transform 1 0 201756 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2185
timestamp 1676037725
transform 1 0 202124 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2191
timestamp 1676037725
transform 1 0 202676 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2199
timestamp 1676037725
transform 1 0 203412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2211
timestamp 1676037725
transform 1 0 204516 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2213
timestamp 1676037725
transform 1 0 204700 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2221
timestamp 1676037725
transform 1 0 205436 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2226
timestamp 1676037725
transform 1 0 205896 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2230
timestamp 1676037725
transform 1 0 206264 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_2234
timestamp 1676037725
transform 1 0 206632 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2241
timestamp 1676037725
transform 1 0 207276 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2246
timestamp 1676037725
transform 1 0 207736 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2253
timestamp 1676037725
transform 1 0 208380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2260
timestamp 1676037725
transform 1 0 209024 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2269
timestamp 1676037725
transform 1 0 209852 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2274
timestamp 1676037725
transform 1 0 210312 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2281
timestamp 1676037725
transform 1 0 210956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2288
timestamp 1676037725
transform 1 0 211600 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2297
timestamp 1676037725
transform 1 0 212428 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2302
timestamp 1676037725
transform 1 0 212888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2309
timestamp 1676037725
transform 1 0 213532 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2316
timestamp 1676037725
transform 1 0 214176 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2325
timestamp 1676037725
transform 1 0 215004 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2330
timestamp 1676037725
transform 1 0 215464 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2337
timestamp 1676037725
transform 1 0 216108 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2344
timestamp 1676037725
transform 1 0 216752 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2353
timestamp 1676037725
transform 1 0 217580 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2358
timestamp 1676037725
transform 1 0 218040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2365
timestamp 1676037725
transform 1 0 218684 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2372
timestamp 1676037725
transform 1 0 219328 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2381
timestamp 1676037725
transform 1 0 220156 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2386
timestamp 1676037725
transform 1 0 220616 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2393
timestamp 1676037725
transform 1 0 221260 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2400
timestamp 1676037725
transform 1 0 221904 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2409
timestamp 1676037725
transform 1 0 222732 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_2414
timestamp 1676037725
transform 1 0 223192 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2420
timestamp 1676037725
transform 1 0 223744 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2425
timestamp 1676037725
transform 1 0 224204 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2432
timestamp 1676037725
transform 1 0 224848 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2437
timestamp 1676037725
transform 1 0 225308 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2449
timestamp 1676037725
transform 1 0 226412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_2461
timestamp 1676037725
transform 1 0 227516 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2465
timestamp 1676037725
transform 1 0 227884 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2471
timestamp 1676037725
transform 1 0 228436 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2479
timestamp 1676037725
transform 1 0 229172 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2483
timestamp 1676037725
transform 1 0 229540 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2488
timestamp 1676037725
transform 1 0 230000 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2493
timestamp 1676037725
transform 1 0 230460 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_2500
timestamp 1676037725
transform 1 0 231104 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2506
timestamp 1676037725
transform 1 0 231656 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2511
timestamp 1676037725
transform 1 0 232116 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2519
timestamp 1676037725
transform 1 0 232852 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2521
timestamp 1676037725
transform 1 0 233036 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2527
timestamp 1676037725
transform 1 0 233588 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_2535
timestamp 1676037725
transform 1 0 234324 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2543
timestamp 1676037725
transform 1 0 235060 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2547
timestamp 1676037725
transform 1 0 235428 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2549
timestamp 1676037725
transform 1 0 235612 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2555
timestamp 1676037725
transform 1 0 236164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2567
timestamp 1676037725
transform 1 0 237268 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2575
timestamp 1676037725
transform 1 0 238004 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2577
timestamp 1676037725
transform 1 0 238188 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2589
timestamp 1676037725
transform 1 0 239292 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2593
timestamp 1676037725
transform 1 0 239660 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_2597
timestamp 1676037725
transform 1 0 240028 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2603
timestamp 1676037725
transform 1 0 240580 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2605
timestamp 1676037725
transform 1 0 240764 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2617
timestamp 1676037725
transform 1 0 241868 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_2625
timestamp 1676037725
transform 1 0 242604 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2631
timestamp 1676037725
transform 1 0 243156 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2633
timestamp 1676037725
transform 1 0 243340 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2639
timestamp 1676037725
transform 1 0 243892 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2647
timestamp 1676037725
transform 1 0 244628 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2655
timestamp 1676037725
transform 1 0 245364 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2659
timestamp 1676037725
transform 1 0 245732 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2661
timestamp 1676037725
transform 1 0 245916 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2665
timestamp 1676037725
transform 1 0 246284 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_2676
timestamp 1676037725
transform 1 0 247296 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2686
timestamp 1676037725
transform 1 0 248216 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2689
timestamp 1676037725
transform 1 0 248492 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2697
timestamp 1676037725
transform 1 0 249228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2708
timestamp 1676037725
transform 1 0 250240 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2717
timestamp 1676037725
transform 1 0 251068 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2721
timestamp 1676037725
transform 1 0 251436 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2732
timestamp 1676037725
transform 1 0 252448 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2745
timestamp 1676037725
transform 1 0 253644 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2757
timestamp 1676037725
transform 1 0 254748 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_2769
timestamp 1676037725
transform 1 0 255852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2773
timestamp 1676037725
transform 1 0 256220 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_2785
timestamp 1676037725
transform 1 0 257324 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2796
timestamp 1676037725
transform 1 0 258336 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2801
timestamp 1676037725
transform 1 0 258796 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_2807
timestamp 1676037725
transform 1 0 259348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2813
timestamp 1676037725
transform 1 0 259900 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2817
timestamp 1676037725
transform 1 0 260268 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2826
timestamp 1676037725
transform 1 0 261096 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2829
timestamp 1676037725
transform 1 0 261372 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2836
timestamp 1676037725
transform 1 0 262016 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2845
timestamp 1676037725
transform 1 0 262844 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2854
timestamp 1676037725
transform 1 0 263672 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2857
timestamp 1676037725
transform 1 0 263948 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2865
timestamp 1676037725
transform 1 0 264684 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2885
timestamp 1676037725
transform 1 0 266524 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2894
timestamp 1676037725
transform 1 0 267352 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2903
timestamp 1676037725
transform 1 0 268180 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2916
timestamp 1676037725
transform 1 0 269376 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2923
timestamp 1676037725
transform 1 0 270020 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2934
timestamp 1676037725
transform 1 0 271032 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1
timestamp 1676037725
transform 1 0 270112 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 264040 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 263396 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1676037725
transform 1 0 264960 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1676037725
transform 1 0 264684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 262108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1676037725
transform 1 0 263028 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1676037725
transform 1 0 262752 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1676037725
transform 1 0 263396 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1676037725
transform 1 0 270756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1676037725
transform 1 0 270756 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1676037725
transform 1 0 270756 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1676037725
transform 1 0 269192 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1676037725
transform 1 0 268548 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1676037725
transform 1 0 268548 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1676037725
transform 1 0 259992 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1676037725
transform 1 0 267904 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1676037725
transform 1 0 265972 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1676037725
transform 1 0 265052 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1676037725
transform 1 0 267904 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1676037725
transform 1 0 267260 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1676037725
transform 1 0 266248 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1676037725
transform 1 0 265328 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1676037725
transform 1 0 268272 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1676037725
transform 1 0 267260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1676037725
transform 1 0 267628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1676037725
transform 1 0 260176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1676037725
transform 1 0 260636 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1676037725
transform 1 0 261740 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1676037725
transform 1 0 264408 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1676037725
transform 1 0 260176 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1676037725
transform 1 0 260820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1676037725
transform 1 0 261464 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1676037725
transform 1 0 262200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1676037725
transform 1 0 18492 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1676037725
transform 1 0 83812 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input37
timestamp 1676037725
transform 1 0 82432 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input38
timestamp 1676037725
transform 1 0 82340 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1676037725
transform 1 0 81604 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1676037725
transform 1 0 80868 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input41
timestamp 1676037725
transform 1 0 79856 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1676037725
transform 1 0 79396 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43
timestamp 1676037725
transform 1 0 78660 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp 1676037725
transform 1 0 77280 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1676037725
transform 1 0 77188 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1676037725
transform 1 0 11684 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input47
timestamp 1676037725
transform 1 0 76452 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input48
timestamp 1676037725
transform 1 0 75716 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1676037725
transform 1 0 74704 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1676037725
transform 1 0 74060 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1676037725
transform 1 0 73508 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1676037725
transform 1 0 72772 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1676037725
transform 1 0 72036 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1676037725
transform 1 0 71300 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input55
timestamp 1676037725
transform 1 0 70932 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1676037725
transform 1 0 69552 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1676037725
transform 1 0 10304 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1676037725
transform 1 0 86756 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1676037725
transform 1 0 86388 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1676037725
transform 1 0 85284 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1676037725
transform 1 0 84548 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input62
timestamp 1676037725
transform 1 0 83812 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1676037725
transform 1 0 82984 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1676037725
transform 1 0 82524 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1676037725
transform 1 0 81604 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1676037725
transform 1 0 81236 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1676037725
transform 1 0 79856 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input68
timestamp 1676037725
transform 1 0 9660 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1676037725
transform 1 0 79120 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input70
timestamp 1676037725
transform 1 0 78660 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input71
timestamp 1676037725
transform 1 0 77280 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input72
timestamp 1676037725
transform 1 0 77188 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input73
timestamp 1676037725
transform 1 0 76452 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input74
timestamp 1676037725
transform 1 0 74704 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input75
timestamp 1676037725
transform 1 0 74704 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1676037725
transform 1 0 74244 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77
timestamp 1676037725
transform 1 0 73416 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input78
timestamp 1676037725
transform 1 0 72128 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input79
timestamp 1676037725
transform 1 0 8372 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input80
timestamp 1676037725
transform 1 0 72036 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1676037725
transform 1 0 71300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input82
timestamp 1676037725
transform 1 0 69552 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1676037725
transform 1 0 69828 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1676037725
transform 1 0 120888 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1676037725
transform 1 0 120152 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1676037725
transform 1 0 119140 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1676037725
transform 1 0 118496 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1676037725
transform 1 0 117852 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1676037725
transform 1 0 117300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input90
timestamp 1676037725
transform 1 0 7728 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1676037725
transform 1 0 117944 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1676037725
transform 1 0 113988 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1676037725
transform 1 0 113344 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1676037725
transform 1 0 118588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1676037725
transform 1 0 120520 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1676037725
transform 1 0 112792 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input97
timestamp 1676037725
transform 1 0 112148 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input98
timestamp 1676037725
transform 1 0 111044 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input99
timestamp 1676037725
transform 1 0 110584 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input100
timestamp 1676037725
transform 1 0 109848 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input101
timestamp 1676037725
transform 1 0 7084 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input102
timestamp 1676037725
transform 1 0 108192 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input103
timestamp 1676037725
transform 1 0 104788 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input104
timestamp 1676037725
transform 1 0 107272 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input105
timestamp 1676037725
transform 1 0 106904 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input106
timestamp 1676037725
transform 1 0 106168 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input107
timestamp 1676037725
transform 1 0 105432 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input108
timestamp 1676037725
transform 1 0 104328 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input109
timestamp 1676037725
transform 1 0 104420 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input110
timestamp 1676037725
transform 1 0 120888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input111
timestamp 1676037725
transform 1 0 120152 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input112
timestamp 1676037725
transform 1 0 6716 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input113
timestamp 1676037725
transform 1 0 119140 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input114
timestamp 1676037725
transform 1 0 118496 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input115
timestamp 1676037725
transform 1 0 117852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input116
timestamp 1676037725
transform 1 0 117300 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input117
timestamp 1676037725
transform 1 0 116472 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input118
timestamp 1676037725
transform 1 0 115736 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input119
timestamp 1676037725
transform 1 0 115000 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input120
timestamp 1676037725
transform 1 0 113988 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input121
timestamp 1676037725
transform 1 0 113344 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input122
timestamp 1676037725
transform 1 0 112700 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input123
timestamp 1676037725
transform 1 0 5152 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input124
timestamp 1676037725
transform 1 0 112148 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input125
timestamp 1676037725
transform 1 0 111320 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input126
timestamp 1676037725
transform 1 0 110584 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input127
timestamp 1676037725
transform 1 0 109848 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input128
timestamp 1676037725
transform 1 0 108836 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input129
timestamp 1676037725
transform 1 0 108192 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input130
timestamp 1676037725
transform 1 0 107548 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input131
timestamp 1676037725
transform 1 0 106996 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input132
timestamp 1676037725
transform 1 0 106168 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input133
timestamp 1676037725
transform 1 0 105432 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input134
timestamp 1676037725
transform 1 0 5152 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input135
timestamp 1676037725
transform 1 0 104696 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input136
timestamp 1676037725
transform 1 0 103684 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input137
timestamp 1676037725
transform 1 0 159160 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input138
timestamp 1676037725
transform 1 0 158516 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input139
timestamp 1676037725
transform 1 0 155020 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input140
timestamp 1676037725
transform 1 0 154652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input141
timestamp 1676037725
transform 1 0 155020 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input142
timestamp 1676037725
transform 1 0 154008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input143
timestamp 1676037725
transform 1 0 154376 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input144
timestamp 1676037725
transform 1 0 154652 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input145
timestamp 1676037725
transform 1 0 4508 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input146
timestamp 1676037725
transform 1 0 17756 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input147
timestamp 1676037725
transform 1 0 153732 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input148
timestamp 1676037725
transform 1 0 154008 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input149
timestamp 1676037725
transform 1 0 153088 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input150
timestamp 1676037725
transform 1 0 153364 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input151
timestamp 1676037725
transform 1 0 152076 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input152
timestamp 1676037725
transform 1 0 151432 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input153
timestamp 1676037725
transform 1 0 148212 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input154
timestamp 1676037725
transform 1 0 150788 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input155
timestamp 1676037725
transform 1 0 146924 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input156
timestamp 1676037725
transform 1 0 146280 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input157
timestamp 1676037725
transform 1 0 3772 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input158
timestamp 1676037725
transform 1 0 145636 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input159
timestamp 1676037725
transform 1 0 138276 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input160
timestamp 1676037725
transform 1 0 138920 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input161
timestamp 1676037725
transform 1 0 139564 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input162
timestamp 1676037725
transform 1 0 139196 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input163
timestamp 1676037725
transform 1 0 138552 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input164
timestamp 1676037725
transform 1 0 155020 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input165
timestamp 1676037725
transform 1 0 154652 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input166
timestamp 1676037725
transform 1 0 154008 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input167
timestamp 1676037725
transform 1 0 153364 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input168
timestamp 1676037725
transform 1 0 2576 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input169
timestamp 1676037725
transform 1 0 152076 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input170
timestamp 1676037725
transform 1 0 151432 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input171
timestamp 1676037725
transform 1 0 150788 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input172
timestamp 1676037725
transform 1 0 149868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input173
timestamp 1676037725
transform 1 0 149500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input174
timestamp 1676037725
transform 1 0 148856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input175
timestamp 1676037725
transform 1 0 148212 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input176
timestamp 1676037725
transform 1 0 146924 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input177
timestamp 1676037725
transform 1 0 146280 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input178
timestamp 1676037725
transform 1 0 145636 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input179
timestamp 1676037725
transform 1 0 1840 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input180
timestamp 1676037725
transform 1 0 144716 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input181
timestamp 1676037725
transform 1 0 144348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input182
timestamp 1676037725
transform 1 0 143704 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input183
timestamp 1676037725
transform 1 0 143060 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input184
timestamp 1676037725
transform 1 0 141772 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input185
timestamp 1676037725
transform 1 0 141128 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input186
timestamp 1676037725
transform 1 0 140484 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input187
timestamp 1676037725
transform 1 0 139564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input188
timestamp 1676037725
transform 1 0 139196 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input189
timestamp 1676037725
transform 1 0 138552 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input190
timestamp 1676037725
transform 1 0 1564 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input191
timestamp 1676037725
transform 1 0 189428 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input192
timestamp 1676037725
transform 1 0 188416 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input193
timestamp 1676037725
transform 1 0 188140 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input194
timestamp 1676037725
transform 1 0 186944 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input195
timestamp 1676037725
transform 1 0 186852 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input196
timestamp 1676037725
transform 1 0 186852 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input197
timestamp 1676037725
transform 1 0 184736 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input198
timestamp 1676037725
transform 1 0 184276 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input199
timestamp 1676037725
transform 1 0 184276 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input200
timestamp 1676037725
transform 1 0 182988 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input201
timestamp 1676037725
transform 1 0 18492 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input202
timestamp 1676037725
transform 1 0 181792 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input203
timestamp 1676037725
transform 1 0 181700 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input204
timestamp 1676037725
transform 1 0 181700 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input205
timestamp 1676037725
transform 1 0 179584 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input206
timestamp 1676037725
transform 1 0 179124 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input207
timestamp 1676037725
transform 1 0 179124 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input208
timestamp 1676037725
transform 1 0 177836 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input209
timestamp 1676037725
transform 1 0 176640 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input210
timestamp 1676037725
transform 1 0 176548 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input211
timestamp 1676037725
transform 1 0 176548 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input212
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input213
timestamp 1676037725
transform 1 0 174432 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input214
timestamp 1676037725
transform 1 0 173972 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input215
timestamp 1676037725
transform 1 0 172960 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input216
timestamp 1676037725
transform 1 0 172224 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input217
timestamp 1676037725
transform 1 0 189428 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input218
timestamp 1676037725
transform 1 0 188416 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input219
timestamp 1676037725
transform 1 0 189428 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input220
timestamp 1676037725
transform 1 0 186944 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input221
timestamp 1676037725
transform 1 0 186852 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input222
timestamp 1676037725
transform 1 0 186852 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input223
timestamp 1676037725
transform 1 0 17020 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input224
timestamp 1676037725
transform 1 0 185564 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input225
timestamp 1676037725
transform 1 0 184276 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input226
timestamp 1676037725
transform 1 0 184276 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input227
timestamp 1676037725
transform 1 0 182528 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input228
timestamp 1676037725
transform 1 0 181792 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input229
timestamp 1676037725
transform 1 0 181700 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input230
timestamp 1676037725
transform 1 0 180320 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input231
timestamp 1676037725
transform 1 0 180412 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input232
timestamp 1676037725
transform 1 0 179124 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input233
timestamp 1676037725
transform 1 0 177744 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input234
timestamp 1676037725
transform 1 0 16008 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input235
timestamp 1676037725
transform 1 0 177376 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input236
timestamp 1676037725
transform 1 0 176640 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input237
timestamp 1676037725
transform 1 0 176548 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input238
timestamp 1676037725
transform 1 0 175168 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input239
timestamp 1676037725
transform 1 0 175260 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input240
timestamp 1676037725
transform 1 0 173972 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input241
timestamp 1676037725
transform 1 0 173972 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input242
timestamp 1676037725
transform 1 0 172224 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input243
timestamp 1676037725
transform 1 0 224480 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input244
timestamp 1676037725
transform 1 0 226964 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input245
timestamp 1676037725
transform 1 0 15272 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input246
timestamp 1676037725
transform 1 0 226320 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input247
timestamp 1676037725
transform 1 0 225676 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input248
timestamp 1676037725
transform 1 0 226228 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input249
timestamp 1676037725
transform 1 0 224756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input250
timestamp 1676037725
transform 1 0 220340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input251
timestamp 1676037725
transform 1 0 222916 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input252
timestamp 1676037725
transform 1 0 220340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input253
timestamp 1676037725
transform 1 0 216936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input254
timestamp 1676037725
transform 1 0 222916 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input255
timestamp 1676037725
transform 1 0 215188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input256
timestamp 1676037725
transform 1 0 14536 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input257
timestamp 1676037725
transform 1 0 17020 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input258
timestamp 1676037725
transform 1 0 220340 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input259
timestamp 1676037725
transform 1 0 219328 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input260
timestamp 1676037725
transform 1 0 218684 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input261
timestamp 1676037725
transform 1 0 214360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input262
timestamp 1676037725
transform 1 0 213716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input263
timestamp 1676037725
transform 1 0 208104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input264
timestamp 1676037725
transform 1 0 207644 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input265
timestamp 1676037725
transform 1 0 208288 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input266
timestamp 1676037725
transform 1 0 208748 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input267
timestamp 1676037725
transform 1 0 208104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input268
timestamp 1676037725
transform 1 0 13432 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input269
timestamp 1676037725
transform 1 0 207460 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input270
timestamp 1676037725
transform 1 0 206356 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input271
timestamp 1676037725
transform 1 0 224572 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input272
timestamp 1676037725
transform 1 0 222916 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input273
timestamp 1676037725
transform 1 0 221812 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input274
timestamp 1676037725
transform 1 0 221628 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input275
timestamp 1676037725
transform 1 0 220984 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input276
timestamp 1676037725
transform 1 0 220340 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input277
timestamp 1676037725
transform 1 0 219052 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input278
timestamp 1676037725
transform 1 0 218408 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input279
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input280
timestamp 1676037725
transform 1 0 217764 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input281
timestamp 1676037725
transform 1 0 216660 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input282
timestamp 1676037725
transform 1 0 216476 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input283
timestamp 1676037725
transform 1 0 215832 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input284
timestamp 1676037725
transform 1 0 215188 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input285
timestamp 1676037725
transform 1 0 213900 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input286
timestamp 1676037725
transform 1 0 213256 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input287
timestamp 1676037725
transform 1 0 212612 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input288
timestamp 1676037725
transform 1 0 211508 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input289
timestamp 1676037725
transform 1 0 211324 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input290
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input291
timestamp 1676037725
transform 1 0 210680 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input292
timestamp 1676037725
transform 1 0 210036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input293
timestamp 1676037725
transform 1 0 208748 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input294
timestamp 1676037725
transform 1 0 208104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input295
timestamp 1676037725
transform 1 0 207460 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input296
timestamp 1676037725
transform 1 0 206356 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input297
timestamp 1676037725
transform 1 0 258704 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input298
timestamp 1676037725
transform 1 0 258980 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input299
timestamp 1676037725
transform 1 0 257416 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input300
timestamp 1676037725
transform 1 0 258980 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input301
timestamp 1676037725
transform 1 0 11868 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input302
timestamp 1676037725
transform 1 0 254840 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input303
timestamp 1676037725
transform 1 0 256404 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input304
timestamp 1676037725
transform 1 0 253828 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input305
timestamp 1676037725
transform 1 0 253552 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input306
timestamp 1676037725
transform 1 0 253828 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input307
timestamp 1676037725
transform 1 0 251252 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input308
timestamp 1676037725
transform 1 0 253828 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input309
timestamp 1676037725
transform 1 0 252264 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input310
timestamp 1676037725
transform 1 0 250976 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input311
timestamp 1676037725
transform 1 0 251252 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input312
timestamp 1676037725
transform 1 0 10856 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input313
timestamp 1676037725
transform 1 0 247020 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input314
timestamp 1676037725
transform 1 0 247204 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input315
timestamp 1676037725
transform 1 0 247112 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input316
timestamp 1676037725
transform 1 0 246100 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input317
timestamp 1676037725
transform 1 0 244720 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input318
timestamp 1676037725
transform 1 0 243432 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input319
timestamp 1676037725
transform 1 0 243524 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input320
timestamp 1676037725
transform 1 0 243524 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input321
timestamp 1676037725
transform 1 0 241224 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input322
timestamp 1676037725
transform 1 0 240948 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input323
timestamp 1676037725
transform 1 0 10120 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input324
timestamp 1676037725
transform 1 0 257692 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input325
timestamp 1676037725
transform 1 0 256680 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input326
timestamp 1676037725
transform 1 0 256404 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input327
timestamp 1676037725
transform 1 0 256404 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input328
timestamp 1676037725
transform 1 0 255024 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input329
timestamp 1676037725
transform 1 0 253736 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input330
timestamp 1676037725
transform 1 0 253828 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input331
timestamp 1676037725
transform 1 0 252264 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input332
timestamp 1676037725
transform 1 0 251528 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input333
timestamp 1676037725
transform 1 0 251252 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input334
timestamp 1676037725
transform 1 0 9384 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input335
timestamp 1676037725
transform 1 0 250056 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input336
timestamp 1676037725
transform 1 0 249320 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input337
timestamp 1676037725
transform 1 0 248584 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input338
timestamp 1676037725
transform 1 0 247848 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input339
timestamp 1676037725
transform 1 0 247112 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input340
timestamp 1676037725
transform 1 0 246376 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input341
timestamp 1676037725
transform 1 0 246100 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input342
timestamp 1676037725
transform 1 0 244904 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input343
timestamp 1676037725
transform 1 0 244996 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input344
timestamp 1676037725
transform 1 0 244260 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input345
timestamp 1676037725
transform 1 0 8280 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input346
timestamp 1676037725
transform 1 0 243524 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input347
timestamp 1676037725
transform 1 0 242236 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input348
timestamp 1676037725
transform 1 0 241224 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input349
timestamp 1676037725
transform 1 0 240948 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input350
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input351
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input352
timestamp 1676037725
transform 1 0 15456 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input353
timestamp 1676037725
transform 1 0 6716 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input354
timestamp 1676037725
transform 1 0 5704 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input355
timestamp 1676037725
transform 1 0 4968 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input356
timestamp 1676037725
transform 1 0 4232 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input357
timestamp 1676037725
transform 1 0 3128 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input358
timestamp 1676037725
transform 1 0 3036 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input359
timestamp 1676037725
transform 1 0 2300 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input360
timestamp 1676037725
transform 1 0 1564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input361
timestamp 1676037725
transform 1 0 52900 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input362
timestamp 1676037725
transform 1 0 51888 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input363
timestamp 1676037725
transform 1 0 15456 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input364
timestamp 1676037725
transform 1 0 51152 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input365
timestamp 1676037725
transform 1 0 50416 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input366
timestamp 1676037725
transform 1 0 49588 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input367
timestamp 1676037725
transform 1 0 48944 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input368
timestamp 1676037725
transform 1 0 48208 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input369
timestamp 1676037725
transform 1 0 47012 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input370
timestamp 1676037725
transform 1 0 46368 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input371
timestamp 1676037725
transform 1 0 45724 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input372
timestamp 1676037725
transform 1 0 45264 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input373
timestamp 1676037725
transform 1 0 44436 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input374
timestamp 1676037725
transform 1 0 14812 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input375
timestamp 1676037725
transform 1 0 43792 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input376
timestamp 1676037725
transform 1 0 43056 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input377
timestamp 1676037725
transform 1 0 41860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input378
timestamp 1676037725
transform 1 0 41216 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input379
timestamp 1676037725
transform 1 0 40572 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input380
timestamp 1676037725
transform 1 0 39284 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input381
timestamp 1676037725
transform 1 0 38640 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input382
timestamp 1676037725
transform 1 0 37996 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input383
timestamp 1676037725
transform 1 0 37904 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input384
timestamp 1676037725
transform 1 0 36708 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input385
timestamp 1676037725
transform 1 0 14076 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input386
timestamp 1676037725
transform 1 0 36064 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input387
timestamp 1676037725
transform 1 0 35420 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input388
timestamp 1676037725
transform 1 0 52900 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input389
timestamp 1676037725
transform 1 0 51888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input390
timestamp 1676037725
transform 1 0 51152 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input391
timestamp 1676037725
transform 1 0 50416 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input392
timestamp 1676037725
transform 1 0 49588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input393
timestamp 1676037725
transform 1 0 48944 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input394
timestamp 1676037725
transform 1 0 48208 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input395
timestamp 1676037725
transform 1 0 47012 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input396
timestamp 1676037725
transform 1 0 13340 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input397
timestamp 1676037725
transform 1 0 46368 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input398
timestamp 1676037725
transform 1 0 45724 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input399
timestamp 1676037725
transform 1 0 45264 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input400
timestamp 1676037725
transform 1 0 44436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input401
timestamp 1676037725
transform 1 0 43792 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input402
timestamp 1676037725
transform 1 0 43056 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input403
timestamp 1676037725
transform 1 0 41860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input404
timestamp 1676037725
transform 1 0 41216 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input405
timestamp 1676037725
transform 1 0 40572 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input406
timestamp 1676037725
transform 1 0 40112 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input407
timestamp 1676037725
transform 1 0 12604 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input408
timestamp 1676037725
transform 1 0 39284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input409
timestamp 1676037725
transform 1 0 38640 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input410
timestamp 1676037725
transform 1 0 37904 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input411
timestamp 1676037725
transform 1 0 36708 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input412
timestamp 1676037725
transform 1 0 36064 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input413
timestamp 1676037725
transform 1 0 35420 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input414
timestamp 1676037725
transform 1 0 86756 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input415
timestamp 1676037725
transform 1 0 86020 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input416
timestamp 1676037725
transform 1 0 85008 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input417
timestamp 1676037725
transform 1 0 84548 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input418
timestamp 1676037725
transform 1 0 11868 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 271492 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 271492 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 271492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 271492 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 271492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 271492 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 271492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 271492 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 271492 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 271492 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 271492 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 271492 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 271492 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 271492 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 271492 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 271492 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1676037725
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1676037725
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1676037725
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1676037725
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1676037725
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1676037725
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1676037725
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1676037725
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1676037725
transform 1 0 26864 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1676037725
transform 1 0 29440 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1676037725
transform 1 0 32016 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1676037725
transform 1 0 34592 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1676037725
transform 1 0 37168 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1676037725
transform 1 0 39744 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1676037725
transform 1 0 42320 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1676037725
transform 1 0 44896 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1676037725
transform 1 0 47472 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1676037725
transform 1 0 50048 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1676037725
transform 1 0 52624 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1676037725
transform 1 0 55200 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1676037725
transform 1 0 57776 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1676037725
transform 1 0 60352 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1676037725
transform 1 0 62928 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1676037725
transform 1 0 65504 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1676037725
transform 1 0 68080 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1676037725
transform 1 0 70656 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1676037725
transform 1 0 73232 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1676037725
transform 1 0 75808 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1676037725
transform 1 0 78384 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1676037725
transform 1 0 80960 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1676037725
transform 1 0 83536 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1676037725
transform 1 0 86112 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1676037725
transform 1 0 88688 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1676037725
transform 1 0 91264 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1676037725
transform 1 0 93840 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1676037725
transform 1 0 96416 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1676037725
transform 1 0 98992 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1676037725
transform 1 0 101568 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1676037725
transform 1 0 104144 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1676037725
transform 1 0 106720 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1676037725
transform 1 0 109296 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1676037725
transform 1 0 111872 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1676037725
transform 1 0 114448 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1676037725
transform 1 0 117024 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1676037725
transform 1 0 119600 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1676037725
transform 1 0 122176 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1676037725
transform 1 0 124752 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1676037725
transform 1 0 127328 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1676037725
transform 1 0 129904 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1676037725
transform 1 0 132480 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 135056 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 137632 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 140208 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 142784 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 145360 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 147936 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 150512 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 153088 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 155664 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 158240 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 160816 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 163392 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 165968 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 168544 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 171120 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 173696 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 176272 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 178848 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 181424 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 184000 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 186576 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 189152 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 191728 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 194304 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 196880 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 199456 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 202032 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 204608 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 207184 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 209760 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 212336 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 214912 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 217488 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 220064 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 222640 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 225216 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 227792 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 230368 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 232944 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 235520 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 238096 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 240672 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 243248 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 245824 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 248400 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 250976 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 253552 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 256128 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 258704 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 261280 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 263856 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 266432 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 269008 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 26864 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 32016 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 37168 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 42320 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 47472 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 52624 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 57776 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 62928 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 68080 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 73232 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 78384 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 83536 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 88688 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 93840 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 98992 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 104144 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 109296 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 114448 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 119600 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 124752 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 129904 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 135056 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 140208 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 145360 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 150512 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 155664 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 160816 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 165968 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 171120 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 176272 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 181424 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 186576 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 191728 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 196880 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 202032 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 207184 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 212336 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 217488 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 222640 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 227792 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 232944 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 238096 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 243248 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 248400 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 253552 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 258704 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 263856 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 269008 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 80960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 86112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 91264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 96416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 101568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 106720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 111872 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 117024 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 122176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 127328 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 132480 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 137632 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 142784 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 147936 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 153088 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 158240 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 163392 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 168544 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 173696 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 178848 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 184000 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 189152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 194304 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 199456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 204608 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 209760 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 214912 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 220064 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 225216 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 230368 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 235520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 240672 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 245824 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 250976 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 256128 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 261280 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 266432 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 83536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 88688 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 93840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 98992 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 104144 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 109296 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 114448 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 119600 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 124752 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 129904 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 135056 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 140208 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 145360 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 150512 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 155664 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 160816 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 165968 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 171120 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 176272 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 181424 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 186576 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 191728 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 196880 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 202032 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 207184 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 212336 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 217488 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 222640 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 227792 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 232944 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 238096 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 243248 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 248400 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 253552 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 258704 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 263856 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 269008 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 80960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 86112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 91264 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 96416 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 101568 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 106720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 111872 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 117024 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 122176 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 127328 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 132480 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 137632 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 142784 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 147936 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 153088 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 158240 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 163392 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 168544 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 173696 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 178848 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 184000 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 189152 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 194304 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 199456 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 204608 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 209760 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 214912 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 220064 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 225216 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 230368 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 235520 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 240672 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 245824 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 250976 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 256128 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 261280 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 266432 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 83536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 88688 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 93840 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 98992 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 104144 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 109296 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 114448 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 119600 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 124752 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 129904 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 135056 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 140208 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 145360 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 150512 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 155664 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 160816 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 165968 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 171120 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 176272 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 181424 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 186576 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 191728 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 196880 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 202032 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 207184 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 212336 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 217488 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 222640 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 227792 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 232944 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 238096 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 243248 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 248400 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 253552 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 258704 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 263856 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 269008 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 80960 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 86112 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 91264 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 96416 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 101568 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 106720 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 111872 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 117024 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 122176 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 127328 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 132480 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 137632 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 142784 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 147936 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 153088 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 158240 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 163392 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 168544 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 173696 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 178848 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 184000 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 189152 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 194304 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 199456 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 204608 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 209760 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 214912 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 220064 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 225216 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 230368 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 235520 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 240672 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 245824 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 250976 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 256128 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 261280 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 266432 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 83536 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 88688 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 93840 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 98992 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 104144 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 109296 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 114448 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 119600 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 124752 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 129904 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 135056 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 140208 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 145360 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 150512 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 155664 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 160816 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 165968 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 171120 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 176272 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 181424 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 186576 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 191728 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 196880 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 202032 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 207184 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 212336 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 217488 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 222640 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 227792 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 232944 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 238096 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 243248 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 248400 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 253552 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 258704 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 263856 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 269008 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 80960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 86112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 91264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 96416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 101568 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 106720 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 111872 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 117024 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 122176 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 127328 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 132480 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 137632 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 142784 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 147936 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 153088 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 158240 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 163392 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 168544 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 173696 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 178848 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 184000 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 189152 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 194304 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 199456 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 204608 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 209760 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 214912 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 220064 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 225216 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 230368 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 235520 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 240672 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 245824 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 250976 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 256128 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 261280 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 266432 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 78384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 83536 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 88688 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 93840 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 98992 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 104144 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 109296 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 114448 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 119600 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 124752 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 129904 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 135056 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 140208 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 145360 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 150512 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 155664 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 160816 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 165968 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 171120 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 176272 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 181424 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 186576 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 191728 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 196880 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 202032 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 207184 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 212336 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 217488 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 222640 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 227792 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 232944 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 238096 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 243248 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 248400 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 253552 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 258704 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 263856 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 269008 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 70656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 75808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 80960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 86112 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 91264 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 96416 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 101568 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 106720 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 111872 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 117024 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 122176 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 127328 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 132480 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 137632 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 142784 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 147936 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1676037725
transform 1 0 153088 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1676037725
transform 1 0 158240 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1676037725
transform 1 0 163392 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1676037725
transform 1 0 168544 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1676037725
transform 1 0 173696 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1676037725
transform 1 0 178848 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1676037725
transform 1 0 184000 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1676037725
transform 1 0 189152 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1676037725
transform 1 0 194304 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1676037725
transform 1 0 199456 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1676037725
transform 1 0 204608 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1676037725
transform 1 0 209760 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1676037725
transform 1 0 214912 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1676037725
transform 1 0 220064 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1676037725
transform 1 0 225216 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1676037725
transform 1 0 230368 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1676037725
transform 1 0 235520 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1676037725
transform 1 0 240672 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1676037725
transform 1 0 245824 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1676037725
transform 1 0 250976 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1676037725
transform 1 0 256128 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1676037725
transform 1 0 261280 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1676037725
transform 1 0 266432 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1676037725
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1676037725
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1676037725
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1676037725
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1676037725
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1676037725
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1676037725
transform 1 0 78384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1676037725
transform 1 0 83536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1676037725
transform 1 0 88688 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1676037725
transform 1 0 93840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1676037725
transform 1 0 98992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1676037725
transform 1 0 104144 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1676037725
transform 1 0 109296 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1676037725
transform 1 0 114448 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1676037725
transform 1 0 119600 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1676037725
transform 1 0 124752 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1676037725
transform 1 0 129904 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1676037725
transform 1 0 135056 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1676037725
transform 1 0 140208 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1676037725
transform 1 0 145360 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1676037725
transform 1 0 150512 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1676037725
transform 1 0 155664 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1676037725
transform 1 0 160816 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1676037725
transform 1 0 165968 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1676037725
transform 1 0 171120 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1676037725
transform 1 0 176272 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1676037725
transform 1 0 181424 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1676037725
transform 1 0 186576 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1676037725
transform 1 0 191728 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1676037725
transform 1 0 196880 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1676037725
transform 1 0 202032 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1676037725
transform 1 0 207184 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1676037725
transform 1 0 212336 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1676037725
transform 1 0 217488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1676037725
transform 1 0 222640 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1676037725
transform 1 0 227792 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1676037725
transform 1 0 232944 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1676037725
transform 1 0 238096 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1676037725
transform 1 0 243248 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1676037725
transform 1 0 248400 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1676037725
transform 1 0 253552 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1676037725
transform 1 0 258704 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1676037725
transform 1 0 263856 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1676037725
transform 1 0 269008 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1676037725
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1676037725
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1676037725
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1676037725
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1676037725
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1676037725
transform 1 0 70656 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1676037725
transform 1 0 75808 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1676037725
transform 1 0 80960 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1676037725
transform 1 0 86112 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1676037725
transform 1 0 91264 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1676037725
transform 1 0 96416 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1676037725
transform 1 0 101568 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1676037725
transform 1 0 106720 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1676037725
transform 1 0 111872 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1676037725
transform 1 0 117024 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1676037725
transform 1 0 122176 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1676037725
transform 1 0 127328 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1676037725
transform 1 0 132480 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1676037725
transform 1 0 137632 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1676037725
transform 1 0 142784 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1676037725
transform 1 0 147936 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1676037725
transform 1 0 153088 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1676037725
transform 1 0 158240 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1676037725
transform 1 0 163392 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1676037725
transform 1 0 168544 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1676037725
transform 1 0 173696 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1676037725
transform 1 0 178848 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1676037725
transform 1 0 184000 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1676037725
transform 1 0 189152 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1676037725
transform 1 0 194304 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1676037725
transform 1 0 199456 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1676037725
transform 1 0 204608 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1676037725
transform 1 0 209760 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1676037725
transform 1 0 214912 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1676037725
transform 1 0 220064 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1676037725
transform 1 0 225216 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1676037725
transform 1 0 230368 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1676037725
transform 1 0 235520 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1676037725
transform 1 0 240672 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1676037725
transform 1 0 245824 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1676037725
transform 1 0 250976 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1676037725
transform 1 0 256128 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1676037725
transform 1 0 261280 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1676037725
transform 1 0 266432 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1676037725
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1676037725
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1676037725
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1676037725
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1676037725
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1676037725
transform 1 0 73232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1676037725
transform 1 0 78384 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1676037725
transform 1 0 83536 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1676037725
transform 1 0 88688 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1676037725
transform 1 0 93840 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1676037725
transform 1 0 98992 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1676037725
transform 1 0 104144 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1676037725
transform 1 0 109296 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1676037725
transform 1 0 114448 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1676037725
transform 1 0 119600 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1676037725
transform 1 0 124752 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1676037725
transform 1 0 129904 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1676037725
transform 1 0 135056 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1676037725
transform 1 0 140208 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1676037725
transform 1 0 145360 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1676037725
transform 1 0 150512 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1676037725
transform 1 0 155664 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1676037725
transform 1 0 160816 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1676037725
transform 1 0 165968 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1676037725
transform 1 0 171120 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1676037725
transform 1 0 176272 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1676037725
transform 1 0 181424 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1676037725
transform 1 0 186576 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1676037725
transform 1 0 191728 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1676037725
transform 1 0 196880 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1676037725
transform 1 0 202032 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1676037725
transform 1 0 207184 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1676037725
transform 1 0 212336 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1676037725
transform 1 0 217488 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1676037725
transform 1 0 222640 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1676037725
transform 1 0 227792 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1676037725
transform 1 0 232944 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1676037725
transform 1 0 238096 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1676037725
transform 1 0 243248 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1676037725
transform 1 0 248400 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1676037725
transform 1 0 253552 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1676037725
transform 1 0 258704 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1676037725
transform 1 0 263856 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1676037725
transform 1 0 269008 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1676037725
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1676037725
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1676037725
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1676037725
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1676037725
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1676037725
transform 1 0 70656 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1676037725
transform 1 0 75808 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1676037725
transform 1 0 80960 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1676037725
transform 1 0 86112 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1676037725
transform 1 0 91264 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1676037725
transform 1 0 96416 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1676037725
transform 1 0 101568 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1676037725
transform 1 0 106720 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1676037725
transform 1 0 111872 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1676037725
transform 1 0 117024 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1676037725
transform 1 0 122176 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1676037725
transform 1 0 127328 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1676037725
transform 1 0 132480 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1676037725
transform 1 0 137632 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1676037725
transform 1 0 142784 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1676037725
transform 1 0 147936 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1676037725
transform 1 0 153088 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1676037725
transform 1 0 158240 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1676037725
transform 1 0 163392 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1676037725
transform 1 0 168544 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1676037725
transform 1 0 173696 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1676037725
transform 1 0 178848 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1676037725
transform 1 0 184000 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1676037725
transform 1 0 189152 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1676037725
transform 1 0 194304 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1676037725
transform 1 0 199456 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1676037725
transform 1 0 204608 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1676037725
transform 1 0 209760 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1676037725
transform 1 0 214912 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1676037725
transform 1 0 220064 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1676037725
transform 1 0 225216 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1676037725
transform 1 0 230368 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1676037725
transform 1 0 235520 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1676037725
transform 1 0 240672 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1676037725
transform 1 0 245824 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1676037725
transform 1 0 250976 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1676037725
transform 1 0 256128 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1676037725
transform 1 0 261280 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1676037725
transform 1 0 266432 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1676037725
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1676037725
transform 1 0 8832 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1676037725
transform 1 0 13984 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1676037725
transform 1 0 19136 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1676037725
transform 1 0 24288 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1676037725
transform 1 0 29440 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1676037725
transform 1 0 34592 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1676037725
transform 1 0 39744 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1676037725
transform 1 0 44896 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1676037725
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1676037725
transform 1 0 50048 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1676037725
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1676037725
transform 1 0 55200 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1676037725
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1676037725
transform 1 0 60352 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1676037725
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1676037725
transform 1 0 65504 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1676037725
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1676037725
transform 1 0 70656 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1676037725
transform 1 0 73232 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1676037725
transform 1 0 75808 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1676037725
transform 1 0 78384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1676037725
transform 1 0 80960 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1676037725
transform 1 0 83536 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1676037725
transform 1 0 86112 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1676037725
transform 1 0 88688 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1676037725
transform 1 0 91264 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1676037725
transform 1 0 93840 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1676037725
transform 1 0 96416 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1676037725
transform 1 0 98992 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1676037725
transform 1 0 101568 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1676037725
transform 1 0 104144 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1676037725
transform 1 0 106720 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1676037725
transform 1 0 109296 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1676037725
transform 1 0 111872 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1676037725
transform 1 0 114448 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1676037725
transform 1 0 117024 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1676037725
transform 1 0 119600 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1676037725
transform 1 0 122176 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1676037725
transform 1 0 124752 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1676037725
transform 1 0 127328 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1676037725
transform 1 0 129904 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1676037725
transform 1 0 132480 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1676037725
transform 1 0 135056 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1676037725
transform 1 0 137632 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1676037725
transform 1 0 140208 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1676037725
transform 1 0 142784 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1676037725
transform 1 0 145360 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1676037725
transform 1 0 147936 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1676037725
transform 1 0 150512 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1676037725
transform 1 0 153088 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1676037725
transform 1 0 155664 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1676037725
transform 1 0 158240 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1676037725
transform 1 0 160816 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1676037725
transform 1 0 163392 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1676037725
transform 1 0 165968 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1676037725
transform 1 0 168544 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1676037725
transform 1 0 171120 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1676037725
transform 1 0 173696 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1676037725
transform 1 0 176272 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1676037725
transform 1 0 178848 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1676037725
transform 1 0 181424 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1676037725
transform 1 0 184000 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1676037725
transform 1 0 186576 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1676037725
transform 1 0 189152 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1676037725
transform 1 0 191728 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1676037725
transform 1 0 194304 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1676037725
transform 1 0 196880 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1676037725
transform 1 0 199456 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1676037725
transform 1 0 202032 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1676037725
transform 1 0 204608 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1676037725
transform 1 0 207184 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1676037725
transform 1 0 209760 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1676037725
transform 1 0 212336 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1676037725
transform 1 0 214912 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1676037725
transform 1 0 217488 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1676037725
transform 1 0 220064 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1676037725
transform 1 0 222640 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1676037725
transform 1 0 225216 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1676037725
transform 1 0 227792 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1676037725
transform 1 0 230368 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1676037725
transform 1 0 232944 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1676037725
transform 1 0 235520 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1676037725
transform 1 0 238096 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1676037725
transform 1 0 240672 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1676037725
transform 1 0 243248 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1676037725
transform 1 0 245824 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1676037725
transform 1 0 248400 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1676037725
transform 1 0 250976 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1676037725
transform 1 0 253552 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1676037725
transform 1 0 256128 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1676037725
transform 1 0 258704 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1676037725
transform 1 0 261280 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1676037725
transform 1 0 263856 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1676037725
transform 1 0 266432 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1676037725
transform 1 0 269008 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  tt_mux_517
timestamp 1676037725
transform 1 0 259348 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_518
timestamp 1676037725
transform 1 0 265604 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_519
timestamp 1676037725
transform 1 0 265972 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_520
timestamp 1676037725
transform 1 0 1564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_521
timestamp 1676037725
transform 1 0 1564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_522
timestamp 1676037725
transform 1 0 34960 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_523
timestamp 1676037725
transform 1 0 34960 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_524
timestamp 1676037725
transform 1 0 68908 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_525
timestamp 1676037725
transform 1 0 68908 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_526
timestamp 1676037725
transform 1 0 103500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_527
timestamp 1676037725
transform 1 0 103040 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_528
timestamp 1676037725
transform 1 0 137908 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_529
timestamp 1676037725
transform 1 0 137908 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_530
timestamp 1676037725
transform 1 0 171488 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_531
timestamp 1676037725
transform 1 0 171488 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_532
timestamp 1676037725
transform 1 0 205620 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_533
timestamp 1676037725
transform 1 0 205620 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_534
timestamp 1676037725
transform 1 0 239752 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_535
timestamp 1676037725
transform 1 0 239752 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_552
timestamp 1676037725
transform 1 0 265972 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 252724 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_8  zbuf_bus_ena_I.genblk1.cell1_I
timestamp 1676037725
transform 1 0 238188 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 267904 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[0\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 267904 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 269284 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[1\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 269284 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 269468 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[2\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 268272 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 267904 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[3\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 267720 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 267076 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[4\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 266800 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 266708 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[5\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 266524 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 266432 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[6\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 265328 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 267352 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[7\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 264316 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 268180 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[8\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 263672 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 264868 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[9\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 264132 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 262752 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[10\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 262844 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 262108 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[11\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 261556 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 260728 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[12\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 261556 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 259900 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[13\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 260268 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 270112 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[14\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 260912 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 266892 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[15\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 259716 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 267720 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[16\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 266800 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 269652 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[17\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 268456 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_sel_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 249964 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_sel_I\[0\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 226596 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_sel_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 252724 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  zbuf_bus_sel_I\[1\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 223744 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  zbuf_bus_sel_I\[2\].genblk1.cell0_I openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 251712 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  zbuf_bus_sel_I\[2\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 213256 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_2  zbuf_bus_sel_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 250792 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  zbuf_bus_sel_I\[3\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 212980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_2  zbuf_bus_sel_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 251252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  zbuf_bus_sel_I\[4\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 212888 0 -1 6528
box -38 -48 1142 592
<< labels >>
flabel metal3 s 272304 9558 272504 9618 0 FreeSans 480 0 0 0 addr[0]
port 0 nsew signal input
flabel metal3 s 272304 9422 272504 9482 0 FreeSans 480 0 0 0 addr[1]
port 1 nsew signal input
flabel metal3 s 272304 9286 272504 9346 0 FreeSans 480 0 0 0 addr[2]
port 2 nsew signal input
flabel metal3 s 272304 9150 272504 9210 0 FreeSans 480 0 0 0 addr[3]
port 3 nsew signal input
flabel metal3 s 272304 9014 272504 9074 0 FreeSans 480 0 0 0 addr[4]
port 4 nsew signal input
flabel metal3 s 272304 8878 272504 8938 0 FreeSans 480 0 0 0 k_one
port 5 nsew signal tristate
flabel metal3 s 272304 8742 272504 8802 0 FreeSans 480 0 0 0 k_zero
port 6 nsew signal tristate
flabel metal3 s 272304 8606 272504 8666 0 FreeSans 480 0 0 0 spine_iw[0]
port 7 nsew signal input
flabel metal3 s 272304 7246 272504 7306 0 FreeSans 480 0 0 0 spine_iw[10]
port 8 nsew signal input
flabel metal3 s 272304 7110 272504 7170 0 FreeSans 480 0 0 0 spine_iw[11]
port 9 nsew signal input
flabel metal3 s 272304 6974 272504 7034 0 FreeSans 480 0 0 0 spine_iw[12]
port 10 nsew signal input
flabel metal3 s 272304 6838 272504 6898 0 FreeSans 480 0 0 0 spine_iw[13]
port 11 nsew signal input
flabel metal3 s 272304 6702 272504 6762 0 FreeSans 480 0 0 0 spine_iw[14]
port 12 nsew signal input
flabel metal3 s 272304 6566 272504 6626 0 FreeSans 480 0 0 0 spine_iw[15]
port 13 nsew signal input
flabel metal3 s 272304 6430 272504 6490 0 FreeSans 480 0 0 0 spine_iw[16]
port 14 nsew signal input
flabel metal3 s 272304 6294 272504 6354 0 FreeSans 480 0 0 0 spine_iw[17]
port 15 nsew signal input
flabel metal3 s 272304 6158 272504 6218 0 FreeSans 480 0 0 0 spine_iw[18]
port 16 nsew signal input
flabel metal3 s 272304 6022 272504 6082 0 FreeSans 480 0 0 0 spine_iw[19]
port 17 nsew signal input
flabel metal3 s 272304 8470 272504 8530 0 FreeSans 480 0 0 0 spine_iw[1]
port 18 nsew signal input
flabel metal3 s 272304 5886 272504 5946 0 FreeSans 480 0 0 0 spine_iw[20]
port 19 nsew signal input
flabel metal3 s 272304 5750 272504 5810 0 FreeSans 480 0 0 0 spine_iw[21]
port 20 nsew signal input
flabel metal3 s 272304 5614 272504 5674 0 FreeSans 480 0 0 0 spine_iw[22]
port 21 nsew signal input
flabel metal3 s 272304 5478 272504 5538 0 FreeSans 480 0 0 0 spine_iw[23]
port 22 nsew signal input
flabel metal3 s 272304 5342 272504 5402 0 FreeSans 480 0 0 0 spine_iw[24]
port 23 nsew signal input
flabel metal3 s 272304 5206 272504 5266 0 FreeSans 480 0 0 0 spine_iw[25]
port 24 nsew signal input
flabel metal3 s 272304 5070 272504 5130 0 FreeSans 480 0 0 0 spine_iw[26]
port 25 nsew signal input
flabel metal3 s 272304 4934 272504 4994 0 FreeSans 480 0 0 0 spine_iw[27]
port 26 nsew signal input
flabel metal3 s 272304 4798 272504 4858 0 FreeSans 480 0 0 0 spine_iw[28]
port 27 nsew signal input
flabel metal3 s 272304 4662 272504 4722 0 FreeSans 480 0 0 0 spine_iw[29]
port 28 nsew signal input
flabel metal3 s 272304 8334 272504 8394 0 FreeSans 480 0 0 0 spine_iw[2]
port 29 nsew signal input
flabel metal3 s 272304 4526 272504 4586 0 FreeSans 480 0 0 0 spine_iw[30]
port 30 nsew signal input
flabel metal3 s 272304 8198 272504 8258 0 FreeSans 480 0 0 0 spine_iw[3]
port 31 nsew signal input
flabel metal3 s 272304 8062 272504 8122 0 FreeSans 480 0 0 0 spine_iw[4]
port 32 nsew signal input
flabel metal3 s 272304 7926 272504 7986 0 FreeSans 480 0 0 0 spine_iw[5]
port 33 nsew signal input
flabel metal3 s 272304 7790 272504 7850 0 FreeSans 480 0 0 0 spine_iw[6]
port 34 nsew signal input
flabel metal3 s 272304 7654 272504 7714 0 FreeSans 480 0 0 0 spine_iw[7]
port 35 nsew signal input
flabel metal3 s 272304 7518 272504 7578 0 FreeSans 480 0 0 0 spine_iw[8]
port 36 nsew signal input
flabel metal3 s 272304 7382 272504 7442 0 FreeSans 480 0 0 0 spine_iw[9]
port 37 nsew signal input
flabel metal3 s 272304 4390 272504 4450 0 FreeSans 480 0 0 0 spine_ow[0]
port 38 nsew signal tristate
flabel metal3 s 272304 3030 272504 3090 0 FreeSans 480 0 0 0 spine_ow[10]
port 39 nsew signal tristate
flabel metal3 s 272304 2894 272504 2954 0 FreeSans 480 0 0 0 spine_ow[11]
port 40 nsew signal tristate
flabel metal3 s 272304 2758 272504 2818 0 FreeSans 480 0 0 0 spine_ow[12]
port 41 nsew signal tristate
flabel metal3 s 272304 2622 272504 2682 0 FreeSans 480 0 0 0 spine_ow[13]
port 42 nsew signal tristate
flabel metal3 s 272304 2486 272504 2546 0 FreeSans 480 0 0 0 spine_ow[14]
port 43 nsew signal tristate
flabel metal3 s 272304 2350 272504 2410 0 FreeSans 480 0 0 0 spine_ow[15]
port 44 nsew signal tristate
flabel metal3 s 272304 2214 272504 2274 0 FreeSans 480 0 0 0 spine_ow[16]
port 45 nsew signal tristate
flabel metal3 s 272304 2078 272504 2138 0 FreeSans 480 0 0 0 spine_ow[17]
port 46 nsew signal tristate
flabel metal3 s 272304 1942 272504 2002 0 FreeSans 480 0 0 0 spine_ow[18]
port 47 nsew signal tristate
flabel metal3 s 272304 1806 272504 1866 0 FreeSans 480 0 0 0 spine_ow[19]
port 48 nsew signal tristate
flabel metal3 s 272304 4254 272504 4314 0 FreeSans 480 0 0 0 spine_ow[1]
port 49 nsew signal tristate
flabel metal3 s 272304 1670 272504 1730 0 FreeSans 480 0 0 0 spine_ow[20]
port 50 nsew signal tristate
flabel metal3 s 272304 1534 272504 1594 0 FreeSans 480 0 0 0 spine_ow[21]
port 51 nsew signal tristate
flabel metal3 s 272304 1398 272504 1458 0 FreeSans 480 0 0 0 spine_ow[22]
port 52 nsew signal tristate
flabel metal3 s 272304 1262 272504 1322 0 FreeSans 480 0 0 0 spine_ow[23]
port 53 nsew signal tristate
flabel metal3 s 272304 1126 272504 1186 0 FreeSans 480 0 0 0 spine_ow[24]
port 54 nsew signal tristate
flabel metal3 s 272304 990 272504 1050 0 FreeSans 480 0 0 0 spine_ow[25]
port 55 nsew signal tristate
flabel metal3 s 272304 4118 272504 4178 0 FreeSans 480 0 0 0 spine_ow[2]
port 56 nsew signal tristate
flabel metal3 s 272304 3982 272504 4042 0 FreeSans 480 0 0 0 spine_ow[3]
port 57 nsew signal tristate
flabel metal3 s 272304 3846 272504 3906 0 FreeSans 480 0 0 0 spine_ow[4]
port 58 nsew signal tristate
flabel metal3 s 272304 3710 272504 3770 0 FreeSans 480 0 0 0 spine_ow[5]
port 59 nsew signal tristate
flabel metal3 s 272304 3574 272504 3634 0 FreeSans 480 0 0 0 spine_ow[6]
port 60 nsew signal tristate
flabel metal3 s 272304 3438 272504 3498 0 FreeSans 480 0 0 0 spine_ow[7]
port 61 nsew signal tristate
flabel metal3 s 272304 3302 272504 3362 0 FreeSans 480 0 0 0 spine_ow[8]
port 62 nsew signal tristate
flabel metal3 s 272304 3166 272504 3226 0 FreeSans 480 0 0 0 spine_ow[9]
port 63 nsew signal tristate
flabel metal4 s 32446 0 32506 200 0 FreeSans 480 90 0 0 um_ena[0]
port 64 nsew signal tristate
flabel metal4 s 203106 0 203166 200 0 FreeSans 480 90 0 0 um_ena[10]
port 65 nsew signal tristate
flabel metal4 s 203106 10680 203166 10880 0 FreeSans 480 90 0 0 um_ena[11]
port 66 nsew signal tristate
flabel metal4 s 237238 0 237298 200 0 FreeSans 480 90 0 0 um_ena[12]
port 67 nsew signal tristate
flabel metal4 s 237238 10680 237298 10880 0 FreeSans 480 90 0 0 um_ena[13]
port 68 nsew signal tristate
flabel metal4 s 271370 0 271430 200 0 FreeSans 480 90 0 0 um_ena[14]
port 69 nsew signal tristate
flabel metal4 s 271370 10680 271430 10880 0 FreeSans 480 90 0 0 um_ena[15]
port 70 nsew signal tristate
flabel metal4 s 32446 10680 32506 10880 0 FreeSans 480 90 0 0 um_ena[1]
port 71 nsew signal tristate
flabel metal4 s 66578 0 66638 200 0 FreeSans 480 90 0 0 um_ena[2]
port 72 nsew signal tristate
flabel metal4 s 66578 10680 66638 10880 0 FreeSans 480 90 0 0 um_ena[3]
port 73 nsew signal tristate
flabel metal4 s 100710 0 100770 200 0 FreeSans 480 90 0 0 um_ena[4]
port 74 nsew signal tristate
flabel metal4 s 100710 10680 100770 10880 0 FreeSans 480 90 0 0 um_ena[5]
port 75 nsew signal tristate
flabel metal4 s 134842 0 134902 200 0 FreeSans 480 90 0 0 um_ena[6]
port 76 nsew signal tristate
flabel metal4 s 134842 10680 134902 10880 0 FreeSans 480 90 0 0 um_ena[7]
port 77 nsew signal tristate
flabel metal4 s 168974 0 169034 200 0 FreeSans 480 90 0 0 um_ena[8]
port 78 nsew signal tristate
flabel metal4 s 168974 10680 169034 10880 0 FreeSans 480 90 0 0 um_ena[9]
port 79 nsew signal tristate
flabel metal4 s 31710 0 31770 200 0 FreeSans 480 90 0 0 um_iw[0]
port 80 nsew signal tristate
flabel metal4 s 92614 10680 92674 10880 0 FreeSans 480 90 0 0 um_iw[100]
port 81 nsew signal tristate
flabel metal4 s 91878 10680 91938 10880 0 FreeSans 480 90 0 0 um_iw[101]
port 82 nsew signal tristate
flabel metal4 s 91142 10680 91202 10880 0 FreeSans 480 90 0 0 um_iw[102]
port 83 nsew signal tristate
flabel metal4 s 90406 10680 90466 10880 0 FreeSans 480 90 0 0 um_iw[103]
port 84 nsew signal tristate
flabel metal4 s 89670 10680 89730 10880 0 FreeSans 480 90 0 0 um_iw[104]
port 85 nsew signal tristate
flabel metal4 s 88934 10680 88994 10880 0 FreeSans 480 90 0 0 um_iw[105]
port 86 nsew signal tristate
flabel metal4 s 88198 10680 88258 10880 0 FreeSans 480 90 0 0 um_iw[106]
port 87 nsew signal tristate
flabel metal4 s 87462 10680 87522 10880 0 FreeSans 480 90 0 0 um_iw[107]
port 88 nsew signal tristate
flabel metal4 s 134106 0 134166 200 0 FreeSans 480 90 0 0 um_iw[108]
port 89 nsew signal tristate
flabel metal4 s 133370 0 133430 200 0 FreeSans 480 90 0 0 um_iw[109]
port 90 nsew signal tristate
flabel metal4 s 24350 0 24410 200 0 FreeSans 480 90 0 0 um_iw[10]
port 91 nsew signal tristate
flabel metal4 s 132634 0 132694 200 0 FreeSans 480 90 0 0 um_iw[110]
port 92 nsew signal tristate
flabel metal4 s 131898 0 131958 200 0 FreeSans 480 90 0 0 um_iw[111]
port 93 nsew signal tristate
flabel metal4 s 131162 0 131222 200 0 FreeSans 480 90 0 0 um_iw[112]
port 94 nsew signal tristate
flabel metal4 s 130426 0 130486 200 0 FreeSans 480 90 0 0 um_iw[113]
port 95 nsew signal tristate
flabel metal4 s 129690 0 129750 200 0 FreeSans 480 90 0 0 um_iw[114]
port 96 nsew signal tristate
flabel metal4 s 128954 0 129014 200 0 FreeSans 480 90 0 0 um_iw[115]
port 97 nsew signal tristate
flabel metal4 s 128218 0 128278 200 0 FreeSans 480 90 0 0 um_iw[116]
port 98 nsew signal tristate
flabel metal4 s 127482 0 127542 200 0 FreeSans 480 90 0 0 um_iw[117]
port 99 nsew signal tristate
flabel metal4 s 126746 0 126806 200 0 FreeSans 480 90 0 0 um_iw[118]
port 100 nsew signal tristate
flabel metal4 s 126010 0 126070 200 0 FreeSans 480 90 0 0 um_iw[119]
port 101 nsew signal tristate
flabel metal4 s 23614 0 23674 200 0 FreeSans 480 90 0 0 um_iw[11]
port 102 nsew signal tristate
flabel metal4 s 125274 0 125334 200 0 FreeSans 480 90 0 0 um_iw[120]
port 103 nsew signal tristate
flabel metal4 s 124538 0 124598 200 0 FreeSans 480 90 0 0 um_iw[121]
port 104 nsew signal tristate
flabel metal4 s 123802 0 123862 200 0 FreeSans 480 90 0 0 um_iw[122]
port 105 nsew signal tristate
flabel metal4 s 123066 0 123126 200 0 FreeSans 480 90 0 0 um_iw[123]
port 106 nsew signal tristate
flabel metal4 s 122330 0 122390 200 0 FreeSans 480 90 0 0 um_iw[124]
port 107 nsew signal tristate
flabel metal4 s 121594 0 121654 200 0 FreeSans 480 90 0 0 um_iw[125]
port 108 nsew signal tristate
flabel metal4 s 134106 10680 134166 10880 0 FreeSans 480 90 0 0 um_iw[126]
port 109 nsew signal tristate
flabel metal4 s 133370 10680 133430 10880 0 FreeSans 480 90 0 0 um_iw[127]
port 110 nsew signal tristate
flabel metal4 s 132634 10680 132694 10880 0 FreeSans 480 90 0 0 um_iw[128]
port 111 nsew signal tristate
flabel metal4 s 131898 10680 131958 10880 0 FreeSans 480 90 0 0 um_iw[129]
port 112 nsew signal tristate
flabel metal4 s 22878 0 22938 200 0 FreeSans 480 90 0 0 um_iw[12]
port 113 nsew signal tristate
flabel metal4 s 131162 10680 131222 10880 0 FreeSans 480 90 0 0 um_iw[130]
port 114 nsew signal tristate
flabel metal4 s 130426 10680 130486 10880 0 FreeSans 480 90 0 0 um_iw[131]
port 115 nsew signal tristate
flabel metal4 s 129690 10680 129750 10880 0 FreeSans 480 90 0 0 um_iw[132]
port 116 nsew signal tristate
flabel metal4 s 128954 10680 129014 10880 0 FreeSans 480 90 0 0 um_iw[133]
port 117 nsew signal tristate
flabel metal4 s 128218 10680 128278 10880 0 FreeSans 480 90 0 0 um_iw[134]
port 118 nsew signal tristate
flabel metal4 s 127482 10680 127542 10880 0 FreeSans 480 90 0 0 um_iw[135]
port 119 nsew signal tristate
flabel metal4 s 126746 10680 126806 10880 0 FreeSans 480 90 0 0 um_iw[136]
port 120 nsew signal tristate
flabel metal4 s 126010 10680 126070 10880 0 FreeSans 480 90 0 0 um_iw[137]
port 121 nsew signal tristate
flabel metal4 s 125274 10680 125334 10880 0 FreeSans 480 90 0 0 um_iw[138]
port 122 nsew signal tristate
flabel metal4 s 124538 10680 124598 10880 0 FreeSans 480 90 0 0 um_iw[139]
port 123 nsew signal tristate
flabel metal4 s 22142 0 22202 200 0 FreeSans 480 90 0 0 um_iw[13]
port 124 nsew signal tristate
flabel metal4 s 123802 10680 123862 10880 0 FreeSans 480 90 0 0 um_iw[140]
port 125 nsew signal tristate
flabel metal4 s 123066 10680 123126 10880 0 FreeSans 480 90 0 0 um_iw[141]
port 126 nsew signal tristate
flabel metal4 s 122330 10680 122390 10880 0 FreeSans 480 90 0 0 um_iw[142]
port 127 nsew signal tristate
flabel metal4 s 121594 10680 121654 10880 0 FreeSans 480 90 0 0 um_iw[143]
port 128 nsew signal tristate
flabel metal4 s 168238 0 168298 200 0 FreeSans 480 90 0 0 um_iw[144]
port 129 nsew signal tristate
flabel metal4 s 167502 0 167562 200 0 FreeSans 480 90 0 0 um_iw[145]
port 130 nsew signal tristate
flabel metal4 s 166766 0 166826 200 0 FreeSans 480 90 0 0 um_iw[146]
port 131 nsew signal tristate
flabel metal4 s 166030 0 166090 200 0 FreeSans 480 90 0 0 um_iw[147]
port 132 nsew signal tristate
flabel metal4 s 165294 0 165354 200 0 FreeSans 480 90 0 0 um_iw[148]
port 133 nsew signal tristate
flabel metal4 s 164558 0 164618 200 0 FreeSans 480 90 0 0 um_iw[149]
port 134 nsew signal tristate
flabel metal4 s 21406 0 21466 200 0 FreeSans 480 90 0 0 um_iw[14]
port 135 nsew signal tristate
flabel metal4 s 163822 0 163882 200 0 FreeSans 480 90 0 0 um_iw[150]
port 136 nsew signal tristate
flabel metal4 s 163086 0 163146 200 0 FreeSans 480 90 0 0 um_iw[151]
port 137 nsew signal tristate
flabel metal4 s 162350 0 162410 200 0 FreeSans 480 90 0 0 um_iw[152]
port 138 nsew signal tristate
flabel metal4 s 161614 0 161674 200 0 FreeSans 480 90 0 0 um_iw[153]
port 139 nsew signal tristate
flabel metal4 s 160878 0 160938 200 0 FreeSans 480 90 0 0 um_iw[154]
port 140 nsew signal tristate
flabel metal4 s 160142 0 160202 200 0 FreeSans 480 90 0 0 um_iw[155]
port 141 nsew signal tristate
flabel metal4 s 159406 0 159466 200 0 FreeSans 480 90 0 0 um_iw[156]
port 142 nsew signal tristate
flabel metal4 s 158670 0 158730 200 0 FreeSans 480 90 0 0 um_iw[157]
port 143 nsew signal tristate
flabel metal4 s 157934 0 157994 200 0 FreeSans 480 90 0 0 um_iw[158]
port 144 nsew signal tristate
flabel metal4 s 157198 0 157258 200 0 FreeSans 480 90 0 0 um_iw[159]
port 145 nsew signal tristate
flabel metal4 s 20670 0 20730 200 0 FreeSans 480 90 0 0 um_iw[15]
port 146 nsew signal tristate
flabel metal4 s 156462 0 156522 200 0 FreeSans 480 90 0 0 um_iw[160]
port 147 nsew signal tristate
flabel metal4 s 155726 0 155786 200 0 FreeSans 480 90 0 0 um_iw[161]
port 148 nsew signal tristate
flabel metal4 s 168238 10680 168298 10880 0 FreeSans 480 90 0 0 um_iw[162]
port 149 nsew signal tristate
flabel metal4 s 167502 10680 167562 10880 0 FreeSans 480 90 0 0 um_iw[163]
port 150 nsew signal tristate
flabel metal4 s 166766 10680 166826 10880 0 FreeSans 480 90 0 0 um_iw[164]
port 151 nsew signal tristate
flabel metal4 s 166030 10680 166090 10880 0 FreeSans 480 90 0 0 um_iw[165]
port 152 nsew signal tristate
flabel metal4 s 165294 10680 165354 10880 0 FreeSans 480 90 0 0 um_iw[166]
port 153 nsew signal tristate
flabel metal4 s 164558 10680 164618 10880 0 FreeSans 480 90 0 0 um_iw[167]
port 154 nsew signal tristate
flabel metal4 s 163822 10680 163882 10880 0 FreeSans 480 90 0 0 um_iw[168]
port 155 nsew signal tristate
flabel metal4 s 163086 10680 163146 10880 0 FreeSans 480 90 0 0 um_iw[169]
port 156 nsew signal tristate
flabel metal4 s 19934 0 19994 200 0 FreeSans 480 90 0 0 um_iw[16]
port 157 nsew signal tristate
flabel metal4 s 162350 10680 162410 10880 0 FreeSans 480 90 0 0 um_iw[170]
port 158 nsew signal tristate
flabel metal4 s 161614 10680 161674 10880 0 FreeSans 480 90 0 0 um_iw[171]
port 159 nsew signal tristate
flabel metal4 s 160878 10680 160938 10880 0 FreeSans 480 90 0 0 um_iw[172]
port 160 nsew signal tristate
flabel metal4 s 160142 10680 160202 10880 0 FreeSans 480 90 0 0 um_iw[173]
port 161 nsew signal tristate
flabel metal4 s 159406 10680 159466 10880 0 FreeSans 480 90 0 0 um_iw[174]
port 162 nsew signal tristate
flabel metal4 s 158670 10680 158730 10880 0 FreeSans 480 90 0 0 um_iw[175]
port 163 nsew signal tristate
flabel metal4 s 157934 10680 157994 10880 0 FreeSans 480 90 0 0 um_iw[176]
port 164 nsew signal tristate
flabel metal4 s 157198 10680 157258 10880 0 FreeSans 480 90 0 0 um_iw[177]
port 165 nsew signal tristate
flabel metal4 s 156462 10680 156522 10880 0 FreeSans 480 90 0 0 um_iw[178]
port 166 nsew signal tristate
flabel metal4 s 155726 10680 155786 10880 0 FreeSans 480 90 0 0 um_iw[179]
port 167 nsew signal tristate
flabel metal4 s 19198 0 19258 200 0 FreeSans 480 90 0 0 um_iw[17]
port 168 nsew signal tristate
flabel metal4 s 202370 0 202430 200 0 FreeSans 480 90 0 0 um_iw[180]
port 169 nsew signal tristate
flabel metal4 s 201634 0 201694 200 0 FreeSans 480 90 0 0 um_iw[181]
port 170 nsew signal tristate
flabel metal4 s 200898 0 200958 200 0 FreeSans 480 90 0 0 um_iw[182]
port 171 nsew signal tristate
flabel metal4 s 200162 0 200222 200 0 FreeSans 480 90 0 0 um_iw[183]
port 172 nsew signal tristate
flabel metal4 s 199426 0 199486 200 0 FreeSans 480 90 0 0 um_iw[184]
port 173 nsew signal tristate
flabel metal4 s 198690 0 198750 200 0 FreeSans 480 90 0 0 um_iw[185]
port 174 nsew signal tristate
flabel metal4 s 197954 0 198014 200 0 FreeSans 480 90 0 0 um_iw[186]
port 175 nsew signal tristate
flabel metal4 s 197218 0 197278 200 0 FreeSans 480 90 0 0 um_iw[187]
port 176 nsew signal tristate
flabel metal4 s 196482 0 196542 200 0 FreeSans 480 90 0 0 um_iw[188]
port 177 nsew signal tristate
flabel metal4 s 195746 0 195806 200 0 FreeSans 480 90 0 0 um_iw[189]
port 178 nsew signal tristate
flabel metal4 s 31710 10680 31770 10880 0 FreeSans 480 90 0 0 um_iw[18]
port 179 nsew signal tristate
flabel metal4 s 195010 0 195070 200 0 FreeSans 480 90 0 0 um_iw[190]
port 180 nsew signal tristate
flabel metal4 s 194274 0 194334 200 0 FreeSans 480 90 0 0 um_iw[191]
port 181 nsew signal tristate
flabel metal4 s 193538 0 193598 200 0 FreeSans 480 90 0 0 um_iw[192]
port 182 nsew signal tristate
flabel metal4 s 192802 0 192862 200 0 FreeSans 480 90 0 0 um_iw[193]
port 183 nsew signal tristate
flabel metal4 s 192066 0 192126 200 0 FreeSans 480 90 0 0 um_iw[194]
port 184 nsew signal tristate
flabel metal4 s 191330 0 191390 200 0 FreeSans 480 90 0 0 um_iw[195]
port 185 nsew signal tristate
flabel metal4 s 190594 0 190654 200 0 FreeSans 480 90 0 0 um_iw[196]
port 186 nsew signal tristate
flabel metal4 s 189858 0 189918 200 0 FreeSans 480 90 0 0 um_iw[197]
port 187 nsew signal tristate
flabel metal4 s 202370 10680 202430 10880 0 FreeSans 480 90 0 0 um_iw[198]
port 188 nsew signal tristate
flabel metal4 s 201634 10680 201694 10880 0 FreeSans 480 90 0 0 um_iw[199]
port 189 nsew signal tristate
flabel metal4 s 30974 10680 31034 10880 0 FreeSans 480 90 0 0 um_iw[19]
port 190 nsew signal tristate
flabel metal4 s 30974 0 31034 200 0 FreeSans 480 90 0 0 um_iw[1]
port 191 nsew signal tristate
flabel metal4 s 200898 10680 200958 10880 0 FreeSans 480 90 0 0 um_iw[200]
port 192 nsew signal tristate
flabel metal4 s 200162 10680 200222 10880 0 FreeSans 480 90 0 0 um_iw[201]
port 193 nsew signal tristate
flabel metal4 s 199426 10680 199486 10880 0 FreeSans 480 90 0 0 um_iw[202]
port 194 nsew signal tristate
flabel metal4 s 198690 10680 198750 10880 0 FreeSans 480 90 0 0 um_iw[203]
port 195 nsew signal tristate
flabel metal4 s 197954 10680 198014 10880 0 FreeSans 480 90 0 0 um_iw[204]
port 196 nsew signal tristate
flabel metal4 s 197218 10680 197278 10880 0 FreeSans 480 90 0 0 um_iw[205]
port 197 nsew signal tristate
flabel metal4 s 196482 10680 196542 10880 0 FreeSans 480 90 0 0 um_iw[206]
port 198 nsew signal tristate
flabel metal4 s 195746 10680 195806 10880 0 FreeSans 480 90 0 0 um_iw[207]
port 199 nsew signal tristate
flabel metal4 s 195010 10680 195070 10880 0 FreeSans 480 90 0 0 um_iw[208]
port 200 nsew signal tristate
flabel metal4 s 194274 10680 194334 10880 0 FreeSans 480 90 0 0 um_iw[209]
port 201 nsew signal tristate
flabel metal4 s 30238 10680 30298 10880 0 FreeSans 480 90 0 0 um_iw[20]
port 202 nsew signal tristate
flabel metal4 s 193538 10680 193598 10880 0 FreeSans 480 90 0 0 um_iw[210]
port 203 nsew signal tristate
flabel metal4 s 192802 10680 192862 10880 0 FreeSans 480 90 0 0 um_iw[211]
port 204 nsew signal tristate
flabel metal4 s 192066 10680 192126 10880 0 FreeSans 480 90 0 0 um_iw[212]
port 205 nsew signal tristate
flabel metal4 s 191330 10680 191390 10880 0 FreeSans 480 90 0 0 um_iw[213]
port 206 nsew signal tristate
flabel metal4 s 190594 10680 190654 10880 0 FreeSans 480 90 0 0 um_iw[214]
port 207 nsew signal tristate
flabel metal4 s 189858 10680 189918 10880 0 FreeSans 480 90 0 0 um_iw[215]
port 208 nsew signal tristate
flabel metal4 s 236502 0 236562 200 0 FreeSans 480 90 0 0 um_iw[216]
port 209 nsew signal tristate
flabel metal4 s 235766 0 235826 200 0 FreeSans 480 90 0 0 um_iw[217]
port 210 nsew signal tristate
flabel metal4 s 235030 0 235090 200 0 FreeSans 480 90 0 0 um_iw[218]
port 211 nsew signal tristate
flabel metal4 s 234294 0 234354 200 0 FreeSans 480 90 0 0 um_iw[219]
port 212 nsew signal tristate
flabel metal4 s 29502 10680 29562 10880 0 FreeSans 480 90 0 0 um_iw[21]
port 213 nsew signal tristate
flabel metal4 s 233558 0 233618 200 0 FreeSans 480 90 0 0 um_iw[220]
port 214 nsew signal tristate
flabel metal4 s 232822 0 232882 200 0 FreeSans 480 90 0 0 um_iw[221]
port 215 nsew signal tristate
flabel metal4 s 232086 0 232146 200 0 FreeSans 480 90 0 0 um_iw[222]
port 216 nsew signal tristate
flabel metal4 s 231350 0 231410 200 0 FreeSans 480 90 0 0 um_iw[223]
port 217 nsew signal tristate
flabel metal4 s 230614 0 230674 200 0 FreeSans 480 90 0 0 um_iw[224]
port 218 nsew signal tristate
flabel metal4 s 229878 0 229938 200 0 FreeSans 480 90 0 0 um_iw[225]
port 219 nsew signal tristate
flabel metal4 s 229142 0 229202 200 0 FreeSans 480 90 0 0 um_iw[226]
port 220 nsew signal tristate
flabel metal4 s 228406 0 228466 200 0 FreeSans 480 90 0 0 um_iw[227]
port 221 nsew signal tristate
flabel metal4 s 227670 0 227730 200 0 FreeSans 480 90 0 0 um_iw[228]
port 222 nsew signal tristate
flabel metal4 s 226934 0 226994 200 0 FreeSans 480 90 0 0 um_iw[229]
port 223 nsew signal tristate
flabel metal4 s 28766 10680 28826 10880 0 FreeSans 480 90 0 0 um_iw[22]
port 224 nsew signal tristate
flabel metal4 s 226198 0 226258 200 0 FreeSans 480 90 0 0 um_iw[230]
port 225 nsew signal tristate
flabel metal4 s 225462 0 225522 200 0 FreeSans 480 90 0 0 um_iw[231]
port 226 nsew signal tristate
flabel metal4 s 224726 0 224786 200 0 FreeSans 480 90 0 0 um_iw[232]
port 227 nsew signal tristate
flabel metal4 s 223990 0 224050 200 0 FreeSans 480 90 0 0 um_iw[233]
port 228 nsew signal tristate
flabel metal4 s 236502 10680 236562 10880 0 FreeSans 480 90 0 0 um_iw[234]
port 229 nsew signal tristate
flabel metal4 s 235766 10680 235826 10880 0 FreeSans 480 90 0 0 um_iw[235]
port 230 nsew signal tristate
flabel metal4 s 235030 10680 235090 10880 0 FreeSans 480 90 0 0 um_iw[236]
port 231 nsew signal tristate
flabel metal4 s 234294 10680 234354 10880 0 FreeSans 480 90 0 0 um_iw[237]
port 232 nsew signal tristate
flabel metal4 s 233558 10680 233618 10880 0 FreeSans 480 90 0 0 um_iw[238]
port 233 nsew signal tristate
flabel metal4 s 232822 10680 232882 10880 0 FreeSans 480 90 0 0 um_iw[239]
port 234 nsew signal tristate
flabel metal4 s 28030 10680 28090 10880 0 FreeSans 480 90 0 0 um_iw[23]
port 235 nsew signal tristate
flabel metal4 s 232086 10680 232146 10880 0 FreeSans 480 90 0 0 um_iw[240]
port 236 nsew signal tristate
flabel metal4 s 231350 10680 231410 10880 0 FreeSans 480 90 0 0 um_iw[241]
port 237 nsew signal tristate
flabel metal4 s 230614 10680 230674 10880 0 FreeSans 480 90 0 0 um_iw[242]
port 238 nsew signal tristate
flabel metal4 s 229878 10680 229938 10880 0 FreeSans 480 90 0 0 um_iw[243]
port 239 nsew signal tristate
flabel metal4 s 229142 10680 229202 10880 0 FreeSans 480 90 0 0 um_iw[244]
port 240 nsew signal tristate
flabel metal4 s 228406 10680 228466 10880 0 FreeSans 480 90 0 0 um_iw[245]
port 241 nsew signal tristate
flabel metal4 s 227670 10680 227730 10880 0 FreeSans 480 90 0 0 um_iw[246]
port 242 nsew signal tristate
flabel metal4 s 226934 10680 226994 10880 0 FreeSans 480 90 0 0 um_iw[247]
port 243 nsew signal tristate
flabel metal4 s 226198 10680 226258 10880 0 FreeSans 480 90 0 0 um_iw[248]
port 244 nsew signal tristate
flabel metal4 s 225462 10680 225522 10880 0 FreeSans 480 90 0 0 um_iw[249]
port 245 nsew signal tristate
flabel metal4 s 27294 10680 27354 10880 0 FreeSans 480 90 0 0 um_iw[24]
port 246 nsew signal tristate
flabel metal4 s 224726 10680 224786 10880 0 FreeSans 480 90 0 0 um_iw[250]
port 247 nsew signal tristate
flabel metal4 s 223990 10680 224050 10880 0 FreeSans 480 90 0 0 um_iw[251]
port 248 nsew signal tristate
flabel metal4 s 270634 0 270694 200 0 FreeSans 480 90 0 0 um_iw[252]
port 249 nsew signal tristate
flabel metal4 s 269898 0 269958 200 0 FreeSans 480 90 0 0 um_iw[253]
port 250 nsew signal tristate
flabel metal4 s 269162 0 269222 200 0 FreeSans 480 90 0 0 um_iw[254]
port 251 nsew signal tristate
flabel metal4 s 268426 0 268486 200 0 FreeSans 480 90 0 0 um_iw[255]
port 252 nsew signal tristate
flabel metal4 s 267690 0 267750 200 0 FreeSans 480 90 0 0 um_iw[256]
port 253 nsew signal tristate
flabel metal4 s 266954 0 267014 200 0 FreeSans 480 90 0 0 um_iw[257]
port 254 nsew signal tristate
flabel metal4 s 266218 0 266278 200 0 FreeSans 480 90 0 0 um_iw[258]
port 255 nsew signal tristate
flabel metal4 s 265482 0 265542 200 0 FreeSans 480 90 0 0 um_iw[259]
port 256 nsew signal tristate
flabel metal4 s 26558 10680 26618 10880 0 FreeSans 480 90 0 0 um_iw[25]
port 257 nsew signal tristate
flabel metal4 s 264746 0 264806 200 0 FreeSans 480 90 0 0 um_iw[260]
port 258 nsew signal tristate
flabel metal4 s 264010 0 264070 200 0 FreeSans 480 90 0 0 um_iw[261]
port 259 nsew signal tristate
flabel metal4 s 263274 0 263334 200 0 FreeSans 480 90 0 0 um_iw[262]
port 260 nsew signal tristate
flabel metal4 s 262538 0 262598 200 0 FreeSans 480 90 0 0 um_iw[263]
port 261 nsew signal tristate
flabel metal4 s 261802 0 261862 200 0 FreeSans 480 90 0 0 um_iw[264]
port 262 nsew signal tristate
flabel metal4 s 261066 0 261126 200 0 FreeSans 480 90 0 0 um_iw[265]
port 263 nsew signal tristate
flabel metal4 s 260330 0 260390 200 0 FreeSans 480 90 0 0 um_iw[266]
port 264 nsew signal tristate
flabel metal4 s 259594 0 259654 200 0 FreeSans 480 90 0 0 um_iw[267]
port 265 nsew signal tristate
flabel metal4 s 258858 0 258918 200 0 FreeSans 480 90 0 0 um_iw[268]
port 266 nsew signal tristate
flabel metal4 s 258122 0 258182 200 0 FreeSans 480 90 0 0 um_iw[269]
port 267 nsew signal tristate
flabel metal4 s 25822 10680 25882 10880 0 FreeSans 480 90 0 0 um_iw[26]
port 268 nsew signal tristate
flabel metal4 s 270634 10680 270694 10880 0 FreeSans 480 90 0 0 um_iw[270]
port 269 nsew signal tristate
flabel metal4 s 269898 10680 269958 10880 0 FreeSans 480 90 0 0 um_iw[271]
port 270 nsew signal tristate
flabel metal4 s 269162 10680 269222 10880 0 FreeSans 480 90 0 0 um_iw[272]
port 271 nsew signal tristate
flabel metal4 s 268426 10680 268486 10880 0 FreeSans 480 90 0 0 um_iw[273]
port 272 nsew signal tristate
flabel metal4 s 267690 10680 267750 10880 0 FreeSans 480 90 0 0 um_iw[274]
port 273 nsew signal tristate
flabel metal4 s 266954 10680 267014 10880 0 FreeSans 480 90 0 0 um_iw[275]
port 274 nsew signal tristate
flabel metal4 s 266218 10680 266278 10880 0 FreeSans 480 90 0 0 um_iw[276]
port 275 nsew signal tristate
flabel metal4 s 265482 10680 265542 10880 0 FreeSans 480 90 0 0 um_iw[277]
port 276 nsew signal tristate
flabel metal4 s 264746 10680 264806 10880 0 FreeSans 480 90 0 0 um_iw[278]
port 277 nsew signal tristate
flabel metal4 s 264010 10680 264070 10880 0 FreeSans 480 90 0 0 um_iw[279]
port 278 nsew signal tristate
flabel metal4 s 25086 10680 25146 10880 0 FreeSans 480 90 0 0 um_iw[27]
port 279 nsew signal tristate
flabel metal4 s 263274 10680 263334 10880 0 FreeSans 480 90 0 0 um_iw[280]
port 280 nsew signal tristate
flabel metal4 s 262538 10680 262598 10880 0 FreeSans 480 90 0 0 um_iw[281]
port 281 nsew signal tristate
flabel metal4 s 261802 10680 261862 10880 0 FreeSans 480 90 0 0 um_iw[282]
port 282 nsew signal tristate
flabel metal4 s 261066 10680 261126 10880 0 FreeSans 480 90 0 0 um_iw[283]
port 283 nsew signal tristate
flabel metal4 s 260330 10680 260390 10880 0 FreeSans 480 90 0 0 um_iw[284]
port 284 nsew signal tristate
flabel metal4 s 259594 10680 259654 10880 0 FreeSans 480 90 0 0 um_iw[285]
port 285 nsew signal tristate
flabel metal4 s 258858 10680 258918 10880 0 FreeSans 480 90 0 0 um_iw[286]
port 286 nsew signal tristate
flabel metal4 s 258122 10680 258182 10880 0 FreeSans 480 90 0 0 um_iw[287]
port 287 nsew signal tristate
flabel metal4 s 24350 10680 24410 10880 0 FreeSans 480 90 0 0 um_iw[28]
port 288 nsew signal tristate
flabel metal4 s 23614 10680 23674 10880 0 FreeSans 480 90 0 0 um_iw[29]
port 289 nsew signal tristate
flabel metal4 s 30238 0 30298 200 0 FreeSans 480 90 0 0 um_iw[2]
port 290 nsew signal tristate
flabel metal4 s 22878 10680 22938 10880 0 FreeSans 480 90 0 0 um_iw[30]
port 291 nsew signal tristate
flabel metal4 s 22142 10680 22202 10880 0 FreeSans 480 90 0 0 um_iw[31]
port 292 nsew signal tristate
flabel metal4 s 21406 10680 21466 10880 0 FreeSans 480 90 0 0 um_iw[32]
port 293 nsew signal tristate
flabel metal4 s 20670 10680 20730 10880 0 FreeSans 480 90 0 0 um_iw[33]
port 294 nsew signal tristate
flabel metal4 s 19934 10680 19994 10880 0 FreeSans 480 90 0 0 um_iw[34]
port 295 nsew signal tristate
flabel metal4 s 19198 10680 19258 10880 0 FreeSans 480 90 0 0 um_iw[35]
port 296 nsew signal tristate
flabel metal4 s 65842 0 65902 200 0 FreeSans 480 90 0 0 um_iw[36]
port 297 nsew signal tristate
flabel metal4 s 65106 0 65166 200 0 FreeSans 480 90 0 0 um_iw[37]
port 298 nsew signal tristate
flabel metal4 s 64370 0 64430 200 0 FreeSans 480 90 0 0 um_iw[38]
port 299 nsew signal tristate
flabel metal4 s 63634 0 63694 200 0 FreeSans 480 90 0 0 um_iw[39]
port 300 nsew signal tristate
flabel metal4 s 29502 0 29562 200 0 FreeSans 480 90 0 0 um_iw[3]
port 301 nsew signal tristate
flabel metal4 s 62898 0 62958 200 0 FreeSans 480 90 0 0 um_iw[40]
port 302 nsew signal tristate
flabel metal4 s 62162 0 62222 200 0 FreeSans 480 90 0 0 um_iw[41]
port 303 nsew signal tristate
flabel metal4 s 61426 0 61486 200 0 FreeSans 480 90 0 0 um_iw[42]
port 304 nsew signal tristate
flabel metal4 s 60690 0 60750 200 0 FreeSans 480 90 0 0 um_iw[43]
port 305 nsew signal tristate
flabel metal4 s 59954 0 60014 200 0 FreeSans 480 90 0 0 um_iw[44]
port 306 nsew signal tristate
flabel metal4 s 59218 0 59278 200 0 FreeSans 480 90 0 0 um_iw[45]
port 307 nsew signal tristate
flabel metal4 s 58482 0 58542 200 0 FreeSans 480 90 0 0 um_iw[46]
port 308 nsew signal tristate
flabel metal4 s 57746 0 57806 200 0 FreeSans 480 90 0 0 um_iw[47]
port 309 nsew signal tristate
flabel metal4 s 57010 0 57070 200 0 FreeSans 480 90 0 0 um_iw[48]
port 310 nsew signal tristate
flabel metal4 s 56274 0 56334 200 0 FreeSans 480 90 0 0 um_iw[49]
port 311 nsew signal tristate
flabel metal4 s 28766 0 28826 200 0 FreeSans 480 90 0 0 um_iw[4]
port 312 nsew signal tristate
flabel metal4 s 55538 0 55598 200 0 FreeSans 480 90 0 0 um_iw[50]
port 313 nsew signal tristate
flabel metal4 s 54802 0 54862 200 0 FreeSans 480 90 0 0 um_iw[51]
port 314 nsew signal tristate
flabel metal4 s 54066 0 54126 200 0 FreeSans 480 90 0 0 um_iw[52]
port 315 nsew signal tristate
flabel metal4 s 53330 0 53390 200 0 FreeSans 480 90 0 0 um_iw[53]
port 316 nsew signal tristate
flabel metal4 s 65842 10680 65902 10880 0 FreeSans 480 90 0 0 um_iw[54]
port 317 nsew signal tristate
flabel metal4 s 65106 10680 65166 10880 0 FreeSans 480 90 0 0 um_iw[55]
port 318 nsew signal tristate
flabel metal4 s 64370 10680 64430 10880 0 FreeSans 480 90 0 0 um_iw[56]
port 319 nsew signal tristate
flabel metal4 s 63634 10680 63694 10880 0 FreeSans 480 90 0 0 um_iw[57]
port 320 nsew signal tristate
flabel metal4 s 62898 10680 62958 10880 0 FreeSans 480 90 0 0 um_iw[58]
port 321 nsew signal tristate
flabel metal4 s 62162 10680 62222 10880 0 FreeSans 480 90 0 0 um_iw[59]
port 322 nsew signal tristate
flabel metal4 s 28030 0 28090 200 0 FreeSans 480 90 0 0 um_iw[5]
port 323 nsew signal tristate
flabel metal4 s 61426 10680 61486 10880 0 FreeSans 480 90 0 0 um_iw[60]
port 324 nsew signal tristate
flabel metal4 s 60690 10680 60750 10880 0 FreeSans 480 90 0 0 um_iw[61]
port 325 nsew signal tristate
flabel metal4 s 59954 10680 60014 10880 0 FreeSans 480 90 0 0 um_iw[62]
port 326 nsew signal tristate
flabel metal4 s 59218 10680 59278 10880 0 FreeSans 480 90 0 0 um_iw[63]
port 327 nsew signal tristate
flabel metal4 s 58482 10680 58542 10880 0 FreeSans 480 90 0 0 um_iw[64]
port 328 nsew signal tristate
flabel metal4 s 57746 10680 57806 10880 0 FreeSans 480 90 0 0 um_iw[65]
port 329 nsew signal tristate
flabel metal4 s 57010 10680 57070 10880 0 FreeSans 480 90 0 0 um_iw[66]
port 330 nsew signal tristate
flabel metal4 s 56274 10680 56334 10880 0 FreeSans 480 90 0 0 um_iw[67]
port 331 nsew signal tristate
flabel metal4 s 55538 10680 55598 10880 0 FreeSans 480 90 0 0 um_iw[68]
port 332 nsew signal tristate
flabel metal4 s 54802 10680 54862 10880 0 FreeSans 480 90 0 0 um_iw[69]
port 333 nsew signal tristate
flabel metal4 s 27294 0 27354 200 0 FreeSans 480 90 0 0 um_iw[6]
port 334 nsew signal tristate
flabel metal4 s 54066 10680 54126 10880 0 FreeSans 480 90 0 0 um_iw[70]
port 335 nsew signal tristate
flabel metal4 s 53330 10680 53390 10880 0 FreeSans 480 90 0 0 um_iw[71]
port 336 nsew signal tristate
flabel metal4 s 99974 0 100034 200 0 FreeSans 480 90 0 0 um_iw[72]
port 337 nsew signal tristate
flabel metal4 s 99238 0 99298 200 0 FreeSans 480 90 0 0 um_iw[73]
port 338 nsew signal tristate
flabel metal4 s 98502 0 98562 200 0 FreeSans 480 90 0 0 um_iw[74]
port 339 nsew signal tristate
flabel metal4 s 97766 0 97826 200 0 FreeSans 480 90 0 0 um_iw[75]
port 340 nsew signal tristate
flabel metal4 s 97030 0 97090 200 0 FreeSans 480 90 0 0 um_iw[76]
port 341 nsew signal tristate
flabel metal4 s 96294 0 96354 200 0 FreeSans 480 90 0 0 um_iw[77]
port 342 nsew signal tristate
flabel metal4 s 95558 0 95618 200 0 FreeSans 480 90 0 0 um_iw[78]
port 343 nsew signal tristate
flabel metal4 s 94822 0 94882 200 0 FreeSans 480 90 0 0 um_iw[79]
port 344 nsew signal tristate
flabel metal4 s 26558 0 26618 200 0 FreeSans 480 90 0 0 um_iw[7]
port 345 nsew signal tristate
flabel metal4 s 94086 0 94146 200 0 FreeSans 480 90 0 0 um_iw[80]
port 346 nsew signal tristate
flabel metal4 s 93350 0 93410 200 0 FreeSans 480 90 0 0 um_iw[81]
port 347 nsew signal tristate
flabel metal4 s 92614 0 92674 200 0 FreeSans 480 90 0 0 um_iw[82]
port 348 nsew signal tristate
flabel metal4 s 91878 0 91938 200 0 FreeSans 480 90 0 0 um_iw[83]
port 349 nsew signal tristate
flabel metal4 s 91142 0 91202 200 0 FreeSans 480 90 0 0 um_iw[84]
port 350 nsew signal tristate
flabel metal4 s 90406 0 90466 200 0 FreeSans 480 90 0 0 um_iw[85]
port 351 nsew signal tristate
flabel metal4 s 89670 0 89730 200 0 FreeSans 480 90 0 0 um_iw[86]
port 352 nsew signal tristate
flabel metal4 s 88934 0 88994 200 0 FreeSans 480 90 0 0 um_iw[87]
port 353 nsew signal tristate
flabel metal4 s 88198 0 88258 200 0 FreeSans 480 90 0 0 um_iw[88]
port 354 nsew signal tristate
flabel metal4 s 87462 0 87522 200 0 FreeSans 480 90 0 0 um_iw[89]
port 355 nsew signal tristate
flabel metal4 s 25822 0 25882 200 0 FreeSans 480 90 0 0 um_iw[8]
port 356 nsew signal tristate
flabel metal4 s 99974 10680 100034 10880 0 FreeSans 480 90 0 0 um_iw[90]
port 357 nsew signal tristate
flabel metal4 s 99238 10680 99298 10880 0 FreeSans 480 90 0 0 um_iw[91]
port 358 nsew signal tristate
flabel metal4 s 98502 10680 98562 10880 0 FreeSans 480 90 0 0 um_iw[92]
port 359 nsew signal tristate
flabel metal4 s 97766 10680 97826 10880 0 FreeSans 480 90 0 0 um_iw[93]
port 360 nsew signal tristate
flabel metal4 s 97030 10680 97090 10880 0 FreeSans 480 90 0 0 um_iw[94]
port 361 nsew signal tristate
flabel metal4 s 96294 10680 96354 10880 0 FreeSans 480 90 0 0 um_iw[95]
port 362 nsew signal tristate
flabel metal4 s 95558 10680 95618 10880 0 FreeSans 480 90 0 0 um_iw[96]
port 363 nsew signal tristate
flabel metal4 s 94822 10680 94882 10880 0 FreeSans 480 90 0 0 um_iw[97]
port 364 nsew signal tristate
flabel metal4 s 94086 10680 94146 10880 0 FreeSans 480 90 0 0 um_iw[98]
port 365 nsew signal tristate
flabel metal4 s 93350 10680 93410 10880 0 FreeSans 480 90 0 0 um_iw[99]
port 366 nsew signal tristate
flabel metal4 s 25086 0 25146 200 0 FreeSans 480 90 0 0 um_iw[9]
port 367 nsew signal tristate
flabel metal4 s 798 0 858 200 0 FreeSans 480 90 0 0 um_k_zero[0]
port 368 nsew signal tristate
flabel metal4 s 171458 0 171518 200 0 FreeSans 480 90 0 0 um_k_zero[10]
port 369 nsew signal tristate
flabel metal4 s 171458 10680 171518 10880 0 FreeSans 480 90 0 0 um_k_zero[11]
port 370 nsew signal tristate
flabel metal4 s 205590 0 205650 200 0 FreeSans 480 90 0 0 um_k_zero[12]
port 371 nsew signal tristate
flabel metal4 s 205590 10680 205650 10880 0 FreeSans 480 90 0 0 um_k_zero[13]
port 372 nsew signal tristate
flabel metal4 s 239722 0 239782 200 0 FreeSans 480 90 0 0 um_k_zero[14]
port 373 nsew signal tristate
flabel metal4 s 239722 10680 239782 10880 0 FreeSans 480 90 0 0 um_k_zero[15]
port 374 nsew signal tristate
flabel metal4 s 798 10680 858 10880 0 FreeSans 480 90 0 0 um_k_zero[1]
port 375 nsew signal tristate
flabel metal4 s 34930 0 34990 200 0 FreeSans 480 90 0 0 um_k_zero[2]
port 376 nsew signal tristate
flabel metal4 s 34930 10680 34990 10880 0 FreeSans 480 90 0 0 um_k_zero[3]
port 377 nsew signal tristate
flabel metal4 s 69062 0 69122 200 0 FreeSans 480 90 0 0 um_k_zero[4]
port 378 nsew signal tristate
flabel metal4 s 69062 10680 69122 10880 0 FreeSans 480 90 0 0 um_k_zero[5]
port 379 nsew signal tristate
flabel metal4 s 103194 0 103254 200 0 FreeSans 480 90 0 0 um_k_zero[6]
port 380 nsew signal tristate
flabel metal4 s 103194 10680 103254 10880 0 FreeSans 480 90 0 0 um_k_zero[7]
port 381 nsew signal tristate
flabel metal4 s 137326 0 137386 200 0 FreeSans 480 90 0 0 um_k_zero[8]
port 382 nsew signal tristate
flabel metal4 s 137326 10680 137386 10880 0 FreeSans 480 90 0 0 um_k_zero[9]
port 383 nsew signal tristate
flabel metal4 s 18462 0 18522 200 0 FreeSans 480 90 0 0 um_ow[0]
port 384 nsew signal input
flabel metal4 s 83782 0 83842 200 0 FreeSans 480 90 0 0 um_ow[100]
port 385 nsew signal input
flabel metal4 s 83046 0 83106 200 0 FreeSans 480 90 0 0 um_ow[101]
port 386 nsew signal input
flabel metal4 s 82310 0 82370 200 0 FreeSans 480 90 0 0 um_ow[102]
port 387 nsew signal input
flabel metal4 s 81574 0 81634 200 0 FreeSans 480 90 0 0 um_ow[103]
port 388 nsew signal input
flabel metal4 s 80838 0 80898 200 0 FreeSans 480 90 0 0 um_ow[104]
port 389 nsew signal input
flabel metal4 s 80102 0 80162 200 0 FreeSans 480 90 0 0 um_ow[105]
port 390 nsew signal input
flabel metal4 s 79366 0 79426 200 0 FreeSans 480 90 0 0 um_ow[106]
port 391 nsew signal input
flabel metal4 s 78630 0 78690 200 0 FreeSans 480 90 0 0 um_ow[107]
port 392 nsew signal input
flabel metal4 s 77894 0 77954 200 0 FreeSans 480 90 0 0 um_ow[108]
port 393 nsew signal input
flabel metal4 s 77158 0 77218 200 0 FreeSans 480 90 0 0 um_ow[109]
port 394 nsew signal input
flabel metal4 s 11102 0 11162 200 0 FreeSans 480 90 0 0 um_ow[10]
port 395 nsew signal input
flabel metal4 s 76422 0 76482 200 0 FreeSans 480 90 0 0 um_ow[110]
port 396 nsew signal input
flabel metal4 s 75686 0 75746 200 0 FreeSans 480 90 0 0 um_ow[111]
port 397 nsew signal input
flabel metal4 s 74950 0 75010 200 0 FreeSans 480 90 0 0 um_ow[112]
port 398 nsew signal input
flabel metal4 s 74214 0 74274 200 0 FreeSans 480 90 0 0 um_ow[113]
port 399 nsew signal input
flabel metal4 s 73478 0 73538 200 0 FreeSans 480 90 0 0 um_ow[114]
port 400 nsew signal input
flabel metal4 s 72742 0 72802 200 0 FreeSans 480 90 0 0 um_ow[115]
port 401 nsew signal input
flabel metal4 s 72006 0 72066 200 0 FreeSans 480 90 0 0 um_ow[116]
port 402 nsew signal input
flabel metal4 s 71270 0 71330 200 0 FreeSans 480 90 0 0 um_ow[117]
port 403 nsew signal input
flabel metal4 s 70534 0 70594 200 0 FreeSans 480 90 0 0 um_ow[118]
port 404 nsew signal input
flabel metal4 s 69798 0 69858 200 0 FreeSans 480 90 0 0 um_ow[119]
port 405 nsew signal input
flabel metal4 s 10366 0 10426 200 0 FreeSans 480 90 0 0 um_ow[11]
port 406 nsew signal input
flabel metal4 s 86726 10680 86786 10880 0 FreeSans 480 90 0 0 um_ow[120]
port 407 nsew signal input
flabel metal4 s 85990 10680 86050 10880 0 FreeSans 480 90 0 0 um_ow[121]
port 408 nsew signal input
flabel metal4 s 85254 10680 85314 10880 0 FreeSans 480 90 0 0 um_ow[122]
port 409 nsew signal input
flabel metal4 s 84518 10680 84578 10880 0 FreeSans 480 90 0 0 um_ow[123]
port 410 nsew signal input
flabel metal4 s 83782 10680 83842 10880 0 FreeSans 480 90 0 0 um_ow[124]
port 411 nsew signal input
flabel metal4 s 83046 10680 83106 10880 0 FreeSans 480 90 0 0 um_ow[125]
port 412 nsew signal input
flabel metal4 s 82310 10680 82370 10880 0 FreeSans 480 90 0 0 um_ow[126]
port 413 nsew signal input
flabel metal4 s 81574 10680 81634 10880 0 FreeSans 480 90 0 0 um_ow[127]
port 414 nsew signal input
flabel metal4 s 80838 10680 80898 10880 0 FreeSans 480 90 0 0 um_ow[128]
port 415 nsew signal input
flabel metal4 s 80102 10680 80162 10880 0 FreeSans 480 90 0 0 um_ow[129]
port 416 nsew signal input
flabel metal4 s 9630 0 9690 200 0 FreeSans 480 90 0 0 um_ow[12]
port 417 nsew signal input
flabel metal4 s 79366 10680 79426 10880 0 FreeSans 480 90 0 0 um_ow[130]
port 418 nsew signal input
flabel metal4 s 78630 10680 78690 10880 0 FreeSans 480 90 0 0 um_ow[131]
port 419 nsew signal input
flabel metal4 s 77894 10680 77954 10880 0 FreeSans 480 90 0 0 um_ow[132]
port 420 nsew signal input
flabel metal4 s 77158 10680 77218 10880 0 FreeSans 480 90 0 0 um_ow[133]
port 421 nsew signal input
flabel metal4 s 76422 10680 76482 10880 0 FreeSans 480 90 0 0 um_ow[134]
port 422 nsew signal input
flabel metal4 s 75686 10680 75746 10880 0 FreeSans 480 90 0 0 um_ow[135]
port 423 nsew signal input
flabel metal4 s 74950 10680 75010 10880 0 FreeSans 480 90 0 0 um_ow[136]
port 424 nsew signal input
flabel metal4 s 74214 10680 74274 10880 0 FreeSans 480 90 0 0 um_ow[137]
port 425 nsew signal input
flabel metal4 s 73478 10680 73538 10880 0 FreeSans 480 90 0 0 um_ow[138]
port 426 nsew signal input
flabel metal4 s 72742 10680 72802 10880 0 FreeSans 480 90 0 0 um_ow[139]
port 427 nsew signal input
flabel metal4 s 8894 0 8954 200 0 FreeSans 480 90 0 0 um_ow[13]
port 428 nsew signal input
flabel metal4 s 72006 10680 72066 10880 0 FreeSans 480 90 0 0 um_ow[140]
port 429 nsew signal input
flabel metal4 s 71270 10680 71330 10880 0 FreeSans 480 90 0 0 um_ow[141]
port 430 nsew signal input
flabel metal4 s 70534 10680 70594 10880 0 FreeSans 480 90 0 0 um_ow[142]
port 431 nsew signal input
flabel metal4 s 69798 10680 69858 10880 0 FreeSans 480 90 0 0 um_ow[143]
port 432 nsew signal input
flabel metal4 s 120858 0 120918 200 0 FreeSans 480 90 0 0 um_ow[144]
port 433 nsew signal input
flabel metal4 s 120122 0 120182 200 0 FreeSans 480 90 0 0 um_ow[145]
port 434 nsew signal input
flabel metal4 s 119386 0 119446 200 0 FreeSans 480 90 0 0 um_ow[146]
port 435 nsew signal input
flabel metal4 s 118650 0 118710 200 0 FreeSans 480 90 0 0 um_ow[147]
port 436 nsew signal input
flabel metal4 s 117914 0 117974 200 0 FreeSans 480 90 0 0 um_ow[148]
port 437 nsew signal input
flabel metal4 s 117178 0 117238 200 0 FreeSans 480 90 0 0 um_ow[149]
port 438 nsew signal input
flabel metal4 s 8158 0 8218 200 0 FreeSans 480 90 0 0 um_ow[14]
port 439 nsew signal input
flabel metal4 s 116442 0 116502 200 0 FreeSans 480 90 0 0 um_ow[150]
port 440 nsew signal input
flabel metal4 s 115706 0 115766 200 0 FreeSans 480 90 0 0 um_ow[151]
port 441 nsew signal input
flabel metal4 s 114970 0 115030 200 0 FreeSans 480 90 0 0 um_ow[152]
port 442 nsew signal input
flabel metal4 s 114234 0 114294 200 0 FreeSans 480 90 0 0 um_ow[153]
port 443 nsew signal input
flabel metal4 s 113498 0 113558 200 0 FreeSans 480 90 0 0 um_ow[154]
port 444 nsew signal input
flabel metal4 s 112762 0 112822 200 0 FreeSans 480 90 0 0 um_ow[155]
port 445 nsew signal input
flabel metal4 s 112026 0 112086 200 0 FreeSans 480 90 0 0 um_ow[156]
port 446 nsew signal input
flabel metal4 s 111290 0 111350 200 0 FreeSans 480 90 0 0 um_ow[157]
port 447 nsew signal input
flabel metal4 s 110554 0 110614 200 0 FreeSans 480 90 0 0 um_ow[158]
port 448 nsew signal input
flabel metal4 s 109818 0 109878 200 0 FreeSans 480 90 0 0 um_ow[159]
port 449 nsew signal input
flabel metal4 s 7422 0 7482 200 0 FreeSans 480 90 0 0 um_ow[15]
port 450 nsew signal input
flabel metal4 s 109082 0 109142 200 0 FreeSans 480 90 0 0 um_ow[160]
port 451 nsew signal input
flabel metal4 s 108346 0 108406 200 0 FreeSans 480 90 0 0 um_ow[161]
port 452 nsew signal input
flabel metal4 s 107610 0 107670 200 0 FreeSans 480 90 0 0 um_ow[162]
port 453 nsew signal input
flabel metal4 s 106874 0 106934 200 0 FreeSans 480 90 0 0 um_ow[163]
port 454 nsew signal input
flabel metal4 s 106138 0 106198 200 0 FreeSans 480 90 0 0 um_ow[164]
port 455 nsew signal input
flabel metal4 s 105402 0 105462 200 0 FreeSans 480 90 0 0 um_ow[165]
port 456 nsew signal input
flabel metal4 s 104666 0 104726 200 0 FreeSans 480 90 0 0 um_ow[166]
port 457 nsew signal input
flabel metal4 s 103930 0 103990 200 0 FreeSans 480 90 0 0 um_ow[167]
port 458 nsew signal input
flabel metal4 s 120858 10680 120918 10880 0 FreeSans 480 90 0 0 um_ow[168]
port 459 nsew signal input
flabel metal4 s 120122 10680 120182 10880 0 FreeSans 480 90 0 0 um_ow[169]
port 460 nsew signal input
flabel metal4 s 6686 0 6746 200 0 FreeSans 480 90 0 0 um_ow[16]
port 461 nsew signal input
flabel metal4 s 119386 10680 119446 10880 0 FreeSans 480 90 0 0 um_ow[170]
port 462 nsew signal input
flabel metal4 s 118650 10680 118710 10880 0 FreeSans 480 90 0 0 um_ow[171]
port 463 nsew signal input
flabel metal4 s 117914 10680 117974 10880 0 FreeSans 480 90 0 0 um_ow[172]
port 464 nsew signal input
flabel metal4 s 117178 10680 117238 10880 0 FreeSans 480 90 0 0 um_ow[173]
port 465 nsew signal input
flabel metal4 s 116442 10680 116502 10880 0 FreeSans 480 90 0 0 um_ow[174]
port 466 nsew signal input
flabel metal4 s 115706 10680 115766 10880 0 FreeSans 480 90 0 0 um_ow[175]
port 467 nsew signal input
flabel metal4 s 114970 10680 115030 10880 0 FreeSans 480 90 0 0 um_ow[176]
port 468 nsew signal input
flabel metal4 s 114234 10680 114294 10880 0 FreeSans 480 90 0 0 um_ow[177]
port 469 nsew signal input
flabel metal4 s 113498 10680 113558 10880 0 FreeSans 480 90 0 0 um_ow[178]
port 470 nsew signal input
flabel metal4 s 112762 10680 112822 10880 0 FreeSans 480 90 0 0 um_ow[179]
port 471 nsew signal input
flabel metal4 s 5950 0 6010 200 0 FreeSans 480 90 0 0 um_ow[17]
port 472 nsew signal input
flabel metal4 s 112026 10680 112086 10880 0 FreeSans 480 90 0 0 um_ow[180]
port 473 nsew signal input
flabel metal4 s 111290 10680 111350 10880 0 FreeSans 480 90 0 0 um_ow[181]
port 474 nsew signal input
flabel metal4 s 110554 10680 110614 10880 0 FreeSans 480 90 0 0 um_ow[182]
port 475 nsew signal input
flabel metal4 s 109818 10680 109878 10880 0 FreeSans 480 90 0 0 um_ow[183]
port 476 nsew signal input
flabel metal4 s 109082 10680 109142 10880 0 FreeSans 480 90 0 0 um_ow[184]
port 477 nsew signal input
flabel metal4 s 108346 10680 108406 10880 0 FreeSans 480 90 0 0 um_ow[185]
port 478 nsew signal input
flabel metal4 s 107610 10680 107670 10880 0 FreeSans 480 90 0 0 um_ow[186]
port 479 nsew signal input
flabel metal4 s 106874 10680 106934 10880 0 FreeSans 480 90 0 0 um_ow[187]
port 480 nsew signal input
flabel metal4 s 106138 10680 106198 10880 0 FreeSans 480 90 0 0 um_ow[188]
port 481 nsew signal input
flabel metal4 s 105402 10680 105462 10880 0 FreeSans 480 90 0 0 um_ow[189]
port 482 nsew signal input
flabel metal4 s 5214 0 5274 200 0 FreeSans 480 90 0 0 um_ow[18]
port 483 nsew signal input
flabel metal4 s 104666 10680 104726 10880 0 FreeSans 480 90 0 0 um_ow[190]
port 484 nsew signal input
flabel metal4 s 103930 10680 103990 10880 0 FreeSans 480 90 0 0 um_ow[191]
port 485 nsew signal input
flabel metal4 s 154990 0 155050 200 0 FreeSans 480 90 0 0 um_ow[192]
port 486 nsew signal input
flabel metal4 s 154254 0 154314 200 0 FreeSans 480 90 0 0 um_ow[193]
port 487 nsew signal input
flabel metal4 s 153518 0 153578 200 0 FreeSans 480 90 0 0 um_ow[194]
port 488 nsew signal input
flabel metal4 s 152782 0 152842 200 0 FreeSans 480 90 0 0 um_ow[195]
port 489 nsew signal input
flabel metal4 s 152046 0 152106 200 0 FreeSans 480 90 0 0 um_ow[196]
port 490 nsew signal input
flabel metal4 s 151310 0 151370 200 0 FreeSans 480 90 0 0 um_ow[197]
port 491 nsew signal input
flabel metal4 s 150574 0 150634 200 0 FreeSans 480 90 0 0 um_ow[198]
port 492 nsew signal input
flabel metal4 s 149838 0 149898 200 0 FreeSans 480 90 0 0 um_ow[199]
port 493 nsew signal input
flabel metal4 s 4478 0 4538 200 0 FreeSans 480 90 0 0 um_ow[19]
port 494 nsew signal input
flabel metal4 s 17726 0 17786 200 0 FreeSans 480 90 0 0 um_ow[1]
port 495 nsew signal input
flabel metal4 s 149102 0 149162 200 0 FreeSans 480 90 0 0 um_ow[200]
port 496 nsew signal input
flabel metal4 s 148366 0 148426 200 0 FreeSans 480 90 0 0 um_ow[201]
port 497 nsew signal input
flabel metal4 s 147630 0 147690 200 0 FreeSans 480 90 0 0 um_ow[202]
port 498 nsew signal input
flabel metal4 s 146894 0 146954 200 0 FreeSans 480 90 0 0 um_ow[203]
port 499 nsew signal input
flabel metal4 s 146158 0 146218 200 0 FreeSans 480 90 0 0 um_ow[204]
port 500 nsew signal input
flabel metal4 s 145422 0 145482 200 0 FreeSans 480 90 0 0 um_ow[205]
port 501 nsew signal input
flabel metal4 s 144686 0 144746 200 0 FreeSans 480 90 0 0 um_ow[206]
port 502 nsew signal input
flabel metal4 s 143950 0 144010 200 0 FreeSans 480 90 0 0 um_ow[207]
port 503 nsew signal input
flabel metal4 s 143214 0 143274 200 0 FreeSans 480 90 0 0 um_ow[208]
port 504 nsew signal input
flabel metal4 s 142478 0 142538 200 0 FreeSans 480 90 0 0 um_ow[209]
port 505 nsew signal input
flabel metal4 s 3742 0 3802 200 0 FreeSans 480 90 0 0 um_ow[20]
port 506 nsew signal input
flabel metal4 s 141742 0 141802 200 0 FreeSans 480 90 0 0 um_ow[210]
port 507 nsew signal input
flabel metal4 s 141006 0 141066 200 0 FreeSans 480 90 0 0 um_ow[211]
port 508 nsew signal input
flabel metal4 s 140270 0 140330 200 0 FreeSans 480 90 0 0 um_ow[212]
port 509 nsew signal input
flabel metal4 s 139534 0 139594 200 0 FreeSans 480 90 0 0 um_ow[213]
port 510 nsew signal input
flabel metal4 s 138798 0 138858 200 0 FreeSans 480 90 0 0 um_ow[214]
port 511 nsew signal input
flabel metal4 s 138062 0 138122 200 0 FreeSans 480 90 0 0 um_ow[215]
port 512 nsew signal input
flabel metal4 s 154990 10680 155050 10880 0 FreeSans 480 90 0 0 um_ow[216]
port 513 nsew signal input
flabel metal4 s 154254 10680 154314 10880 0 FreeSans 480 90 0 0 um_ow[217]
port 514 nsew signal input
flabel metal4 s 153518 10680 153578 10880 0 FreeSans 480 90 0 0 um_ow[218]
port 515 nsew signal input
flabel metal4 s 152782 10680 152842 10880 0 FreeSans 480 90 0 0 um_ow[219]
port 516 nsew signal input
flabel metal4 s 3006 0 3066 200 0 FreeSans 480 90 0 0 um_ow[21]
port 517 nsew signal input
flabel metal4 s 152046 10680 152106 10880 0 FreeSans 480 90 0 0 um_ow[220]
port 518 nsew signal input
flabel metal4 s 151310 10680 151370 10880 0 FreeSans 480 90 0 0 um_ow[221]
port 519 nsew signal input
flabel metal4 s 150574 10680 150634 10880 0 FreeSans 480 90 0 0 um_ow[222]
port 520 nsew signal input
flabel metal4 s 149838 10680 149898 10880 0 FreeSans 480 90 0 0 um_ow[223]
port 521 nsew signal input
flabel metal4 s 149102 10680 149162 10880 0 FreeSans 480 90 0 0 um_ow[224]
port 522 nsew signal input
flabel metal4 s 148366 10680 148426 10880 0 FreeSans 480 90 0 0 um_ow[225]
port 523 nsew signal input
flabel metal4 s 147630 10680 147690 10880 0 FreeSans 480 90 0 0 um_ow[226]
port 524 nsew signal input
flabel metal4 s 146894 10680 146954 10880 0 FreeSans 480 90 0 0 um_ow[227]
port 525 nsew signal input
flabel metal4 s 146158 10680 146218 10880 0 FreeSans 480 90 0 0 um_ow[228]
port 526 nsew signal input
flabel metal4 s 145422 10680 145482 10880 0 FreeSans 480 90 0 0 um_ow[229]
port 527 nsew signal input
flabel metal4 s 2270 0 2330 200 0 FreeSans 480 90 0 0 um_ow[22]
port 528 nsew signal input
flabel metal4 s 144686 10680 144746 10880 0 FreeSans 480 90 0 0 um_ow[230]
port 529 nsew signal input
flabel metal4 s 143950 10680 144010 10880 0 FreeSans 480 90 0 0 um_ow[231]
port 530 nsew signal input
flabel metal4 s 143214 10680 143274 10880 0 FreeSans 480 90 0 0 um_ow[232]
port 531 nsew signal input
flabel metal4 s 142478 10680 142538 10880 0 FreeSans 480 90 0 0 um_ow[233]
port 532 nsew signal input
flabel metal4 s 141742 10680 141802 10880 0 FreeSans 480 90 0 0 um_ow[234]
port 533 nsew signal input
flabel metal4 s 141006 10680 141066 10880 0 FreeSans 480 90 0 0 um_ow[235]
port 534 nsew signal input
flabel metal4 s 140270 10680 140330 10880 0 FreeSans 480 90 0 0 um_ow[236]
port 535 nsew signal input
flabel metal4 s 139534 10680 139594 10880 0 FreeSans 480 90 0 0 um_ow[237]
port 536 nsew signal input
flabel metal4 s 138798 10680 138858 10880 0 FreeSans 480 90 0 0 um_ow[238]
port 537 nsew signal input
flabel metal4 s 138062 10680 138122 10880 0 FreeSans 480 90 0 0 um_ow[239]
port 538 nsew signal input
flabel metal4 s 1534 0 1594 200 0 FreeSans 480 90 0 0 um_ow[23]
port 539 nsew signal input
flabel metal4 s 189122 0 189182 200 0 FreeSans 480 90 0 0 um_ow[240]
port 540 nsew signal input
flabel metal4 s 188386 0 188446 200 0 FreeSans 480 90 0 0 um_ow[241]
port 541 nsew signal input
flabel metal4 s 187650 0 187710 200 0 FreeSans 480 90 0 0 um_ow[242]
port 542 nsew signal input
flabel metal4 s 186914 0 186974 200 0 FreeSans 480 90 0 0 um_ow[243]
port 543 nsew signal input
flabel metal4 s 186178 0 186238 200 0 FreeSans 480 90 0 0 um_ow[244]
port 544 nsew signal input
flabel metal4 s 185442 0 185502 200 0 FreeSans 480 90 0 0 um_ow[245]
port 545 nsew signal input
flabel metal4 s 184706 0 184766 200 0 FreeSans 480 90 0 0 um_ow[246]
port 546 nsew signal input
flabel metal4 s 183970 0 184030 200 0 FreeSans 480 90 0 0 um_ow[247]
port 547 nsew signal input
flabel metal4 s 183234 0 183294 200 0 FreeSans 480 90 0 0 um_ow[248]
port 548 nsew signal input
flabel metal4 s 182498 0 182558 200 0 FreeSans 480 90 0 0 um_ow[249]
port 549 nsew signal input
flabel metal4 s 18462 10680 18522 10880 0 FreeSans 480 90 0 0 um_ow[24]
port 550 nsew signal input
flabel metal4 s 181762 0 181822 200 0 FreeSans 480 90 0 0 um_ow[250]
port 551 nsew signal input
flabel metal4 s 181026 0 181086 200 0 FreeSans 480 90 0 0 um_ow[251]
port 552 nsew signal input
flabel metal4 s 180290 0 180350 200 0 FreeSans 480 90 0 0 um_ow[252]
port 553 nsew signal input
flabel metal4 s 179554 0 179614 200 0 FreeSans 480 90 0 0 um_ow[253]
port 554 nsew signal input
flabel metal4 s 178818 0 178878 200 0 FreeSans 480 90 0 0 um_ow[254]
port 555 nsew signal input
flabel metal4 s 178082 0 178142 200 0 FreeSans 480 90 0 0 um_ow[255]
port 556 nsew signal input
flabel metal4 s 177346 0 177406 200 0 FreeSans 480 90 0 0 um_ow[256]
port 557 nsew signal input
flabel metal4 s 176610 0 176670 200 0 FreeSans 480 90 0 0 um_ow[257]
port 558 nsew signal input
flabel metal4 s 175874 0 175934 200 0 FreeSans 480 90 0 0 um_ow[258]
port 559 nsew signal input
flabel metal4 s 175138 0 175198 200 0 FreeSans 480 90 0 0 um_ow[259]
port 560 nsew signal input
flabel metal4 s 17726 10680 17786 10880 0 FreeSans 480 90 0 0 um_ow[25]
port 561 nsew signal input
flabel metal4 s 174402 0 174462 200 0 FreeSans 480 90 0 0 um_ow[260]
port 562 nsew signal input
flabel metal4 s 173666 0 173726 200 0 FreeSans 480 90 0 0 um_ow[261]
port 563 nsew signal input
flabel metal4 s 172930 0 172990 200 0 FreeSans 480 90 0 0 um_ow[262]
port 564 nsew signal input
flabel metal4 s 172194 0 172254 200 0 FreeSans 480 90 0 0 um_ow[263]
port 565 nsew signal input
flabel metal4 s 189122 10680 189182 10880 0 FreeSans 480 90 0 0 um_ow[264]
port 566 nsew signal input
flabel metal4 s 188386 10680 188446 10880 0 FreeSans 480 90 0 0 um_ow[265]
port 567 nsew signal input
flabel metal4 s 187650 10680 187710 10880 0 FreeSans 480 90 0 0 um_ow[266]
port 568 nsew signal input
flabel metal4 s 186914 10680 186974 10880 0 FreeSans 480 90 0 0 um_ow[267]
port 569 nsew signal input
flabel metal4 s 186178 10680 186238 10880 0 FreeSans 480 90 0 0 um_ow[268]
port 570 nsew signal input
flabel metal4 s 185442 10680 185502 10880 0 FreeSans 480 90 0 0 um_ow[269]
port 571 nsew signal input
flabel metal4 s 16990 10680 17050 10880 0 FreeSans 480 90 0 0 um_ow[26]
port 572 nsew signal input
flabel metal4 s 184706 10680 184766 10880 0 FreeSans 480 90 0 0 um_ow[270]
port 573 nsew signal input
flabel metal4 s 183970 10680 184030 10880 0 FreeSans 480 90 0 0 um_ow[271]
port 574 nsew signal input
flabel metal4 s 183234 10680 183294 10880 0 FreeSans 480 90 0 0 um_ow[272]
port 575 nsew signal input
flabel metal4 s 182498 10680 182558 10880 0 FreeSans 480 90 0 0 um_ow[273]
port 576 nsew signal input
flabel metal4 s 181762 10680 181822 10880 0 FreeSans 480 90 0 0 um_ow[274]
port 577 nsew signal input
flabel metal4 s 181026 10680 181086 10880 0 FreeSans 480 90 0 0 um_ow[275]
port 578 nsew signal input
flabel metal4 s 180290 10680 180350 10880 0 FreeSans 480 90 0 0 um_ow[276]
port 579 nsew signal input
flabel metal4 s 179554 10680 179614 10880 0 FreeSans 480 90 0 0 um_ow[277]
port 580 nsew signal input
flabel metal4 s 178818 10680 178878 10880 0 FreeSans 480 90 0 0 um_ow[278]
port 581 nsew signal input
flabel metal4 s 178082 10680 178142 10880 0 FreeSans 480 90 0 0 um_ow[279]
port 582 nsew signal input
flabel metal4 s 16254 10680 16314 10880 0 FreeSans 480 90 0 0 um_ow[27]
port 583 nsew signal input
flabel metal4 s 177346 10680 177406 10880 0 FreeSans 480 90 0 0 um_ow[280]
port 584 nsew signal input
flabel metal4 s 176610 10680 176670 10880 0 FreeSans 480 90 0 0 um_ow[281]
port 585 nsew signal input
flabel metal4 s 175874 10680 175934 10880 0 FreeSans 480 90 0 0 um_ow[282]
port 586 nsew signal input
flabel metal4 s 175138 10680 175198 10880 0 FreeSans 480 90 0 0 um_ow[283]
port 587 nsew signal input
flabel metal4 s 174402 10680 174462 10880 0 FreeSans 480 90 0 0 um_ow[284]
port 588 nsew signal input
flabel metal4 s 173666 10680 173726 10880 0 FreeSans 480 90 0 0 um_ow[285]
port 589 nsew signal input
flabel metal4 s 172930 10680 172990 10880 0 FreeSans 480 90 0 0 um_ow[286]
port 590 nsew signal input
flabel metal4 s 172194 10680 172254 10880 0 FreeSans 480 90 0 0 um_ow[287]
port 591 nsew signal input
flabel metal4 s 223254 0 223314 200 0 FreeSans 480 90 0 0 um_ow[288]
port 592 nsew signal input
flabel metal4 s 222518 0 222578 200 0 FreeSans 480 90 0 0 um_ow[289]
port 593 nsew signal input
flabel metal4 s 15518 10680 15578 10880 0 FreeSans 480 90 0 0 um_ow[28]
port 594 nsew signal input
flabel metal4 s 221782 0 221842 200 0 FreeSans 480 90 0 0 um_ow[290]
port 595 nsew signal input
flabel metal4 s 221046 0 221106 200 0 FreeSans 480 90 0 0 um_ow[291]
port 596 nsew signal input
flabel metal4 s 220310 0 220370 200 0 FreeSans 480 90 0 0 um_ow[292]
port 597 nsew signal input
flabel metal4 s 219574 0 219634 200 0 FreeSans 480 90 0 0 um_ow[293]
port 598 nsew signal input
flabel metal4 s 218838 0 218898 200 0 FreeSans 480 90 0 0 um_ow[294]
port 599 nsew signal input
flabel metal4 s 218102 0 218162 200 0 FreeSans 480 90 0 0 um_ow[295]
port 600 nsew signal input
flabel metal4 s 217366 0 217426 200 0 FreeSans 480 90 0 0 um_ow[296]
port 601 nsew signal input
flabel metal4 s 216630 0 216690 200 0 FreeSans 480 90 0 0 um_ow[297]
port 602 nsew signal input
flabel metal4 s 215894 0 215954 200 0 FreeSans 480 90 0 0 um_ow[298]
port 603 nsew signal input
flabel metal4 s 215158 0 215218 200 0 FreeSans 480 90 0 0 um_ow[299]
port 604 nsew signal input
flabel metal4 s 14782 10680 14842 10880 0 FreeSans 480 90 0 0 um_ow[29]
port 605 nsew signal input
flabel metal4 s 16990 0 17050 200 0 FreeSans 480 90 0 0 um_ow[2]
port 606 nsew signal input
flabel metal4 s 214422 0 214482 200 0 FreeSans 480 90 0 0 um_ow[300]
port 607 nsew signal input
flabel metal4 s 213686 0 213746 200 0 FreeSans 480 90 0 0 um_ow[301]
port 608 nsew signal input
flabel metal4 s 212950 0 213010 200 0 FreeSans 480 90 0 0 um_ow[302]
port 609 nsew signal input
flabel metal4 s 212214 0 212274 200 0 FreeSans 480 90 0 0 um_ow[303]
port 610 nsew signal input
flabel metal4 s 211478 0 211538 200 0 FreeSans 480 90 0 0 um_ow[304]
port 611 nsew signal input
flabel metal4 s 210742 0 210802 200 0 FreeSans 480 90 0 0 um_ow[305]
port 612 nsew signal input
flabel metal4 s 210006 0 210066 200 0 FreeSans 480 90 0 0 um_ow[306]
port 613 nsew signal input
flabel metal4 s 209270 0 209330 200 0 FreeSans 480 90 0 0 um_ow[307]
port 614 nsew signal input
flabel metal4 s 208534 0 208594 200 0 FreeSans 480 90 0 0 um_ow[308]
port 615 nsew signal input
flabel metal4 s 207798 0 207858 200 0 FreeSans 480 90 0 0 um_ow[309]
port 616 nsew signal input
flabel metal4 s 14046 10680 14106 10880 0 FreeSans 480 90 0 0 um_ow[30]
port 617 nsew signal input
flabel metal4 s 207062 0 207122 200 0 FreeSans 480 90 0 0 um_ow[310]
port 618 nsew signal input
flabel metal4 s 206326 0 206386 200 0 FreeSans 480 90 0 0 um_ow[311]
port 619 nsew signal input
flabel metal4 s 223254 10680 223314 10880 0 FreeSans 480 90 0 0 um_ow[312]
port 620 nsew signal input
flabel metal4 s 222518 10680 222578 10880 0 FreeSans 480 90 0 0 um_ow[313]
port 621 nsew signal input
flabel metal4 s 221782 10680 221842 10880 0 FreeSans 480 90 0 0 um_ow[314]
port 622 nsew signal input
flabel metal4 s 221046 10680 221106 10880 0 FreeSans 480 90 0 0 um_ow[315]
port 623 nsew signal input
flabel metal4 s 220310 10680 220370 10880 0 FreeSans 480 90 0 0 um_ow[316]
port 624 nsew signal input
flabel metal4 s 219574 10680 219634 10880 0 FreeSans 480 90 0 0 um_ow[317]
port 625 nsew signal input
flabel metal4 s 218838 10680 218898 10880 0 FreeSans 480 90 0 0 um_ow[318]
port 626 nsew signal input
flabel metal4 s 218102 10680 218162 10880 0 FreeSans 480 90 0 0 um_ow[319]
port 627 nsew signal input
flabel metal4 s 13310 10680 13370 10880 0 FreeSans 480 90 0 0 um_ow[31]
port 628 nsew signal input
flabel metal4 s 217366 10680 217426 10880 0 FreeSans 480 90 0 0 um_ow[320]
port 629 nsew signal input
flabel metal4 s 216630 10680 216690 10880 0 FreeSans 480 90 0 0 um_ow[321]
port 630 nsew signal input
flabel metal4 s 215894 10680 215954 10880 0 FreeSans 480 90 0 0 um_ow[322]
port 631 nsew signal input
flabel metal4 s 215158 10680 215218 10880 0 FreeSans 480 90 0 0 um_ow[323]
port 632 nsew signal input
flabel metal4 s 214422 10680 214482 10880 0 FreeSans 480 90 0 0 um_ow[324]
port 633 nsew signal input
flabel metal4 s 213686 10680 213746 10880 0 FreeSans 480 90 0 0 um_ow[325]
port 634 nsew signal input
flabel metal4 s 212950 10680 213010 10880 0 FreeSans 480 90 0 0 um_ow[326]
port 635 nsew signal input
flabel metal4 s 212214 10680 212274 10880 0 FreeSans 480 90 0 0 um_ow[327]
port 636 nsew signal input
flabel metal4 s 211478 10680 211538 10880 0 FreeSans 480 90 0 0 um_ow[328]
port 637 nsew signal input
flabel metal4 s 210742 10680 210802 10880 0 FreeSans 480 90 0 0 um_ow[329]
port 638 nsew signal input
flabel metal4 s 12574 10680 12634 10880 0 FreeSans 480 90 0 0 um_ow[32]
port 639 nsew signal input
flabel metal4 s 210006 10680 210066 10880 0 FreeSans 480 90 0 0 um_ow[330]
port 640 nsew signal input
flabel metal4 s 209270 10680 209330 10880 0 FreeSans 480 90 0 0 um_ow[331]
port 641 nsew signal input
flabel metal4 s 208534 10680 208594 10880 0 FreeSans 480 90 0 0 um_ow[332]
port 642 nsew signal input
flabel metal4 s 207798 10680 207858 10880 0 FreeSans 480 90 0 0 um_ow[333]
port 643 nsew signal input
flabel metal4 s 207062 10680 207122 10880 0 FreeSans 480 90 0 0 um_ow[334]
port 644 nsew signal input
flabel metal4 s 206326 10680 206386 10880 0 FreeSans 480 90 0 0 um_ow[335]
port 645 nsew signal input
flabel metal4 s 257386 0 257446 200 0 FreeSans 480 90 0 0 um_ow[336]
port 646 nsew signal input
flabel metal4 s 256650 0 256710 200 0 FreeSans 480 90 0 0 um_ow[337]
port 647 nsew signal input
flabel metal4 s 255914 0 255974 200 0 FreeSans 480 90 0 0 um_ow[338]
port 648 nsew signal input
flabel metal4 s 255178 0 255238 200 0 FreeSans 480 90 0 0 um_ow[339]
port 649 nsew signal input
flabel metal4 s 11838 10680 11898 10880 0 FreeSans 480 90 0 0 um_ow[33]
port 650 nsew signal input
flabel metal4 s 254442 0 254502 200 0 FreeSans 480 90 0 0 um_ow[340]
port 651 nsew signal input
flabel metal4 s 253706 0 253766 200 0 FreeSans 480 90 0 0 um_ow[341]
port 652 nsew signal input
flabel metal4 s 252970 0 253030 200 0 FreeSans 480 90 0 0 um_ow[342]
port 653 nsew signal input
flabel metal4 s 252234 0 252294 200 0 FreeSans 480 90 0 0 um_ow[343]
port 654 nsew signal input
flabel metal4 s 251498 0 251558 200 0 FreeSans 480 90 0 0 um_ow[344]
port 655 nsew signal input
flabel metal4 s 250762 0 250822 200 0 FreeSans 480 90 0 0 um_ow[345]
port 656 nsew signal input
flabel metal4 s 250026 0 250086 200 0 FreeSans 480 90 0 0 um_ow[346]
port 657 nsew signal input
flabel metal4 s 249290 0 249350 200 0 FreeSans 480 90 0 0 um_ow[347]
port 658 nsew signal input
flabel metal4 s 248554 0 248614 200 0 FreeSans 480 90 0 0 um_ow[348]
port 659 nsew signal input
flabel metal4 s 247818 0 247878 200 0 FreeSans 480 90 0 0 um_ow[349]
port 660 nsew signal input
flabel metal4 s 11102 10680 11162 10880 0 FreeSans 480 90 0 0 um_ow[34]
port 661 nsew signal input
flabel metal4 s 247082 0 247142 200 0 FreeSans 480 90 0 0 um_ow[350]
port 662 nsew signal input
flabel metal4 s 246346 0 246406 200 0 FreeSans 480 90 0 0 um_ow[351]
port 663 nsew signal input
flabel metal4 s 245610 0 245670 200 0 FreeSans 480 90 0 0 um_ow[352]
port 664 nsew signal input
flabel metal4 s 244874 0 244934 200 0 FreeSans 480 90 0 0 um_ow[353]
port 665 nsew signal input
flabel metal4 s 244138 0 244198 200 0 FreeSans 480 90 0 0 um_ow[354]
port 666 nsew signal input
flabel metal4 s 243402 0 243462 200 0 FreeSans 480 90 0 0 um_ow[355]
port 667 nsew signal input
flabel metal4 s 242666 0 242726 200 0 FreeSans 480 90 0 0 um_ow[356]
port 668 nsew signal input
flabel metal4 s 241930 0 241990 200 0 FreeSans 480 90 0 0 um_ow[357]
port 669 nsew signal input
flabel metal4 s 241194 0 241254 200 0 FreeSans 480 90 0 0 um_ow[358]
port 670 nsew signal input
flabel metal4 s 240458 0 240518 200 0 FreeSans 480 90 0 0 um_ow[359]
port 671 nsew signal input
flabel metal4 s 10366 10680 10426 10880 0 FreeSans 480 90 0 0 um_ow[35]
port 672 nsew signal input
flabel metal4 s 257386 10680 257446 10880 0 FreeSans 480 90 0 0 um_ow[360]
port 673 nsew signal input
flabel metal4 s 256650 10680 256710 10880 0 FreeSans 480 90 0 0 um_ow[361]
port 674 nsew signal input
flabel metal4 s 255914 10680 255974 10880 0 FreeSans 480 90 0 0 um_ow[362]
port 675 nsew signal input
flabel metal4 s 255178 10680 255238 10880 0 FreeSans 480 90 0 0 um_ow[363]
port 676 nsew signal input
flabel metal4 s 254442 10680 254502 10880 0 FreeSans 480 90 0 0 um_ow[364]
port 677 nsew signal input
flabel metal4 s 253706 10680 253766 10880 0 FreeSans 480 90 0 0 um_ow[365]
port 678 nsew signal input
flabel metal4 s 252970 10680 253030 10880 0 FreeSans 480 90 0 0 um_ow[366]
port 679 nsew signal input
flabel metal4 s 252234 10680 252294 10880 0 FreeSans 480 90 0 0 um_ow[367]
port 680 nsew signal input
flabel metal4 s 251498 10680 251558 10880 0 FreeSans 480 90 0 0 um_ow[368]
port 681 nsew signal input
flabel metal4 s 250762 10680 250822 10880 0 FreeSans 480 90 0 0 um_ow[369]
port 682 nsew signal input
flabel metal4 s 9630 10680 9690 10880 0 FreeSans 480 90 0 0 um_ow[36]
port 683 nsew signal input
flabel metal4 s 250026 10680 250086 10880 0 FreeSans 480 90 0 0 um_ow[370]
port 684 nsew signal input
flabel metal4 s 249290 10680 249350 10880 0 FreeSans 480 90 0 0 um_ow[371]
port 685 nsew signal input
flabel metal4 s 248554 10680 248614 10880 0 FreeSans 480 90 0 0 um_ow[372]
port 686 nsew signal input
flabel metal4 s 247818 10680 247878 10880 0 FreeSans 480 90 0 0 um_ow[373]
port 687 nsew signal input
flabel metal4 s 247082 10680 247142 10880 0 FreeSans 480 90 0 0 um_ow[374]
port 688 nsew signal input
flabel metal4 s 246346 10680 246406 10880 0 FreeSans 480 90 0 0 um_ow[375]
port 689 nsew signal input
flabel metal4 s 245610 10680 245670 10880 0 FreeSans 480 90 0 0 um_ow[376]
port 690 nsew signal input
flabel metal4 s 244874 10680 244934 10880 0 FreeSans 480 90 0 0 um_ow[377]
port 691 nsew signal input
flabel metal4 s 244138 10680 244198 10880 0 FreeSans 480 90 0 0 um_ow[378]
port 692 nsew signal input
flabel metal4 s 243402 10680 243462 10880 0 FreeSans 480 90 0 0 um_ow[379]
port 693 nsew signal input
flabel metal4 s 8894 10680 8954 10880 0 FreeSans 480 90 0 0 um_ow[37]
port 694 nsew signal input
flabel metal4 s 242666 10680 242726 10880 0 FreeSans 480 90 0 0 um_ow[380]
port 695 nsew signal input
flabel metal4 s 241930 10680 241990 10880 0 FreeSans 480 90 0 0 um_ow[381]
port 696 nsew signal input
flabel metal4 s 241194 10680 241254 10880 0 FreeSans 480 90 0 0 um_ow[382]
port 697 nsew signal input
flabel metal4 s 240458 10680 240518 10880 0 FreeSans 480 90 0 0 um_ow[383]
port 698 nsew signal input
flabel metal4 s 8158 10680 8218 10880 0 FreeSans 480 90 0 0 um_ow[38]
port 699 nsew signal input
flabel metal4 s 7422 10680 7482 10880 0 FreeSans 480 90 0 0 um_ow[39]
port 700 nsew signal input
flabel metal4 s 16254 0 16314 200 0 FreeSans 480 90 0 0 um_ow[3]
port 701 nsew signal input
flabel metal4 s 6686 10680 6746 10880 0 FreeSans 480 90 0 0 um_ow[40]
port 702 nsew signal input
flabel metal4 s 5950 10680 6010 10880 0 FreeSans 480 90 0 0 um_ow[41]
port 703 nsew signal input
flabel metal4 s 5214 10680 5274 10880 0 FreeSans 480 90 0 0 um_ow[42]
port 704 nsew signal input
flabel metal4 s 4478 10680 4538 10880 0 FreeSans 480 90 0 0 um_ow[43]
port 705 nsew signal input
flabel metal4 s 3742 10680 3802 10880 0 FreeSans 480 90 0 0 um_ow[44]
port 706 nsew signal input
flabel metal4 s 3006 10680 3066 10880 0 FreeSans 480 90 0 0 um_ow[45]
port 707 nsew signal input
flabel metal4 s 2270 10680 2330 10880 0 FreeSans 480 90 0 0 um_ow[46]
port 708 nsew signal input
flabel metal4 s 1534 10680 1594 10880 0 FreeSans 480 90 0 0 um_ow[47]
port 709 nsew signal input
flabel metal4 s 52594 0 52654 200 0 FreeSans 480 90 0 0 um_ow[48]
port 710 nsew signal input
flabel metal4 s 51858 0 51918 200 0 FreeSans 480 90 0 0 um_ow[49]
port 711 nsew signal input
flabel metal4 s 15518 0 15578 200 0 FreeSans 480 90 0 0 um_ow[4]
port 712 nsew signal input
flabel metal4 s 51122 0 51182 200 0 FreeSans 480 90 0 0 um_ow[50]
port 713 nsew signal input
flabel metal4 s 50386 0 50446 200 0 FreeSans 480 90 0 0 um_ow[51]
port 714 nsew signal input
flabel metal4 s 49650 0 49710 200 0 FreeSans 480 90 0 0 um_ow[52]
port 715 nsew signal input
flabel metal4 s 48914 0 48974 200 0 FreeSans 480 90 0 0 um_ow[53]
port 716 nsew signal input
flabel metal4 s 48178 0 48238 200 0 FreeSans 480 90 0 0 um_ow[54]
port 717 nsew signal input
flabel metal4 s 47442 0 47502 200 0 FreeSans 480 90 0 0 um_ow[55]
port 718 nsew signal input
flabel metal4 s 46706 0 46766 200 0 FreeSans 480 90 0 0 um_ow[56]
port 719 nsew signal input
flabel metal4 s 45970 0 46030 200 0 FreeSans 480 90 0 0 um_ow[57]
port 720 nsew signal input
flabel metal4 s 45234 0 45294 200 0 FreeSans 480 90 0 0 um_ow[58]
port 721 nsew signal input
flabel metal4 s 44498 0 44558 200 0 FreeSans 480 90 0 0 um_ow[59]
port 722 nsew signal input
flabel metal4 s 14782 0 14842 200 0 FreeSans 480 90 0 0 um_ow[5]
port 723 nsew signal input
flabel metal4 s 43762 0 43822 200 0 FreeSans 480 90 0 0 um_ow[60]
port 724 nsew signal input
flabel metal4 s 43026 0 43086 200 0 FreeSans 480 90 0 0 um_ow[61]
port 725 nsew signal input
flabel metal4 s 42290 0 42350 200 0 FreeSans 480 90 0 0 um_ow[62]
port 726 nsew signal input
flabel metal4 s 41554 0 41614 200 0 FreeSans 480 90 0 0 um_ow[63]
port 727 nsew signal input
flabel metal4 s 40818 0 40878 200 0 FreeSans 480 90 0 0 um_ow[64]
port 728 nsew signal input
flabel metal4 s 40082 0 40142 200 0 FreeSans 480 90 0 0 um_ow[65]
port 729 nsew signal input
flabel metal4 s 39346 0 39406 200 0 FreeSans 480 90 0 0 um_ow[66]
port 730 nsew signal input
flabel metal4 s 38610 0 38670 200 0 FreeSans 480 90 0 0 um_ow[67]
port 731 nsew signal input
flabel metal4 s 37874 0 37934 200 0 FreeSans 480 90 0 0 um_ow[68]
port 732 nsew signal input
flabel metal4 s 37138 0 37198 200 0 FreeSans 480 90 0 0 um_ow[69]
port 733 nsew signal input
flabel metal4 s 14046 0 14106 200 0 FreeSans 480 90 0 0 um_ow[6]
port 734 nsew signal input
flabel metal4 s 36402 0 36462 200 0 FreeSans 480 90 0 0 um_ow[70]
port 735 nsew signal input
flabel metal4 s 35666 0 35726 200 0 FreeSans 480 90 0 0 um_ow[71]
port 736 nsew signal input
flabel metal4 s 52594 10680 52654 10880 0 FreeSans 480 90 0 0 um_ow[72]
port 737 nsew signal input
flabel metal4 s 51858 10680 51918 10880 0 FreeSans 480 90 0 0 um_ow[73]
port 738 nsew signal input
flabel metal4 s 51122 10680 51182 10880 0 FreeSans 480 90 0 0 um_ow[74]
port 739 nsew signal input
flabel metal4 s 50386 10680 50446 10880 0 FreeSans 480 90 0 0 um_ow[75]
port 740 nsew signal input
flabel metal4 s 49650 10680 49710 10880 0 FreeSans 480 90 0 0 um_ow[76]
port 741 nsew signal input
flabel metal4 s 48914 10680 48974 10880 0 FreeSans 480 90 0 0 um_ow[77]
port 742 nsew signal input
flabel metal4 s 48178 10680 48238 10880 0 FreeSans 480 90 0 0 um_ow[78]
port 743 nsew signal input
flabel metal4 s 47442 10680 47502 10880 0 FreeSans 480 90 0 0 um_ow[79]
port 744 nsew signal input
flabel metal4 s 13310 0 13370 200 0 FreeSans 480 90 0 0 um_ow[7]
port 745 nsew signal input
flabel metal4 s 46706 10680 46766 10880 0 FreeSans 480 90 0 0 um_ow[80]
port 746 nsew signal input
flabel metal4 s 45970 10680 46030 10880 0 FreeSans 480 90 0 0 um_ow[81]
port 747 nsew signal input
flabel metal4 s 45234 10680 45294 10880 0 FreeSans 480 90 0 0 um_ow[82]
port 748 nsew signal input
flabel metal4 s 44498 10680 44558 10880 0 FreeSans 480 90 0 0 um_ow[83]
port 749 nsew signal input
flabel metal4 s 43762 10680 43822 10880 0 FreeSans 480 90 0 0 um_ow[84]
port 750 nsew signal input
flabel metal4 s 43026 10680 43086 10880 0 FreeSans 480 90 0 0 um_ow[85]
port 751 nsew signal input
flabel metal4 s 42290 10680 42350 10880 0 FreeSans 480 90 0 0 um_ow[86]
port 752 nsew signal input
flabel metal4 s 41554 10680 41614 10880 0 FreeSans 480 90 0 0 um_ow[87]
port 753 nsew signal input
flabel metal4 s 40818 10680 40878 10880 0 FreeSans 480 90 0 0 um_ow[88]
port 754 nsew signal input
flabel metal4 s 40082 10680 40142 10880 0 FreeSans 480 90 0 0 um_ow[89]
port 755 nsew signal input
flabel metal4 s 12574 0 12634 200 0 FreeSans 480 90 0 0 um_ow[8]
port 756 nsew signal input
flabel metal4 s 39346 10680 39406 10880 0 FreeSans 480 90 0 0 um_ow[90]
port 757 nsew signal input
flabel metal4 s 38610 10680 38670 10880 0 FreeSans 480 90 0 0 um_ow[91]
port 758 nsew signal input
flabel metal4 s 37874 10680 37934 10880 0 FreeSans 480 90 0 0 um_ow[92]
port 759 nsew signal input
flabel metal4 s 37138 10680 37198 10880 0 FreeSans 480 90 0 0 um_ow[93]
port 760 nsew signal input
flabel metal4 s 36402 10680 36462 10880 0 FreeSans 480 90 0 0 um_ow[94]
port 761 nsew signal input
flabel metal4 s 35666 10680 35726 10880 0 FreeSans 480 90 0 0 um_ow[95]
port 762 nsew signal input
flabel metal4 s 86726 0 86786 200 0 FreeSans 480 90 0 0 um_ow[96]
port 763 nsew signal input
flabel metal4 s 85990 0 86050 200 0 FreeSans 480 90 0 0 um_ow[97]
port 764 nsew signal input
flabel metal4 s 85254 0 85314 200 0 FreeSans 480 90 0 0 um_ow[98]
port 765 nsew signal input
flabel metal4 s 84518 0 84578 200 0 FreeSans 480 90 0 0 um_ow[99]
port 766 nsew signal input
flabel metal4 s 11838 0 11898 200 0 FreeSans 480 90 0 0 um_ow[9]
port 767 nsew signal input
flabel metal4 s 34742 1040 35062 9840 0 FreeSans 1920 90 0 0 vccd1
port 768 nsew power bidirectional
flabel metal4 s 102339 1040 102659 9840 0 FreeSans 1920 90 0 0 vccd1
port 768 nsew power bidirectional
flabel metal4 s 169936 1040 170256 9840 0 FreeSans 1920 90 0 0 vccd1
port 768 nsew power bidirectional
flabel metal4 s 237533 1040 237853 9840 0 FreeSans 1920 90 0 0 vccd1
port 768 nsew power bidirectional
flabel metal4 s 68540 1040 68860 9840 0 FreeSans 1920 90 0 0 vssd1
port 769 nsew ground bidirectional
flabel metal4 s 136137 1040 136457 9840 0 FreeSans 1920 90 0 0 vssd1
port 769 nsew ground bidirectional
flabel metal4 s 203734 1040 204054 9840 0 FreeSans 1920 90 0 0 vssd1
port 769 nsew ground bidirectional
flabel metal4 s 271331 1040 271651 9840 0 FreeSans 1920 90 0 0 vssd1
port 769 nsew ground bidirectional
rlabel metal1 136298 9248 136298 9248 0 vccd1
rlabel via1 136377 9792 136377 9792 0 vssd1
rlabel metal1 270802 7514 270802 7514 0 _0000_
rlabel metal2 267122 9418 267122 9418 0 _0001_
rlabel metal2 253874 4658 253874 4658 0 _0002_
rlabel metal1 270388 6834 270388 6834 0 _0003_
rlabel metal1 269698 7786 269698 7786 0 _0004_
rlabel metal1 251436 5270 251436 5270 0 _0005_
rlabel metal2 252862 4250 252862 4250 0 _0006_
rlabel metal2 269238 7242 269238 7242 0 _0007_
rlabel metal2 249826 5916 249826 5916 0 _0008_
rlabel metal1 252908 4658 252908 4658 0 _0009_
rlabel metal1 270158 7446 270158 7446 0 _0010_
rlabel via1 269600 7378 269600 7378 0 _0011_
rlabel metal1 253414 5712 253414 5712 0 _0012_
rlabel metal1 253322 4182 253322 4182 0 _0013_
rlabel metal2 255898 4794 255898 4794 0 _0014_
rlabel metal1 258106 4114 258106 4114 0 _0015_
rlabel metal2 254058 5100 254058 5100 0 _0016_
rlabel metal2 253874 6154 253874 6154 0 _0017_
rlabel metal1 259072 3366 259072 3366 0 _0018_
rlabel metal2 259210 5236 259210 5236 0 _0019_
rlabel metal1 259026 4080 259026 4080 0 _0020_
rlabel metal2 256726 6596 256726 6596 0 _0021_
rlabel metal1 253322 5134 253322 5134 0 _0022_
rlabel metal2 247250 1156 247250 1156 0 _0023_
rlabel metal1 246974 1530 246974 1530 0 _0024_
rlabel metal1 251574 4658 251574 4658 0 _0025_
rlabel metal1 247296 1326 247296 1326 0 _0026_
rlabel metal1 244766 4114 244766 4114 0 _0027_
rlabel metal2 248262 6086 248262 6086 0 _0028_
rlabel metal1 253184 3638 253184 3638 0 _0029_
rlabel metal1 252264 4454 252264 4454 0 _0030_
rlabel metal2 246698 4454 246698 4454 0 _0031_
rlabel metal2 245594 3978 245594 3978 0 _0032_
rlabel metal2 244674 4828 244674 4828 0 _0033_
rlabel metal1 251942 5270 251942 5270 0 _0034_
rlabel metal1 244720 3162 244720 3162 0 _0035_
rlabel metal1 245778 1326 245778 1326 0 _0036_
rlabel metal2 249366 6596 249366 6596 0 _0037_
rlabel metal2 250746 5610 250746 5610 0 _0038_
rlabel metal2 259854 5066 259854 5066 0 _0039_
rlabel metal2 248170 5746 248170 5746 0 _0040_
rlabel metal2 116794 6630 116794 6630 0 _0041_
rlabel metal1 135930 5780 135930 5780 0 _0042_
rlabel metal1 108284 6222 108284 6222 0 _0043_
rlabel metal2 133262 6222 133262 6222 0 _0044_
rlabel metal1 136114 5542 136114 5542 0 _0045_
rlabel metal2 128110 6154 128110 6154 0 _0046_
rlabel metal2 167026 1343 167026 1343 0 _0047_
rlabel metal1 112378 4624 112378 4624 0 _0048_
rlabel metal2 114494 4930 114494 4930 0 _0049_
rlabel metal1 113068 4590 113068 4590 0 _0050_
rlabel metal2 114218 4556 114218 4556 0 _0051_
rlabel metal1 113666 4624 113666 4624 0 _0052_
rlabel metal2 108606 6528 108606 6528 0 _0053_
rlabel metal1 109802 7412 109802 7412 0 _0054_
rlabel metal1 106490 5712 106490 5712 0 _0055_
rlabel metal2 109066 7174 109066 7174 0 _0056_
rlabel metal2 109342 7140 109342 7140 0 _0057_
rlabel metal1 97152 5678 97152 5678 0 _0058_
rlabel metal2 96646 5474 96646 5474 0 _0059_
rlabel metal1 101614 6154 101614 6154 0 _0060_
rlabel metal2 102350 6562 102350 6562 0 _0061_
rlabel metal1 101522 5814 101522 5814 0 _0062_
rlabel metal1 103040 5202 103040 5202 0 _0063_
rlabel metal1 103638 5712 103638 5712 0 _0064_
rlabel metal1 102120 3706 102120 3706 0 _0065_
rlabel metal2 116058 5712 116058 5712 0 _0066_
rlabel metal2 98762 6902 98762 6902 0 _0067_
rlabel metal1 92782 3468 92782 3468 0 _0068_
rlabel metal2 92966 4063 92966 4063 0 _0069_
rlabel metal2 98670 6120 98670 6120 0 _0070_
rlabel metal1 93610 5168 93610 5168 0 _0071_
rlabel metal2 94714 6188 94714 6188 0 _0072_
rlabel metal2 96186 6324 96186 6324 0 _0073_
rlabel metal2 118174 6562 118174 6562 0 _0074_
rlabel metal1 137678 5066 137678 5066 0 _0075_
rlabel metal2 137494 4998 137494 4998 0 _0076_
rlabel metal2 168314 4828 168314 4828 0 _0077_
rlabel metal1 122866 3502 122866 3502 0 _0078_
rlabel metal2 121854 4998 121854 4998 0 _0079_
rlabel metal1 121486 3978 121486 3978 0 _0080_
rlabel metal1 118910 4624 118910 4624 0 _0081_
rlabel metal1 120152 1938 120152 1938 0 _0082_
rlabel metal2 110538 3502 110538 3502 0 _0083_
rlabel metal1 104742 4148 104742 4148 0 _0084_
rlabel metal1 111228 4250 111228 4250 0 _0085_
rlabel metal1 109894 4114 109894 4114 0 _0086_
rlabel metal1 109802 2992 109802 2992 0 _0087_
rlabel metal1 109204 3910 109204 3910 0 _0088_
rlabel metal2 107226 6392 107226 6392 0 _0089_
rlabel metal1 105478 4624 105478 4624 0 _0090_
rlabel metal1 107548 4454 107548 4454 0 _0091_
rlabel metal1 104880 4590 104880 4590 0 _0092_
rlabel metal1 106444 3706 106444 3706 0 _0093_
rlabel metal2 106490 5508 106490 5508 0 _0094_
rlabel metal2 105294 4828 105294 4828 0 _0095_
rlabel metal2 148534 5899 148534 5899 0 _0096_
rlabel metal1 116886 5848 116886 5848 0 _0097_
rlabel metal1 101292 4794 101292 4794 0 _0098_
rlabel metal1 101660 5338 101660 5338 0 _0099_
rlabel metal1 98854 6392 98854 6392 0 _0100_
rlabel metal1 100464 5338 100464 5338 0 _0101_
rlabel metal2 95266 6562 95266 6562 0 _0102_
rlabel metal2 97934 6052 97934 6052 0 _0103_
rlabel metal1 98992 5338 98992 5338 0 _0104_
rlabel metal1 169188 4590 169188 4590 0 _0105_
rlabel metal2 148810 6732 148810 6732 0 _0106_
rlabel metal1 149592 5814 149592 5814 0 _0107_
rlabel metal1 147706 3910 147706 3910 0 _0108_
rlabel metal2 147982 4896 147982 4896 0 _0109_
rlabel metal1 150374 5066 150374 5066 0 _0110_
rlabel metal1 148672 4046 148672 4046 0 _0111_
rlabel metal1 152674 2482 152674 2482 0 _0112_
rlabel metal1 154652 3026 154652 3026 0 _0113_
rlabel viali 150282 6289 150282 6289 0 _0114_
rlabel metal1 149546 5712 149546 5712 0 _0115_
rlabel metal1 150512 4114 150512 4114 0 _0116_
rlabel metal1 152950 3026 152950 3026 0 _0117_
rlabel metal1 153962 3060 153962 3060 0 _0118_
rlabel metal2 152766 3706 152766 3706 0 _0119_
rlabel metal1 148488 4250 148488 4250 0 _0120_
rlabel metal1 139610 3944 139610 3944 0 _0121_
rlabel metal1 138920 4114 138920 4114 0 _0122_
rlabel metal2 143658 4998 143658 4998 0 _0123_
rlabel metal1 138782 5066 138782 5066 0 _0124_
rlabel metal1 145038 4148 145038 4148 0 _0125_
rlabel metal1 145038 5236 145038 5236 0 _0126_
rlabel metal1 143842 3978 143842 3978 0 _0127_
rlabel metal1 139840 2278 139840 2278 0 _0128_
rlabel metal1 141588 2278 141588 2278 0 _0129_
rlabel metal2 139058 3196 139058 3196 0 _0130_
rlabel metal1 138736 3502 138736 3502 0 _0131_
rlabel metal2 139150 4148 139150 4148 0 _0132_
rlabel metal2 139702 3468 139702 3468 0 _0133_
rlabel metal1 223008 3502 223008 3502 0 _0134_
rlabel metal1 223606 3060 223606 3060 0 _0135_
rlabel metal2 222778 3196 222778 3196 0 _0136_
rlabel metal1 208794 2414 208794 2414 0 _0137_
rlabel metal1 209116 2414 209116 2414 0 _0138_
rlabel metal2 208978 2587 208978 2587 0 _0139_
rlabel metal1 248860 5814 248860 5814 0 _0140_
rlabel metal1 138092 5066 138092 5066 0 _0141_
rlabel metal1 113022 6256 113022 6256 0 _0142_
rlabel metal1 111136 6766 111136 6766 0 _0143_
rlabel metal1 68770 3536 68770 3536 0 _0144_
rlabel metal2 137218 5984 137218 5984 0 _0145_
rlabel via1 115782 7786 115782 7786 0 _0146_
rlabel metal2 135562 6018 135562 6018 0 _0147_
rlabel metal2 189382 6562 189382 6562 0 _0148_
rlabel metal2 78798 7327 78798 7327 0 _0149_
rlabel metal1 66930 4080 66930 4080 0 _0150_
rlabel via2 76590 7395 76590 7395 0 _0151_
rlabel metal2 99314 7650 99314 7650 0 _0152_
rlabel metal2 118174 7004 118174 7004 0 _0153_
rlabel metal1 109802 8024 109802 8024 0 _0154_
rlabel metal1 120842 5678 120842 5678 0 _0155_
rlabel metal1 119646 6426 119646 6426 0 _0156_
rlabel metal1 167992 3502 167992 3502 0 _0157_
rlabel metal2 189566 5950 189566 5950 0 _0158_
rlabel metal2 169050 6766 169050 6766 0 _0159_
rlabel metal2 190486 4964 190486 4964 0 _0160_
rlabel metal2 189750 6596 189750 6596 0 _0161_
rlabel metal1 224342 3502 224342 3502 0 _0162_
rlabel via1 217074 6630 217074 6630 0 _0163_
rlabel metal1 217718 5882 217718 5882 0 _0164_
rlabel metal2 227286 6579 227286 6579 0 _0165_
rlabel metal2 216890 7106 216890 7106 0 _0166_
rlabel metal2 248906 5950 248906 5950 0 _0167_
rlabel metal1 253759 4522 253759 4522 0 _0168_
rlabel metal1 256174 4046 256174 4046 0 _0169_
rlabel metal2 255346 5848 255346 5848 0 _0170_
rlabel metal2 254242 5457 254242 5457 0 _0171_
rlabel metal1 256542 2516 256542 2516 0 _0172_
rlabel metal1 256726 5542 256726 5542 0 _0173_
rlabel metal1 255346 2924 255346 2924 0 _0174_
rlabel metal2 256634 5644 256634 5644 0 _0175_
rlabel metal2 253966 4216 253966 4216 0 _0176_
rlabel metal1 244812 4046 244812 4046 0 _0177_
rlabel metal1 248768 3094 248768 3094 0 _0178_
rlabel metal1 248814 2482 248814 2482 0 _0179_
rlabel metal1 251896 1190 251896 1190 0 _0180_
rlabel metal2 245134 4046 245134 4046 0 _0181_
rlabel metal1 245226 2006 245226 2006 0 _0182_
rlabel metal1 250976 6086 250976 6086 0 _0183_
rlabel metal1 250378 918 250378 918 0 _0184_
rlabel metal1 248216 1870 248216 1870 0 _0185_
rlabel metal1 245824 1190 245824 1190 0 _0186_
rlabel metal1 248998 3570 248998 3570 0 _0187_
rlabel metal1 249182 4046 249182 4046 0 _0188_
rlabel metal2 259854 4318 259854 4318 0 _0189_
rlabel metal2 249090 5372 249090 5372 0 _0190_
rlabel metal2 110998 5950 110998 5950 0 _0191_
rlabel metal2 117530 7684 117530 7684 0 _0192_
rlabel metal1 114448 2482 114448 2482 0 _0193_
rlabel metal2 115230 4148 115230 4148 0 _0194_
rlabel metal1 114264 4522 114264 4522 0 _0195_
rlabel metal1 114954 4012 114954 4012 0 _0196_
rlabel metal1 115000 3570 115000 3570 0 _0197_
rlabel metal2 109250 6460 109250 6460 0 _0198_
rlabel metal1 108698 4726 108698 4726 0 _0199_
rlabel metal2 109802 6800 109802 6800 0 _0200_
rlabel metal1 109342 7718 109342 7718 0 _0201_
rlabel metal1 101844 3094 101844 3094 0 _0202_
rlabel metal1 101614 1870 101614 1870 0 _0203_
rlabel metal1 102350 6630 102350 6630 0 _0204_
rlabel metal1 102856 4658 102856 4658 0 _0205_
rlabel metal1 102626 4046 102626 4046 0 _0206_
rlabel metal2 99774 4590 99774 4590 0 _0207_
rlabel metal2 99314 5372 99314 5372 0 _0208_
rlabel via2 92598 3723 92598 3723 0 _0209_
rlabel metal1 96232 3094 96232 3094 0 _0210_
rlabel via1 96646 5797 96646 5797 0 _0211_
rlabel metal2 94530 4828 94530 4828 0 _0212_
rlabel metal2 97474 5338 97474 5338 0 _0213_
rlabel metal1 95266 5134 95266 5134 0 _0214_
rlabel metal1 113390 6426 113390 6426 0 _0215_
rlabel metal2 117530 5440 117530 5440 0 _0216_
rlabel metal2 122498 3876 122498 3876 0 _0217_
rlabel metal1 121302 2958 121302 2958 0 _0218_
rlabel metal1 121302 3570 121302 3570 0 _0219_
rlabel metal1 119232 2482 119232 2482 0 _0220_
rlabel metal1 119278 1734 119278 1734 0 _0221_
rlabel metal2 111826 4250 111826 4250 0 _0222_
rlabel metal1 112286 3434 112286 3434 0 _0223_
rlabel metal1 112010 2924 112010 2924 0 _0224_
rlabel metal2 112378 2553 112378 2553 0 _0225_
rlabel metal1 105777 4454 105777 4454 0 _0226_
rlabel metal1 107686 2006 107686 2006 0 _0227_
rlabel metal1 106812 3094 106812 3094 0 _0228_
rlabel metal2 106122 4063 106122 4063 0 _0229_
rlabel metal2 105938 5066 105938 5066 0 _0230_
rlabel metal1 104926 5542 104926 5542 0 _0231_
rlabel metal2 99682 4556 99682 4556 0 _0232_
rlabel metal1 99728 2006 99728 2006 0 _0233_
rlabel metal1 97060 2482 97060 2482 0 _0234_
rlabel metal1 97106 4012 97106 4012 0 _0235_
rlabel metal2 94806 5066 94806 5066 0 _0236_
rlabel metal2 97750 5916 97750 5916 0 _0237_
rlabel metal1 96140 6358 96140 6358 0 _0238_
rlabel metal1 140484 5746 140484 5746 0 _0239_
rlabel metal1 169510 4726 169510 4726 0 _0240_
rlabel metal2 158470 5100 158470 5100 0 _0241_
rlabel metal1 156078 2958 156078 2958 0 _0242_
rlabel metal2 153410 6052 153410 6052 0 _0243_
rlabel metal1 153594 2618 153594 2618 0 _0244_
rlabel metal1 155342 3162 155342 3162 0 _0245_
rlabel metal2 153594 5083 153594 5083 0 _0246_
rlabel metal1 152996 5270 152996 5270 0 _0247_
rlabel metal1 150558 4046 150558 4046 0 _0248_
rlabel metal1 151018 2924 151018 2924 0 _0249_
rlabel metal1 152122 3162 152122 3162 0 _0250_
rlabel metal1 150972 2482 150972 2482 0 _0251_
rlabel metal1 148534 4454 148534 4454 0 _0252_
rlabel metal1 145866 5100 145866 5100 0 _0253_
rlabel metal2 145590 3672 145590 3672 0 _0254_
rlabel metal1 145774 3094 145774 3094 0 _0255_
rlabel metal1 144486 2482 144486 2482 0 _0256_
rlabel metal1 139334 2618 139334 2618 0 _0257_
rlabel metal2 138276 2516 138276 2516 0 _0258_
rlabel metal1 141082 2822 141082 2822 0 _0259_
rlabel metal1 139518 3094 139518 3094 0 _0260_
rlabel metal1 139840 3706 139840 3706 0 _0261_
rlabel metal2 139518 3162 139518 3162 0 _0262_
rlabel metal2 216522 5474 216522 5474 0 _0263_
rlabel metal1 213302 5644 213302 5644 0 _0264_
rlabel metal2 221582 4590 221582 4590 0 _0265_
rlabel metal1 223836 1258 223836 1258 0 _0266_
rlabel metal1 224940 4522 224940 4522 0 _0267_
rlabel metal2 223146 5678 223146 5678 0 _0268_
rlabel metal2 220938 3298 220938 3298 0 _0269_
rlabel metal1 220248 5270 220248 5270 0 _0270_
rlabel metal2 218178 5372 218178 5372 0 _0271_
rlabel metal1 217258 3434 217258 3434 0 _0272_
rlabel metal1 218362 1190 218362 1190 0 _0273_
rlabel metal1 221260 2346 221260 2346 0 _0274_
rlabel metal1 213440 2958 213440 2958 0 _0275_
rlabel metal2 215142 3264 215142 3264 0 _0276_
rlabel metal1 212750 4046 212750 4046 0 _0277_
rlabel via2 214774 4675 214774 4675 0 _0278_
rlabel metal1 212428 3094 212428 3094 0 _0279_
rlabel metal1 212474 3026 212474 3026 0 _0280_
rlabel metal1 210174 2346 210174 2346 0 _0281_
rlabel metal1 208748 1870 208748 1870 0 _0282_
rlabel metal2 209990 4250 209990 4250 0 _0283_
rlabel metal1 207690 4012 207690 4012 0 _0284_
rlabel metal1 207230 5338 207230 5338 0 _0285_
rlabel metal1 206356 4522 206356 4522 0 _0286_
rlabel metal1 270342 9554 270342 9554 0 addr[0]
rlabel metal3 272282 9452 272282 9452 0 addr[1]
rlabel metal3 270212 9316 270212 9316 0 addr[2]
rlabel metal3 270580 9180 270580 9180 0 addr[3]
rlabel metal3 270534 9044 270534 9044 0 addr[4]
rlabel metal2 114586 6103 114586 6103 0 bus_ow\[0\]
rlabel metal1 111918 2482 111918 2482 0 bus_ow\[10\]
rlabel metal1 180780 6936 180780 6936 0 bus_ow\[11\]
rlabel metal2 213486 714 213486 714 0 bus_ow\[12\]
rlabel metal4 110308 4012 110308 4012 0 bus_ow\[13\]
rlabel metal2 226320 1292 226320 1292 0 bus_ow\[14\]
rlabel metal2 244858 1054 244858 1054 0 bus_ow\[15\]
rlabel metal2 248538 1649 248538 1649 0 bus_ow\[16\]
rlabel metal2 230598 1428 230598 1428 0 bus_ow\[17\]
rlabel metal2 177054 1054 177054 1054 0 bus_ow\[18\]
rlabel metal2 209806 1445 209806 1445 0 bus_ow\[19\]
rlabel metal3 243524 2448 243524 2448 0 bus_ow\[1\]
rlabel metal3 122820 748 122820 748 0 bus_ow\[20\]
rlabel metal2 176686 3655 176686 3655 0 bus_ow\[21\]
rlabel metal2 98486 5474 98486 5474 0 bus_ow\[22\]
rlabel metal2 214590 1071 214590 1071 0 bus_ow\[23\]
rlabel metal1 121532 2482 121532 2482 0 bus_ow\[2\]
rlabel metal1 133630 2040 133630 2040 0 bus_ow\[3\]
rlabel metal2 167946 5236 167946 5236 0 bus_ow\[4\]
rlabel metal1 116610 3978 116610 3978 0 bus_ow\[5\]
rlabel metal3 152674 1156 152674 1156 0 bus_ow\[6\]
rlabel metal1 112056 4046 112056 4046 0 bus_ow\[7\]
rlabel metal2 154790 6613 154790 6613 0 bus_ow\[8\]
rlabel metal1 112378 6358 112378 6358 0 bus_ow\[9\]
rlabel metal2 53314 5593 53314 5593 0 col\[0\].genblk1.mux4_I\[0\].x
rlabel metal2 108514 1581 108514 1581 0 col\[0\].genblk1.mux4_I\[10\].x
rlabel metal1 64860 3468 64860 3468 0 col\[0\].genblk1.mux4_I\[11\].x
rlabel metal3 93840 2380 93840 2380 0 col\[0\].genblk1.mux4_I\[12\].x
rlabel metal1 101016 2482 101016 2482 0 col\[0\].genblk1.mux4_I\[13\].x
rlabel metal2 42826 5355 42826 5355 0 col\[0\].genblk1.mux4_I\[14\].x
rlabel metal2 92690 3859 92690 3859 0 col\[0\].genblk1.mux4_I\[15\].x
rlabel metal2 41538 2176 41538 2176 0 col\[0\].genblk1.mux4_I\[16\].x
rlabel via2 40434 1717 40434 1717 0 col\[0\].genblk1.mux4_I\[17\].x
rlabel metal2 39882 1377 39882 1377 0 col\[0\].genblk1.mux4_I\[18\].x
rlabel via2 38962 3995 38962 3995 0 col\[0\].genblk1.mux4_I\[19\].x
rlabel metal1 52256 5066 52256 5066 0 col\[0\].genblk1.mux4_I\[1\].x
rlabel metal1 39054 3162 39054 3162 0 col\[0\].genblk1.mux4_I\[20\].x
rlabel metal2 39514 3264 39514 3264 0 col\[0\].genblk1.mux4_I\[21\].x
rlabel via2 36846 4981 36846 4981 0 col\[0\].genblk1.mux4_I\[22\].x
rlabel metal2 37030 5066 37030 5066 0 col\[0\].genblk1.mux4_I\[23\].x
rlabel metal3 96094 2652 96094 2652 0 col\[0\].genblk1.mux4_I\[2\].x
rlabel metal2 51842 3417 51842 3417 0 col\[0\].genblk1.mux4_I\[3\].x
rlabel metal2 55890 4386 55890 4386 0 col\[0\].genblk1.mux4_I\[4\].x
rlabel metal3 93840 1020 93840 1020 0 col\[0\].genblk1.mux4_I\[5\].x
rlabel metal2 114954 3213 114954 3213 0 col\[0\].genblk1.mux4_I\[6\].x
rlabel metal1 51382 6256 51382 6256 0 col\[0\].genblk1.mux4_I\[7\].x
rlabel metal2 109158 4845 109158 4845 0 col\[0\].genblk1.mux4_I\[8\].x
rlabel metal1 60720 6732 60720 6732 0 col\[0\].genblk1.mux4_I\[9\].x
rlabel metal2 67666 3349 67666 3349 0 col\[0\].zbuf_bot_ena_I.e
rlabel metal1 32936 1938 32936 1938 0 col\[0\].zbuf_bot_ena_I.z
rlabel metal2 179446 7871 179446 7871 0 col\[0\].zbuf_bot_iw_I\[0\].a
rlabel metal2 32338 1530 32338 1530 0 col\[0\].zbuf_bot_iw_I\[0\].z
rlabel metal2 180550 816 180550 816 0 col\[0\].zbuf_bot_iw_I\[10\].a
rlabel metal1 23736 2618 23736 2618 0 col\[0\].zbuf_bot_iw_I\[10\].z
rlabel metal2 170798 6936 170798 6936 0 col\[0\].zbuf_bot_iw_I\[11\].a
rlabel metal1 23322 3502 23322 3502 0 col\[0\].zbuf_bot_iw_I\[11\].z
rlabel metal2 194534 9214 194534 9214 0 col\[0\].zbuf_bot_iw_I\[12\].a
rlabel metal1 21988 2414 21988 2414 0 col\[0\].zbuf_bot_iw_I\[12\].z
rlabel metal2 229034 9860 229034 9860 0 col\[0\].zbuf_bot_iw_I\[13\].a
rlabel metal1 21712 1938 21712 1938 0 col\[0\].zbuf_bot_iw_I\[13\].z
rlabel metal2 168406 833 168406 833 0 col\[0\].zbuf_bot_iw_I\[14\].a
rlabel metal2 22126 1530 22126 1530 0 col\[0\].zbuf_bot_iw_I\[14\].z
rlabel metal2 230414 1088 230414 1088 0 col\[0\].zbuf_bot_iw_I\[15\].a
rlabel metal1 23782 1938 23782 1938 0 col\[0\].zbuf_bot_iw_I\[15\].z
rlabel metal1 209760 748 209760 748 0 col\[0\].zbuf_bot_iw_I\[16\].a
rlabel metal1 24518 1326 24518 1326 0 col\[0\].zbuf_bot_iw_I\[16\].z
rlabel metal3 233703 1292 233703 1292 0 col\[0\].zbuf_bot_iw_I\[17\].a
rlabel metal2 25898 2142 25898 2142 0 col\[0\].zbuf_bot_iw_I\[17\].z
rlabel metal1 180780 8500 180780 8500 0 col\[0\].zbuf_bot_iw_I\[1\].a
rlabel metal2 31050 1530 31050 1530 0 col\[0\].zbuf_bot_iw_I\[1\].z
rlabel via2 215234 9707 215234 9707 0 col\[0\].zbuf_bot_iw_I\[2\].a
rlabel metal1 30360 1326 30360 1326 0 col\[0\].zbuf_bot_iw_I\[2\].z
rlabel metal2 246974 8483 246974 8483 0 col\[0\].zbuf_bot_iw_I\[3\].a
rlabel metal2 29762 2142 29762 2142 0 col\[0\].zbuf_bot_iw_I\[3\].z
rlabel metal2 226550 1564 226550 1564 0 col\[0\].zbuf_bot_iw_I\[4\].a
rlabel metal2 28842 1530 28842 1530 0 col\[0\].zbuf_bot_iw_I\[4\].z
rlabel metal2 168866 8568 168866 8568 0 col\[0\].zbuf_bot_iw_I\[5\].a
rlabel metal2 28014 1530 28014 1530 0 col\[0\].zbuf_bot_iw_I\[5\].z
rlabel metal2 228390 8143 228390 8143 0 col\[0\].zbuf_bot_iw_I\[6\].a
rlabel metal1 27508 1530 27508 1530 0 col\[0\].zbuf_bot_iw_I\[6\].z
rlabel metal2 230322 867 230322 867 0 col\[0\].zbuf_bot_iw_I\[7\].a
rlabel metal1 26312 3026 26312 3026 0 col\[0\].zbuf_bot_iw_I\[7\].z
rlabel metal1 228758 10540 228758 10540 0 col\[0\].zbuf_bot_iw_I\[8\].a
rlabel metal1 25530 3026 25530 3026 0 col\[0\].zbuf_bot_iw_I\[8\].z
rlabel metal1 214038 8466 214038 8466 0 col\[0\].zbuf_bot_iw_I\[9\].a
rlabel metal1 24610 2822 24610 2822 0 col\[0\].zbuf_bot_iw_I\[9\].z
rlabel metal1 64860 7208 64860 7208 0 col\[0\].zbuf_top_ena_I.e
rlabel metal2 33166 8772 33166 8772 0 col\[0\].zbuf_top_ena_I.z
rlabel metal2 32154 9350 32154 9350 0 col\[0\].zbuf_top_iw_I\[0\].z
rlabel metal2 24058 8772 24058 8772 0 col\[0\].zbuf_top_iw_I\[10\].z
rlabel metal2 23506 8092 23506 8092 0 col\[0\].zbuf_top_iw_I\[11\].z
rlabel metal2 22770 8330 22770 8330 0 col\[0\].zbuf_top_iw_I\[12\].z
rlabel metal2 20286 9146 20286 9146 0 col\[0\].zbuf_top_iw_I\[13\].z
rlabel metal1 21643 8466 21643 8466 0 col\[0\].zbuf_top_iw_I\[14\].z
rlabel metal1 21712 7854 21712 7854 0 col\[0\].zbuf_top_iw_I\[15\].z
rlabel metal2 22954 9146 22954 9146 0 col\[0\].zbuf_top_iw_I\[16\].z
rlabel metal2 24702 9146 24702 9146 0 col\[0\].zbuf_top_iw_I\[17\].z
rlabel metal2 30866 8636 30866 8636 0 col\[0\].zbuf_top_iw_I\[1\].z
rlabel metal2 30406 9350 30406 9350 0 col\[0\].zbuf_top_iw_I\[2\].z
rlabel metal2 29854 9078 29854 9078 0 col\[0\].zbuf_top_iw_I\[3\].z
rlabel metal2 28750 8636 28750 8636 0 col\[0\].zbuf_top_iw_I\[4\].z
rlabel metal2 28014 8636 28014 8636 0 col\[0\].zbuf_top_iw_I\[5\].z
rlabel metal2 27278 8636 27278 8636 0 col\[0\].zbuf_top_iw_I\[6\].z
rlabel metal2 26542 9078 26542 9078 0 col\[0\].zbuf_top_iw_I\[7\].z
rlabel metal1 26128 9554 26128 9554 0 col\[0\].zbuf_top_iw_I\[8\].z
rlabel metal2 25070 8058 25070 8058 0 col\[0\].zbuf_top_iw_I\[9\].z
rlabel metal1 66562 2380 66562 2380 0 col\[1\].zbuf_bot_ena_I.e
rlabel metal1 66884 1938 66884 1938 0 col\[1\].zbuf_bot_ena_I.z
rlabel metal1 66608 1326 66608 1326 0 col\[1\].zbuf_bot_iw_I\[0\].z
rlabel metal1 58420 1530 58420 1530 0 col\[1\].zbuf_bot_iw_I\[10\].z
rlabel metal2 57546 2210 57546 2210 0 col\[1\].zbuf_bot_iw_I\[11\].z
rlabel metal2 56994 1530 56994 1530 0 col\[1\].zbuf_bot_iw_I\[12\].z
rlabel metal2 56258 1530 56258 1530 0 col\[1\].zbuf_bot_iw_I\[13\].z
rlabel metal2 55062 1530 55062 1530 0 col\[1\].zbuf_bot_iw_I\[14\].z
rlabel metal2 55522 2210 55522 2210 0 col\[1\].zbuf_bot_iw_I\[15\].z
rlabel metal1 54510 3026 54510 3026 0 col\[1\].zbuf_bot_iw_I\[16\].z
rlabel metal1 53268 1938 53268 1938 0 col\[1\].zbuf_bot_iw_I\[17\].z
rlabel metal2 65458 2210 65458 2210 0 col\[1\].zbuf_bot_iw_I\[1\].z
rlabel metal2 64446 1530 64446 1530 0 col\[1\].zbuf_bot_iw_I\[2\].z
rlabel metal2 63710 1530 63710 1530 0 col\[1\].zbuf_bot_iw_I\[3\].z
rlabel metal2 62698 2210 62698 2210 0 col\[1\].zbuf_bot_iw_I\[4\].z
rlabel metal1 62330 1530 62330 1530 0 col\[1\].zbuf_bot_iw_I\[5\].z
rlabel metal2 61686 2210 61686 2210 0 col\[1\].zbuf_bot_iw_I\[6\].z
rlabel metal2 60766 1530 60766 1530 0 col\[1\].zbuf_bot_iw_I\[7\].z
rlabel metal2 59846 1530 59846 1530 0 col\[1\].zbuf_bot_iw_I\[8\].z
rlabel metal2 59202 2210 59202 2210 0 col\[1\].zbuf_bot_iw_I\[9\].z
rlabel metal2 76406 8568 76406 8568 0 col\[1\].zbuf_top_ena_I.e
rlabel metal1 67160 8058 67160 8058 0 col\[1\].zbuf_top_ena_I.z
rlabel metal2 66102 8636 66102 8636 0 col\[1\].zbuf_top_iw_I\[0\].z
rlabel metal1 58466 8466 58466 8466 0 col\[1\].zbuf_top_iw_I\[10\].z
rlabel metal1 57684 9146 57684 9146 0 col\[1\].zbuf_top_iw_I\[11\].z
rlabel metal2 57362 9078 57362 9078 0 col\[1\].zbuf_top_iw_I\[12\].z
rlabel metal2 56626 9350 56626 9350 0 col\[1\].zbuf_top_iw_I\[13\].z
rlabel metal2 55890 8772 55890 8772 0 col\[1\].zbuf_top_iw_I\[14\].z
rlabel metal2 54970 9350 54970 9350 0 col\[1\].zbuf_top_iw_I\[15\].z
rlabel metal1 54280 8602 54280 8602 0 col\[1\].zbuf_top_iw_I\[16\].z
rlabel metal2 53130 9146 53130 9146 0 col\[1\].zbuf_top_iw_I\[17\].z
rlabel metal2 65366 8636 65366 8636 0 col\[1\].zbuf_top_iw_I\[1\].z
rlabel metal2 64538 8636 64538 8636 0 col\[1\].zbuf_top_iw_I\[2\].z
rlabel metal2 63802 8636 63802 8636 0 col\[1\].zbuf_top_iw_I\[3\].z
rlabel metal2 62790 9350 62790 9350 0 col\[1\].zbuf_top_iw_I\[4\].z
rlabel metal2 62606 9078 62606 9078 0 col\[1\].zbuf_top_iw_I\[5\].z
rlabel metal2 62238 9350 62238 9350 0 col\[1\].zbuf_top_iw_I\[6\].z
rlabel metal2 60858 8636 60858 8636 0 col\[1\].zbuf_top_iw_I\[7\].z
rlabel metal2 60122 8636 60122 8636 0 col\[1\].zbuf_top_iw_I\[8\].z
rlabel metal2 59386 8636 59386 8636 0 col\[1\].zbuf_top_iw_I\[9\].z
rlabel metal2 113758 7004 113758 7004 0 col\[2\].genblk1.mux4_I\[0\].x
rlabel metal1 113114 1190 113114 1190 0 col\[2\].genblk1.mux4_I\[10\].x
rlabel metal2 109066 1972 109066 1972 0 col\[2\].genblk1.mux4_I\[11\].x
rlabel metal1 106996 1870 106996 1870 0 col\[2\].genblk1.mux4_I\[12\].x
rlabel metal1 106858 2958 106858 2958 0 col\[2\].genblk1.mux4_I\[13\].x
rlabel metal2 106306 3332 106306 3332 0 col\[2\].genblk1.mux4_I\[14\].x
rlabel metal2 105386 3876 105386 3876 0 col\[2\].genblk1.mux4_I\[15\].x
rlabel metal2 101522 1836 101522 1836 0 col\[2\].genblk1.mux4_I\[16\].x
rlabel metal2 98762 2244 98762 2244 0 col\[2\].genblk1.mux4_I\[17\].x
rlabel metal1 98946 1530 98946 1530 0 col\[2\].genblk1.mux4_I\[18\].x
rlabel metal1 96692 2414 96692 2414 0 col\[2\].genblk1.mux4_I\[19\].x
rlabel metal2 117346 5916 117346 5916 0 col\[2\].genblk1.mux4_I\[1\].x
rlabel metal1 96370 3706 96370 3706 0 col\[2\].genblk1.mux4_I\[20\].x
rlabel metal2 94622 4284 94622 4284 0 col\[2\].genblk1.mux4_I\[21\].x
rlabel metal1 97336 5746 97336 5746 0 col\[2\].genblk1.mux4_I\[22\].x
rlabel metal1 94484 6222 94484 6222 0 col\[2\].genblk1.mux4_I\[23\].x
rlabel metal1 120566 3706 120566 3706 0 col\[2\].genblk1.mux4_I\[2\].x
rlabel metal1 120060 2074 120060 2074 0 col\[2\].genblk1.mux4_I\[3\].x
rlabel metal2 120106 3740 120106 3740 0 col\[2\].genblk1.mux4_I\[4\].x
rlabel metal2 119002 2244 119002 2244 0 col\[2\].genblk1.mux4_I\[5\].x
rlabel metal1 117162 1326 117162 1326 0 col\[2\].genblk1.mux4_I\[6\].x
rlabel metal2 111642 3876 111642 3876 0 col\[2\].genblk1.mux4_I\[7\].x
rlabel metal1 112378 3570 112378 3570 0 col\[2\].genblk1.mux4_I\[8\].x
rlabel metal1 111734 2958 111734 2958 0 col\[2\].genblk1.mux4_I\[9\].x
rlabel metal1 93058 3638 93058 3638 0 col\[2\].zbuf_bot_ena_I.e
rlabel via2 96462 2091 96462 2091 0 col\[2\].zbuf_bot_ena_I.z
rlabel metal1 98670 1292 98670 1292 0 col\[2\].zbuf_bot_iw_I\[0\].z
rlabel metal2 91678 1530 91678 1530 0 col\[2\].zbuf_bot_iw_I\[10\].z
rlabel metal1 91908 2074 91908 2074 0 col\[2\].zbuf_bot_iw_I\[11\].z
rlabel metal2 91126 2244 91126 2244 0 col\[2\].zbuf_bot_iw_I\[12\].z
rlabel metal1 90804 3026 90804 3026 0 col\[2\].zbuf_bot_iw_I\[13\].z
rlabel metal2 90298 2244 90298 2244 0 col\[2\].zbuf_bot_iw_I\[14\].z
rlabel metal1 89332 2074 89332 2074 0 col\[2\].zbuf_bot_iw_I\[15\].z
rlabel metal1 88964 1190 88964 1190 0 col\[2\].zbuf_bot_iw_I\[16\].z
rlabel metal1 88504 1326 88504 1326 0 col\[2\].zbuf_bot_iw_I\[17\].z
rlabel metal1 98854 1768 98854 1768 0 col\[2\].zbuf_bot_iw_I\[1\].z
rlabel metal1 95358 1258 95358 1258 0 col\[2\].zbuf_bot_iw_I\[2\].z
rlabel metal2 96462 3876 96462 3876 0 col\[2\].zbuf_bot_iw_I\[3\].z
rlabel metal1 94392 2074 94392 2074 0 col\[2\].zbuf_bot_iw_I\[4\].z
rlabel metal1 94116 1530 94116 1530 0 col\[2\].zbuf_bot_iw_I\[5\].z
rlabel metal1 93334 3060 93334 3060 0 col\[2\].zbuf_bot_iw_I\[6\].z
rlabel metal1 92736 1326 92736 1326 0 col\[2\].zbuf_bot_iw_I\[7\].z
rlabel metal1 93426 2074 93426 2074 0 col\[2\].zbuf_bot_iw_I\[8\].z
rlabel metal1 93472 1326 93472 1326 0 col\[2\].zbuf_bot_iw_I\[9\].z
rlabel metal2 94806 10200 94806 10200 0 col\[2\].zbuf_top_ena_I.e
rlabel metal1 100970 8058 100970 8058 0 col\[2\].zbuf_top_ena_I.z
rlabel metal2 100602 9350 100602 9350 0 col\[2\].zbuf_top_iw_I\[0\].z
rlabel metal1 93012 8602 93012 8602 0 col\[2\].zbuf_top_iw_I\[10\].z
rlabel metal1 91586 8908 91586 8908 0 col\[2\].zbuf_top_iw_I\[11\].z
rlabel metal1 91770 8602 91770 8602 0 col\[2\].zbuf_top_iw_I\[12\].z
rlabel metal2 90666 8636 90666 8636 0 col\[2\].zbuf_top_iw_I\[13\].z
rlabel metal1 90160 9146 90160 9146 0 col\[2\].zbuf_top_iw_I\[14\].z
rlabel metal2 90114 8058 90114 8058 0 col\[2\].zbuf_top_iw_I\[15\].z
rlabel metal1 88274 8908 88274 8908 0 col\[2\].zbuf_top_iw_I\[16\].z
rlabel metal2 88826 8908 88826 8908 0 col\[2\].zbuf_top_iw_I\[17\].z
rlabel metal2 99682 8636 99682 8636 0 col\[2\].zbuf_top_iw_I\[1\].z
rlabel metal2 98946 9350 98946 9350 0 col\[2\].zbuf_top_iw_I\[2\].z
rlabel metal2 98118 8704 98118 8704 0 col\[2\].zbuf_top_iw_I\[3\].z
rlabel metal1 97382 8534 97382 8534 0 col\[2\].zbuf_top_iw_I\[4\].z
rlabel metal2 96922 9078 96922 9078 0 col\[2\].zbuf_top_iw_I\[5\].z
rlabel metal2 96186 9078 96186 9078 0 col\[2\].zbuf_top_iw_I\[6\].z
rlabel metal2 94898 8636 94898 8636 0 col\[2\].zbuf_top_iw_I\[7\].z
rlabel metal2 94438 8636 94438 8636 0 col\[2\].zbuf_top_iw_I\[8\].z
rlabel metal2 93702 9350 93702 9350 0 col\[2\].zbuf_top_iw_I\[9\].z
rlabel metal1 121900 2414 121900 2414 0 col\[3\].zbuf_bot_ena_I.e
rlabel metal2 135378 2108 135378 2108 0 col\[3\].zbuf_bot_ena_I.z
rlabel metal2 134366 1530 134366 1530 0 col\[3\].zbuf_bot_iw_I\[0\].z
rlabel metal2 126730 2244 126730 2244 0 col\[3\].zbuf_bot_iw_I\[10\].z
rlabel metal1 126316 1530 126316 1530 0 col\[3\].zbuf_bot_iw_I\[11\].z
rlabel metal1 125626 1326 125626 1326 0 col\[3\].zbuf_bot_iw_I\[12\].z
rlabel metal1 124706 1326 124706 1326 0 col\[3\].zbuf_bot_iw_I\[13\].z
rlabel metal2 124338 2244 124338 2244 0 col\[3\].zbuf_bot_iw_I\[14\].z
rlabel metal2 123234 1530 123234 1530 0 col\[3\].zbuf_bot_iw_I\[15\].z
rlabel metal2 122498 1530 122498 1530 0 col\[3\].zbuf_bot_iw_I\[16\].z
rlabel metal2 121670 1530 121670 1530 0 col\[3\].zbuf_bot_iw_I\[17\].z
rlabel metal2 133722 2244 133722 2244 0 col\[3\].zbuf_bot_iw_I\[1\].z
rlabel metal2 133538 1938 133538 1938 0 col\[3\].zbuf_bot_iw_I\[2\].z
rlabel metal2 132710 1530 132710 1530 0 col\[3\].zbuf_bot_iw_I\[3\].z
rlabel metal2 131790 2210 131790 2210 0 col\[3\].zbuf_bot_iw_I\[4\].z
rlabel metal2 130686 1530 130686 1530 0 col\[3\].zbuf_bot_iw_I\[5\].z
rlabel metal1 130364 2414 130364 2414 0 col\[3\].zbuf_bot_iw_I\[6\].z
rlabel metal1 129168 1530 129168 1530 0 col\[3\].zbuf_bot_iw_I\[7\].z
rlabel metal2 128386 2244 128386 2244 0 col\[3\].zbuf_bot_iw_I\[8\].z
rlabel metal2 127650 1530 127650 1530 0 col\[3\].zbuf_bot_iw_I\[9\].z
rlabel metal1 128570 9044 128570 9044 0 col\[3\].zbuf_top_ena_I.e
rlabel metal2 134550 8772 134550 8772 0 col\[3\].zbuf_top_ena_I.z
rlabel metal2 134090 9350 134090 9350 0 col\[3\].zbuf_top_iw_I\[0\].z
rlabel metal2 126822 8636 126822 8636 0 col\[3\].zbuf_top_iw_I\[10\].z
rlabel metal2 126270 9350 126270 9350 0 col\[3\].zbuf_top_iw_I\[11\].z
rlabel metal2 125442 8636 125442 8636 0 col\[3\].zbuf_top_iw_I\[12\].z
rlabel metal2 124430 9350 124430 9350 0 col\[3\].zbuf_top_iw_I\[13\].z
rlabel metal2 123878 8636 123878 8636 0 col\[3\].zbuf_top_iw_I\[14\].z
rlabel metal2 123050 8636 123050 8636 0 col\[3\].zbuf_top_iw_I\[15\].z
rlabel metal2 122222 8636 122222 8636 0 col\[3\].zbuf_top_iw_I\[16\].z
rlabel metal2 121670 9078 121670 9078 0 col\[3\].zbuf_top_iw_I\[17\].z
rlabel metal2 133078 9350 133078 9350 0 col\[3\].zbuf_top_iw_I\[1\].z
rlabel metal2 132802 8058 132802 8058 0 col\[3\].zbuf_top_iw_I\[2\].z
rlabel metal2 131974 8636 131974 8636 0 col\[3\].zbuf_top_iw_I\[3\].z
rlabel metal2 131422 9350 131422 9350 0 col\[3\].zbuf_top_iw_I\[4\].z
rlabel metal2 130594 9350 130594 9350 0 col\[3\].zbuf_top_iw_I\[5\].z
rlabel metal1 129996 8602 129996 8602 0 col\[3\].zbuf_top_iw_I\[6\].z
rlabel metal2 129122 8058 129122 8058 0 col\[3\].zbuf_top_iw_I\[7\].z
rlabel metal2 128110 8908 128110 8908 0 col\[3\].zbuf_top_iw_I\[8\].z
rlabel metal2 127558 8636 127558 8636 0 col\[3\].zbuf_top_iw_I\[9\].z
rlabel metal2 145130 7123 145130 7123 0 col\[4\].genblk1.mux4_I\[0\].x
rlabel metal1 150558 2958 150558 2958 0 col\[4\].genblk1.mux4_I\[10\].x
rlabel metal1 152628 2074 152628 2074 0 col\[4\].genblk1.mux4_I\[11\].x
rlabel metal1 150512 1326 150512 1326 0 col\[4\].genblk1.mux4_I\[12\].x
rlabel metal1 149224 2074 149224 2074 0 col\[4\].genblk1.mux4_I\[13\].x
rlabel metal2 147522 4692 147522 4692 0 col\[4\].genblk1.mux4_I\[14\].x
rlabel metal1 145406 3434 145406 3434 0 col\[4\].genblk1.mux4_I\[15\].x
rlabel metal1 147476 2074 147476 2074 0 col\[4\].genblk1.mux4_I\[16\].x
rlabel metal1 145176 1530 145176 1530 0 col\[4\].genblk1.mux4_I\[17\].x
rlabel metal1 143796 2890 143796 2890 0 col\[4\].genblk1.mux4_I\[18\].x
rlabel metal2 142186 1972 142186 1972 0 col\[4\].genblk1.mux4_I\[19\].x
rlabel metal2 168130 4964 168130 4964 0 col\[4\].genblk1.mux4_I\[1\].x
rlabel metal1 142738 3502 142738 3502 0 col\[4\].genblk1.mux4_I\[20\].x
rlabel metal1 140852 2958 140852 2958 0 col\[4\].genblk1.mux4_I\[21\].x
rlabel metal1 140530 4012 140530 4012 0 col\[4\].genblk1.mux4_I\[22\].x
rlabel metal2 139610 3757 139610 3757 0 col\[4\].genblk1.mux4_I\[23\].x
rlabel metal1 158286 4012 158286 4012 0 col\[4\].genblk1.mux4_I\[2\].x
rlabel metal2 156170 3196 156170 3196 0 col\[4\].genblk1.mux4_I\[3\].x
rlabel metal2 155986 5406 155986 5406 0 col\[4\].genblk1.mux4_I\[4\].x
rlabel metal1 155388 4250 155388 4250 0 col\[4\].genblk1.mux4_I\[5\].x
rlabel metal2 155250 3876 155250 3876 0 col\[4\].genblk1.mux4_I\[6\].x
rlabel metal1 153134 4658 153134 4658 0 col\[4\].genblk1.mux4_I\[7\].x
rlabel metal1 152996 5134 152996 5134 0 col\[4\].genblk1.mux4_I\[8\].x
rlabel metal2 150834 4284 150834 4284 0 col\[4\].genblk1.mux4_I\[9\].x
rlabel viali 168866 2415 168866 2415 0 col\[4\].zbuf_bot_ena_I.e
rlabel metal1 168544 1326 168544 1326 0 col\[4\].zbuf_bot_ena_I.z
rlabel metal1 168544 1938 168544 1938 0 col\[4\].zbuf_bot_iw_I\[0\].z
rlabel metal1 161322 1326 161322 1326 0 col\[4\].zbuf_bot_iw_I\[10\].z
rlabel metal1 160448 2414 160448 2414 0 col\[4\].zbuf_bot_iw_I\[11\].z
rlabel metal1 159988 1326 159988 1326 0 col\[4\].zbuf_bot_iw_I\[12\].z
rlabel metal1 159758 3026 159758 3026 0 col\[4\].zbuf_bot_iw_I\[13\].z
rlabel metal1 159298 2074 159298 2074 0 col\[4\].zbuf_bot_iw_I\[14\].z
rlabel metal1 158332 1258 158332 1258 0 col\[4\].zbuf_bot_iw_I\[15\].z
rlabel metal2 155618 1836 155618 1836 0 col\[4\].zbuf_bot_iw_I\[16\].z
rlabel metal1 156584 1530 156584 1530 0 col\[4\].zbuf_bot_iw_I\[17\].z
rlabel metal1 167532 1326 167532 1326 0 col\[4\].zbuf_bot_iw_I\[1\].z
rlabel metal2 167486 2244 167486 2244 0 col\[4\].zbuf_bot_iw_I\[2\].z
rlabel metal1 166244 2074 166244 2074 0 col\[4\].zbuf_bot_iw_I\[3\].z
rlabel metal2 165646 2244 165646 2244 0 col\[4\].zbuf_bot_iw_I\[4\].z
rlabel metal2 164450 1530 164450 1530 0 col\[4\].zbuf_bot_iw_I\[5\].z
rlabel metal2 163990 2244 163990 2244 0 col\[4\].zbuf_bot_iw_I\[6\].z
rlabel metal1 163392 1326 163392 1326 0 col\[4\].zbuf_bot_iw_I\[7\].z
rlabel metal1 162380 1326 162380 1326 0 col\[4\].zbuf_bot_iw_I\[8\].z
rlabel metal1 161920 2074 161920 2074 0 col\[4\].zbuf_bot_iw_I\[9\].z
rlabel metal1 168636 7514 168636 7514 0 col\[4\].zbuf_top_ena_I.e
rlabel metal2 169234 8772 169234 8772 0 col\[4\].zbuf_top_ena_I.z
rlabel metal1 168636 7990 168636 7990 0 col\[4\].zbuf_top_iw_I\[0\].z
rlabel metal2 161506 8092 161506 8092 0 col\[4\].zbuf_top_iw_I\[10\].z
rlabel metal2 160770 8058 160770 8058 0 col\[4\].zbuf_top_iw_I\[11\].z
rlabel metal2 160034 8602 160034 8602 0 col\[4\].zbuf_top_iw_I\[12\].z
rlabel metal2 159298 8092 159298 8092 0 col\[4\].zbuf_top_iw_I\[13\].z
rlabel metal2 158562 8602 158562 8602 0 col\[4\].zbuf_top_iw_I\[14\].z
rlabel metal2 157090 8058 157090 8058 0 col\[4\].zbuf_top_iw_I\[15\].z
rlabel metal2 157366 9282 157366 9282 0 col\[4\].zbuf_top_iw_I\[16\].z
rlabel metal2 155986 8636 155986 8636 0 col\[4\].zbuf_top_iw_I\[17\].z
rlabel metal1 168268 9554 168268 9554 0 col\[4\].zbuf_top_iw_I\[1\].z
rlabel metal2 166750 8364 166750 8364 0 col\[4\].zbuf_top_iw_I\[2\].z
rlabel metal1 166606 7854 166606 7854 0 col\[4\].zbuf_top_iw_I\[3\].z
rlabel metal2 165922 8602 165922 8602 0 col\[4\].zbuf_top_iw_I\[4\].z
rlabel metal2 165186 8602 165186 8602 0 col\[4\].zbuf_top_iw_I\[5\].z
rlabel metal2 164450 8602 164450 8602 0 col\[4\].zbuf_top_iw_I\[6\].z
rlabel metal2 163714 8602 163714 8602 0 col\[4\].zbuf_top_iw_I\[7\].z
rlabel metal2 162978 8364 162978 8364 0 col\[4\].zbuf_top_iw_I\[8\].z
rlabel metal2 162242 8602 162242 8602 0 col\[4\].zbuf_top_iw_I\[9\].z
rlabel metal2 191222 2074 191222 2074 0 col\[5\].zbuf_bot_ena_I.e
rlabel metal1 203688 2414 203688 2414 0 col\[5\].zbuf_bot_ena_I.z
rlabel metal1 203504 1326 203504 1326 0 col\[5\].zbuf_bot_iw_I\[0\].z
rlabel metal1 195776 1326 195776 1326 0 col\[5\].zbuf_bot_iw_I\[10\].z
rlabel metal2 195730 2176 195730 2176 0 col\[5\].zbuf_bot_iw_I\[11\].z
rlabel metal2 194626 1530 194626 1530 0 col\[5\].zbuf_bot_iw_I\[12\].z
rlabel metal1 193614 1326 193614 1326 0 col\[5\].zbuf_bot_iw_I\[13\].z
rlabel metal1 192418 1292 192418 1292 0 col\[5\].zbuf_bot_iw_I\[14\].z
rlabel metal2 192234 2244 192234 2244 0 col\[5\].zbuf_bot_iw_I\[15\].z
rlabel metal2 191314 2176 191314 2176 0 col\[5\].zbuf_bot_iw_I\[16\].z
rlabel metal2 190946 2244 190946 2244 0 col\[5\].zbuf_bot_iw_I\[17\].z
rlabel metal1 203780 1938 203780 1938 0 col\[5\].zbuf_bot_iw_I\[1\].z
rlabel metal2 202722 2210 202722 2210 0 col\[5\].zbuf_bot_iw_I\[2\].z
rlabel metal1 201388 1258 201388 1258 0 col\[5\].zbuf_bot_iw_I\[3\].z
rlabel metal1 200836 2006 200836 2006 0 col\[5\].zbuf_bot_iw_I\[4\].z
rlabel metal2 200606 1530 200606 1530 0 col\[5\].zbuf_bot_iw_I\[5\].z
rlabel metal2 199778 2244 199778 2244 0 col\[5\].zbuf_bot_iw_I\[6\].z
rlabel metal2 198306 1938 198306 1938 0 col\[5\].zbuf_bot_iw_I\[7\].z
rlabel metal2 197570 2244 197570 2244 0 col\[5\].zbuf_bot_iw_I\[8\].z
rlabel metal1 196420 1462 196420 1462 0 col\[5\].zbuf_bot_iw_I\[9\].z
rlabel metal2 190854 9282 190854 9282 0 col\[5\].zbuf_top_ena_I.e
rlabel metal2 203550 8704 203550 8704 0 col\[5\].zbuf_top_ena_I.z
rlabel metal2 203458 9350 203458 9350 0 col\[5\].zbuf_top_iw_I\[0\].z
rlabel metal2 195638 9010 195638 9010 0 col\[5\].zbuf_top_iw_I\[10\].z
rlabel metal1 195224 9146 195224 9146 0 col\[5\].zbuf_top_iw_I\[11\].z
rlabel metal2 193890 8636 193890 8636 0 col\[5\].zbuf_top_iw_I\[12\].z
rlabel metal2 193154 8636 193154 8636 0 col\[5\].zbuf_top_iw_I\[13\].z
rlabel metal2 192694 9010 192694 9010 0 col\[5\].zbuf_top_iw_I\[14\].z
rlabel metal1 192418 9146 192418 9146 0 col\[5\].zbuf_top_iw_I\[15\].z
rlabel metal1 191544 8466 191544 8466 0 col\[5\].zbuf_top_iw_I\[16\].z
rlabel metal2 190394 8636 190394 8636 0 col\[5\].zbuf_top_iw_I\[17\].z
rlabel metal2 202722 9010 202722 9010 0 col\[5\].zbuf_top_iw_I\[1\].z
rlabel metal1 201618 8466 201618 8466 0 col\[5\].zbuf_top_iw_I\[2\].z
rlabel metal1 200836 8466 200836 8466 0 col\[5\].zbuf_top_iw_I\[3\].z
rlabel metal1 200008 8466 200008 8466 0 col\[5\].zbuf_top_iw_I\[4\].z
rlabel metal1 199134 8466 199134 8466 0 col\[5\].zbuf_top_iw_I\[5\].z
rlabel metal2 198582 8704 198582 8704 0 col\[5\].zbuf_top_iw_I\[6\].z
rlabel metal1 198076 9554 198076 9554 0 col\[5\].zbuf_top_iw_I\[7\].z
rlabel metal2 197570 9010 197570 9010 0 col\[5\].zbuf_top_iw_I\[8\].z
rlabel metal2 196098 8636 196098 8636 0 col\[5\].zbuf_top_iw_I\[9\].z
rlabel metal2 227102 5848 227102 5848 0 col\[6\].genblk1.mux4_I\[0\].x
rlabel metal1 219328 2618 219328 2618 0 col\[6\].genblk1.mux4_I\[10\].x
rlabel metal1 221674 2074 221674 2074 0 col\[6\].genblk1.mux4_I\[11\].x
rlabel metal2 219650 2176 219650 2176 0 col\[6\].genblk1.mux4_I\[12\].x
rlabel metal2 214958 1972 214958 1972 0 col\[6\].genblk1.mux4_I\[13\].x
rlabel metal2 213210 4046 213210 4046 0 col\[6\].genblk1.mux4_I\[14\].x
rlabel metal1 214958 4590 214958 4590 0 col\[6\].genblk1.mux4_I\[15\].x
rlabel metal1 212934 2924 212934 2924 0 col\[6\].genblk1.mux4_I\[16\].x
rlabel metal1 213348 1190 213348 1190 0 col\[6\].genblk1.mux4_I\[17\].x
rlabel metal2 214498 2142 214498 2142 0 col\[6\].genblk1.mux4_I\[18\].x
rlabel metal1 210841 1190 210841 1190 0 col\[6\].genblk1.mux4_I\[19\].x
rlabel metal2 222778 6052 222778 6052 0 col\[6\].genblk1.mux4_I\[1\].x
rlabel metal1 210312 3162 210312 3162 0 col\[6\].genblk1.mux4_I\[20\].x
rlabel metal1 208196 3706 208196 3706 0 col\[6\].genblk1.mux4_I\[21\].x
rlabel metal2 207322 5882 207322 5882 0 col\[6\].genblk1.mux4_I\[22\].x
rlabel metal2 206494 4828 206494 4828 0 col\[6\].genblk1.mux4_I\[23\].x
rlabel metal2 225262 4114 225262 4114 0 col\[6\].genblk1.mux4_I\[2\].x
rlabel metal2 227378 3808 227378 3808 0 col\[6\].genblk1.mux4_I\[3\].x
rlabel metal2 224802 4352 224802 4352 0 col\[6\].genblk1.mux4_I\[4\].x
rlabel metal2 222962 4964 222962 4964 0 col\[6\].genblk1.mux4_I\[5\].x
rlabel metal2 221122 3740 221122 3740 0 col\[6\].genblk1.mux4_I\[6\].x
rlabel metal2 220202 5644 220202 5644 0 col\[6\].genblk1.mux4_I\[7\].x
rlabel metal2 217994 4828 217994 4828 0 col\[6\].genblk1.mux4_I\[8\].x
rlabel metal2 217442 3740 217442 3740 0 col\[6\].genblk1.mux4_I\[9\].x
rlabel metal1 224112 1326 224112 1326 0 col\[6\].zbuf_bot_ena_I.e
rlabel metal1 237406 1972 237406 1972 0 col\[6\].zbuf_bot_ena_I.z
rlabel metal2 236946 2244 236946 2244 0 col\[6\].zbuf_bot_iw_I\[0\].z
rlabel metal1 229724 1326 229724 1326 0 col\[6\].zbuf_bot_iw_I\[10\].z
rlabel metal2 228574 1530 228574 1530 0 col\[6\].zbuf_bot_iw_I\[11\].z
rlabel metal2 228482 2244 228482 2244 0 col\[6\].zbuf_bot_iw_I\[12\].z
rlabel metal2 227286 1666 227286 1666 0 col\[6\].zbuf_bot_iw_I\[13\].z
rlabel metal2 226826 2244 226826 2244 0 col\[6\].zbuf_bot_iw_I\[14\].z
rlabel metal2 225814 2244 225814 2244 0 col\[6\].zbuf_bot_iw_I\[15\].z
rlabel metal2 225538 1530 225538 1530 0 col\[6\].zbuf_bot_iw_I\[16\].z
rlabel metal2 224158 2244 224158 2244 0 col\[6\].zbuf_bot_iw_I\[17\].z
rlabel metal1 236440 1326 236440 1326 0 col\[6\].zbuf_bot_iw_I\[1\].z
rlabel metal1 235566 2074 235566 2074 0 col\[6\].zbuf_bot_iw_I\[2\].z
rlabel metal1 234876 1326 234876 1326 0 col\[6\].zbuf_bot_iw_I\[3\].z
rlabel metal2 233726 1530 233726 1530 0 col\[6\].zbuf_bot_iw_I\[4\].z
rlabel metal1 233312 2074 233312 2074 0 col\[6\].zbuf_bot_iw_I\[5\].z
rlabel metal2 232622 2244 232622 2244 0 col\[6\].zbuf_bot_iw_I\[6\].z
rlabel metal1 231932 1326 231932 1326 0 col\[6\].zbuf_bot_iw_I\[7\].z
rlabel metal2 231794 2244 231794 2244 0 col\[6\].zbuf_bot_iw_I\[8\].z
rlabel metal2 230966 2244 230966 2244 0 col\[6\].zbuf_bot_iw_I\[9\].z
rlabel metal1 222594 8466 222594 8466 0 col\[6\].zbuf_top_ena_I.e
rlabel metal1 235796 8466 235796 8466 0 col\[6\].zbuf_top_ena_I.z
rlabel metal1 236440 8942 236440 8942 0 col\[6\].zbuf_top_iw_I\[0\].z
rlabel metal2 229034 8636 229034 8636 0 col\[6\].zbuf_top_iw_I\[10\].z
rlabel metal2 228482 9078 228482 9078 0 col\[6\].zbuf_top_iw_I\[11\].z
rlabel metal2 228390 9350 228390 9350 0 col\[6\].zbuf_top_iw_I\[12\].z
rlabel metal2 226826 8636 226826 8636 0 col\[6\].zbuf_top_iw_I\[13\].z
rlabel metal2 226090 8636 226090 8636 0 col\[6\].zbuf_top_iw_I\[14\].z
rlabel metal2 225354 8636 225354 8636 0 col\[6\].zbuf_top_iw_I\[15\].z
rlabel metal2 224526 8636 224526 8636 0 col\[6\].zbuf_top_iw_I\[16\].z
rlabel metal2 223790 9316 223790 9316 0 col\[6\].zbuf_top_iw_I\[17\].z
rlabel metal1 235428 9554 235428 9554 0 col\[6\].zbuf_top_iw_I\[1\].z
rlabel metal2 234738 8330 234738 8330 0 col\[6\].zbuf_top_iw_I\[2\].z
rlabel metal1 234048 8466 234048 8466 0 col\[6\].zbuf_top_iw_I\[3\].z
rlabel metal2 234002 9350 234002 9350 0 col\[6\].zbuf_top_iw_I\[4\].z
rlabel metal2 232438 8636 232438 8636 0 col\[6\].zbuf_top_iw_I\[5\].z
rlabel metal2 232346 9248 232346 9248 0 col\[6\].zbuf_top_iw_I\[6\].z
rlabel metal2 231518 8908 231518 8908 0 col\[6\].zbuf_top_iw_I\[7\].z
rlabel metal1 230552 8466 230552 8466 0 col\[6\].zbuf_top_iw_I\[8\].z
rlabel metal2 230046 9248 230046 9248 0 col\[6\].zbuf_top_iw_I\[9\].z
rlabel metal1 264086 2448 264086 2448 0 col\[7\].zbuf_bot_ena_I.e
rlabel metal1 270020 2618 270020 2618 0 col\[7\].zbuf_bot_ena_I.z
rlabel metal1 269882 1326 269882 1326 0 col\[7\].zbuf_bot_iw_I\[0\].z
rlabel metal1 263258 2074 263258 2074 0 col\[7\].zbuf_bot_iw_I\[10\].z
rlabel metal2 263166 1530 263166 1530 0 col\[7\].zbuf_bot_iw_I\[11\].z
rlabel metal1 262200 2414 262200 2414 0 col\[7\].zbuf_bot_iw_I\[12\].z
rlabel metal1 262200 1326 262200 1326 0 col\[7\].zbuf_bot_iw_I\[13\].z
rlabel metal1 261878 2992 261878 2992 0 col\[7\].zbuf_bot_iw_I\[14\].z
rlabel metal1 261418 2074 261418 2074 0 col\[7\].zbuf_bot_iw_I\[15\].z
rlabel metal1 260544 3502 260544 3502 0 col\[7\].zbuf_bot_iw_I\[16\].z
rlabel metal2 255622 1173 255622 1173 0 col\[7\].zbuf_bot_iw_I\[17\].z
rlabel metal2 270158 1802 270158 1802 0 col\[7\].zbuf_bot_iw_I\[1\].z
rlabel metal1 269928 1938 269928 1938 0 col\[7\].zbuf_bot_iw_I\[2\].z
rlabel metal2 268226 1530 268226 1530 0 col\[7\].zbuf_bot_iw_I\[3\].z
rlabel metal1 267674 1326 267674 1326 0 col\[7\].zbuf_bot_iw_I\[4\].z
rlabel metal2 267030 2176 267030 2176 0 col\[7\].zbuf_bot_iw_I\[5\].z
rlabel metal2 266754 1530 266754 1530 0 col\[7\].zbuf_bot_iw_I\[6\].z
rlabel metal2 265650 1530 265650 1530 0 col\[7\].zbuf_bot_iw_I\[7\].z
rlabel metal2 264914 1802 264914 1802 0 col\[7\].zbuf_bot_iw_I\[8\].z
rlabel metal2 264178 1530 264178 1530 0 col\[7\].zbuf_bot_iw_I\[9\].z
rlabel metal2 263902 8738 263902 8738 0 col\[7\].zbuf_top_ena_I.e
rlabel metal1 270250 3502 270250 3502 0 col\[7\].zbuf_top_ena_I.z
rlabel metal1 270480 4114 270480 4114 0 col\[7\].zbuf_top_iw_I\[0\].z
rlabel metal2 263166 8330 263166 8330 0 col\[7\].zbuf_top_iw_I\[10\].z
rlabel metal2 262338 8602 262338 8602 0 col\[7\].zbuf_top_iw_I\[11\].z
rlabel metal1 261832 8466 261832 8466 0 col\[7\].zbuf_top_iw_I\[12\].z
rlabel metal2 261602 8602 261602 8602 0 col\[7\].zbuf_top_iw_I\[13\].z
rlabel metal2 260314 8636 260314 8636 0 col\[7\].zbuf_top_iw_I\[14\].z
rlabel metal2 259762 8636 259762 8636 0 col\[7\].zbuf_top_iw_I\[15\].z
rlabel metal2 259394 9350 259394 9350 0 col\[7\].zbuf_top_iw_I\[16\].z
rlabel metal2 258106 8908 258106 8908 0 col\[7\].zbuf_top_iw_I\[17\].z
rlabel metal1 270802 4590 270802 4590 0 col\[7\].zbuf_top_iw_I\[1\].z
rlabel metal2 269330 6256 269330 6256 0 col\[7\].zbuf_top_iw_I\[2\].z
rlabel metal1 270158 5678 270158 5678 0 col\[7\].zbuf_top_iw_I\[3\].z
rlabel metal1 266846 9350 266846 9350 0 col\[7\].zbuf_top_iw_I\[4\].z
rlabel metal2 265926 7650 265926 7650 0 col\[7\].zbuf_top_iw_I\[5\].z
rlabel via1 266021 7378 266021 7378 0 col\[7\].zbuf_top_iw_I\[6\].z
rlabel metal1 266110 9520 266110 9520 0 col\[7\].zbuf_top_iw_I\[7\].z
rlabel metal1 264592 7854 264592 7854 0 col\[7\].zbuf_top_iw_I\[8\].z
rlabel metal2 264178 8364 264178 8364 0 col\[7\].zbuf_top_iw_I\[9\].z
rlabel metal2 269882 8670 269882 8670 0 net1
rlabel metal1 270204 3162 270204 3162 0 net10
rlabel metal1 109894 7956 109894 7956 0 net100
rlabel metal1 38778 3434 38778 3434 0 net101
rlabel metal1 102856 1326 102856 1326 0 net102
rlabel viali 97969 1938 97969 1938 0 net103
rlabel metal2 97842 1088 97842 1088 0 net104
rlabel metal1 97152 2550 97152 2550 0 net105
rlabel metal2 95082 4811 95082 4811 0 net106
rlabel metal1 94438 4692 94438 4692 0 net107
rlabel metal2 95910 7446 95910 7446 0 net108
rlabel metal1 101430 6120 101430 6120 0 net109
rlabel metal2 270802 5746 270802 5746 0 net11
rlabel metal2 112838 7650 112838 7650 0 net110
rlabel via1 115966 6307 115966 6307 0 net111
rlabel metal2 41354 1462 41354 1462 0 net112
rlabel metal1 118956 3570 118956 3570 0 net113
rlabel metal2 118266 1700 118266 1700 0 net114
rlabel metal2 117990 6698 117990 6698 0 net115
rlabel metal2 115966 3995 115966 3995 0 net116
rlabel metal1 116196 9350 116196 9350 0 net117
rlabel metal2 110722 3723 110722 3723 0 net118
rlabel metal1 111550 1870 111550 1870 0 net119
rlabel metal1 270802 3400 270802 3400 0 net12
rlabel metal2 110722 1904 110722 1904 0 net120
rlabel metal2 113160 1326 113160 1326 0 net121
rlabel metal1 112700 9350 112700 9350 0 net122
rlabel metal2 5474 850 5474 850 0 net123
rlabel metal2 112194 7837 112194 7837 0 net124
rlabel metal1 110538 9418 110538 9418 0 net125
rlabel metal2 110630 9112 110630 9112 0 net126
rlabel metal2 108974 9214 108974 9214 0 net127
rlabel metal2 100694 1394 100694 1394 0 net128
rlabel via1 97851 1938 97851 1938 0 net129
rlabel metal1 269192 3706 269192 3706 0 net13
rlabel metal1 107594 9656 107594 9656 0 net130
rlabel metal2 95312 2482 95312 2482 0 net131
rlabel metal2 94898 5287 94898 5287 0 net132
rlabel metal1 92414 4658 92414 4658 0 net133
rlabel metal2 38410 2040 38410 2040 0 net134
rlabel metal1 96554 7208 96554 7208 0 net135
rlabel metal2 92690 6018 92690 6018 0 net136
rlabel metal1 158930 3366 158930 3366 0 net137
rlabel metal2 158562 3638 158562 3638 0 net138
rlabel metal1 155112 2822 155112 2822 0 net139
rlabel metal1 268594 3604 268594 3604 0 net14
rlabel metal1 154974 2618 154974 2618 0 net140
rlabel metal1 155020 2074 155020 2074 0 net141
rlabel metal1 153778 2278 153778 2278 0 net142
rlabel metal1 154192 2074 154192 2074 0 net143
rlabel metal2 154698 986 154698 986 0 net144
rlabel via2 4830 2499 4830 2499 0 net145
rlabel metal2 18078 3026 18078 3026 0 net146
rlabel metal1 153824 2074 153824 2074 0 net147
rlabel metal1 154008 1190 154008 1190 0 net148
rlabel metal1 152950 2074 152950 2074 0 net149
rlabel metal1 268226 3162 268226 3162 0 net15
rlabel metal1 152858 1190 152858 1190 0 net150
rlabel metal1 148442 1258 148442 1258 0 net151
rlabel metal1 151386 1530 151386 1530 0 net152
rlabel metal2 145866 3876 145866 3876 0 net153
rlabel metal2 150834 782 150834 782 0 net154
rlabel metal1 146694 1462 146694 1462 0 net155
rlabel metal1 143290 1258 143290 1258 0 net156
rlabel metal2 5566 2210 5566 2210 0 net157
rlabel metal1 145268 1190 145268 1190 0 net158
rlabel metal1 140530 1360 140530 1360 0 net159
rlabel metal1 252862 6324 252862 6324 0 net16
rlabel metal1 139840 1870 139840 1870 0 net160
rlabel metal1 139564 2074 139564 2074 0 net161
rlabel metal3 139564 4420 139564 4420 0 net162
rlabel metal1 138506 1190 138506 1190 0 net163
rlabel metal1 157228 5610 157228 5610 0 net164
rlabel metal1 155894 9554 155894 9554 0 net165
rlabel metal2 156538 6596 156538 6596 0 net166
rlabel metal1 155664 3502 155664 3502 0 net167
rlabel metal2 2898 884 2898 884 0 net168
rlabel metal1 153548 5746 153548 5746 0 net169
rlabel metal1 268088 3706 268088 3706 0 net17
rlabel metal2 153226 6766 153226 6766 0 net170
rlabel metal2 153410 4352 153410 4352 0 net171
rlabel metal1 150696 5678 150696 5678 0 net172
rlabel metal1 150696 5202 150696 5202 0 net173
rlabel metal1 148948 4658 148948 4658 0 net174
rlabel metal1 148350 3026 148350 3026 0 net175
rlabel metal1 150742 1938 150742 1938 0 net176
rlabel metal1 148166 1326 148166 1326 0 net177
rlabel metal1 147821 1938 147821 1938 0 net178
rlabel metal2 2070 1088 2070 1088 0 net179
rlabel metal1 265880 4794 265880 4794 0 net18
rlabel metal1 145222 4046 145222 4046 0 net180
rlabel metal1 144440 4658 144440 4658 0 net181
rlabel metal1 145452 1938 145452 1938 0 net182
rlabel metal2 143106 5338 143106 5338 0 net183
rlabel metal2 142784 6052 142784 6052 0 net184
rlabel metal1 140392 1326 140392 1326 0 net185
rlabel metal2 140530 5644 140530 5644 0 net186
rlabel metal1 139472 8806 139472 8806 0 net187
rlabel metal1 140484 4658 140484 4658 0 net188
rlabel metal1 138414 4658 138414 4658 0 net189
rlabel metal1 265052 5338 265052 5338 0 net19
rlabel metal1 1840 2074 1840 2074 0 net190
rlabel metal2 189750 2448 189750 2448 0 net191
rlabel metal1 188048 1190 188048 1190 0 net192
rlabel metal2 182114 2822 182114 2822 0 net193
rlabel metal1 184874 2482 184874 2482 0 net194
rlabel metal2 187174 2686 187174 2686 0 net195
rlabel metal2 187174 918 187174 918 0 net196
rlabel metal1 185058 2550 185058 2550 0 net197
rlabel metal2 184598 3468 184598 3468 0 net198
rlabel metal2 184598 816 184598 816 0 net199
rlabel metal1 269882 7378 269882 7378 0 net2
rlabel via2 267950 2805 267950 2805 0 net20
rlabel metal1 177307 2006 177307 2006 0 net200
rlabel metal2 18722 7718 18722 7718 0 net201
rlabel metal1 153272 2550 153272 2550 0 net202
rlabel metal1 182022 1836 182022 1836 0 net203
rlabel metal2 182022 680 182022 680 0 net204
rlabel metal2 172454 1394 172454 1394 0 net205
rlabel metal2 179446 2023 179446 2023 0 net206
rlabel metal2 179446 1156 179446 1156 0 net207
rlabel metal2 178158 1666 178158 1666 0 net208
rlabel metal2 176962 1972 176962 1972 0 net209
rlabel metal1 265466 3400 265466 3400 0 net21
rlabel metal2 176870 2091 176870 2091 0 net210
rlabel metal3 173972 408 173972 408 0 net211
rlabel metal2 18078 9758 18078 9758 0 net212
rlabel via2 174754 1853 174754 1853 0 net213
rlabel metal2 174294 765 174294 765 0 net214
rlabel metal1 171534 1938 171534 1938 0 net215
rlabel metal2 172546 850 172546 850 0 net216
rlabel metal2 189750 8330 189750 8330 0 net217
rlabel metal1 187404 9350 187404 9350 0 net218
rlabel metal1 187312 9418 187312 9418 0 net219
rlabel metal1 265006 4046 265006 4046 0 net22
rlabel metal1 180780 8330 180780 8330 0 net220
rlabel metal2 182114 8398 182114 8398 0 net221
rlabel metal1 186806 9486 186806 9486 0 net222
rlabel metal1 20746 8296 20746 8296 0 net223
rlabel metal2 185886 7701 185886 7701 0 net224
rlabel metal2 177698 8432 177698 8432 0 net225
rlabel metal1 180780 9112 180780 9112 0 net226
rlabel metal2 178434 7021 178434 7021 0 net227
rlabel metal2 182114 9792 182114 9792 0 net228
rlabel metal1 179262 9520 179262 9520 0 net229
rlabel metal2 265374 4930 265374 4930 0 net23
rlabel metal2 149178 2043 149178 2043 0 net230
rlabel metal2 180734 10064 180734 10064 0 net231
rlabel metal1 179446 9452 179446 9452 0 net232
rlabel metal2 178066 9996 178066 9996 0 net233
rlabel metal2 19182 8568 19182 8568 0 net234
rlabel metal2 177606 9962 177606 9962 0 net235
rlabel metal2 176870 9520 176870 9520 0 net236
rlabel metal2 152490 8840 152490 8840 0 net237
rlabel metal2 172730 6256 172730 6256 0 net238
rlabel metal2 175582 9894 175582 9894 0 net239
rlabel metal1 267674 2618 267674 2618 0 net24
rlabel metal2 174294 9690 174294 9690 0 net240
rlabel metal2 169694 9214 169694 9214 0 net241
rlabel metal2 171166 8449 171166 8449 0 net242
rlabel metal1 224710 4794 224710 4794 0 net243
rlabel metal2 227010 3400 227010 3400 0 net244
rlabel metal2 15594 7854 15594 7854 0 net245
rlabel metal1 223606 2890 223606 2890 0 net246
rlabel metal2 225722 3332 225722 3332 0 net247
rlabel metal2 226274 1088 226274 1088 0 net248
rlabel metal2 222134 4182 222134 4182 0 net249
rlabel metal2 267306 3604 267306 3604 0 net25
rlabel metal2 220294 4284 220294 4284 0 net250
rlabel metal1 222824 2074 222824 2074 0 net251
rlabel metal1 220156 3638 220156 3638 0 net252
rlabel metal1 217488 4114 217488 4114 0 net253
rlabel metal2 222962 884 222962 884 0 net254
rlabel metal1 220248 1938 220248 1938 0 net255
rlabel metal2 18446 8364 18446 8364 0 net256
rlabel metal2 17342 1122 17342 1122 0 net257
rlabel metal1 219972 1530 219972 1530 0 net258
rlabel metal1 215418 1258 215418 1258 0 net259
rlabel metal1 268456 2278 268456 2278 0 net26
rlabel metal2 213670 1105 213670 1105 0 net260
rlabel metal1 213716 3706 213716 3706 0 net261
rlabel metal1 214820 1870 214820 1870 0 net262
rlabel metal2 212658 952 212658 952 0 net263
rlabel metal1 212842 1836 212842 1836 0 net264
rlabel metal2 210266 1530 210266 1530 0 net265
rlabel metal1 208978 1190 208978 1190 0 net266
rlabel metal1 207874 1190 207874 1190 0 net267
rlabel metal2 13754 7786 13754 7786 0 net268
rlabel metal1 207506 1224 207506 1224 0 net269
rlabel metal2 252862 7276 252862 7276 0 net27
rlabel metal1 206770 1190 206770 1190 0 net270
rlabel metal2 225262 7786 225262 7786 0 net271
rlabel metal1 223054 5746 223054 5746 0 net272
rlabel metal2 223422 5916 223422 5916 0 net273
rlabel metal2 225446 8177 225446 8177 0 net274
rlabel metal1 222640 4114 222640 4114 0 net275
rlabel metal1 220754 4658 220754 4658 0 net276
rlabel metal1 219742 4046 219742 4046 0 net277
rlabel metal1 218638 6290 218638 6290 0 net278
rlabel metal2 13662 7548 13662 7548 0 net279
rlabel metal1 251758 7276 251758 7276 0 net28
rlabel metal1 217856 5202 217856 5202 0 net280
rlabel metal1 217764 4046 217764 4046 0 net281
rlabel metal1 217028 9350 217028 9350 0 net282
rlabel metal1 219834 1870 219834 1870 0 net283
rlabel metal1 215050 9350 215050 9350 0 net284
rlabel metal1 215142 1326 215142 1326 0 net285
rlabel metal1 213394 5202 213394 5202 0 net286
rlabel metal1 212750 4658 212750 4658 0 net287
rlabel metal1 214820 1938 214820 1938 0 net288
rlabel metal1 211922 9350 211922 9350 0 net289
rlabel metal2 251666 7038 251666 7038 0 net29
rlabel metal2 12926 7922 12926 7922 0 net290
rlabel metal1 211232 2006 211232 2006 0 net291
rlabel metal2 210082 5338 210082 5338 0 net292
rlabel metal1 208886 3026 208886 3026 0 net293
rlabel metal2 207046 6494 207046 6494 0 net294
rlabel metal1 207874 6290 207874 6290 0 net295
rlabel metal1 207184 5202 207184 5202 0 net296
rlabel metal1 258704 2346 258704 2346 0 net297
rlabel metal2 226090 5406 226090 5406 0 net298
rlabel metal1 225170 2924 225170 2924 0 net299
rlabel metal2 263718 6052 263718 6052 0 net3
rlabel metal1 252586 6222 252586 6222 0 net30
rlabel metal1 243823 714 243823 714 0 net300
rlabel metal2 16514 8704 16514 8704 0 net301
rlabel metal1 255162 2346 255162 2346 0 net302
rlabel metal2 246882 1530 246882 1530 0 net303
rlabel metal1 228114 3672 228114 3672 0 net304
rlabel metal1 253690 2482 253690 2482 0 net305
rlabel metal1 246100 1870 246100 1870 0 net306
rlabel metal1 225630 3128 225630 3128 0 net307
rlabel metal2 223054 408 223054 408 0 net308
rlabel metal1 244260 1768 244260 1768 0 net309
rlabel via2 267766 7939 267766 7939 0 net31
rlabel via2 251298 1853 251298 1853 0 net310
rlabel metal2 251574 884 251574 884 0 net311
rlabel metal2 20746 7582 20746 7582 0 net312
rlabel metal2 213210 5355 213210 5355 0 net313
rlabel metal1 213728 4658 213728 4658 0 net314
rlabel metal3 245364 2176 245364 2176 0 net315
rlabel metal2 213578 1088 213578 1088 0 net316
rlabel metal2 213670 2091 213670 2091 0 net317
rlabel via1 211106 1326 211106 1326 0 net318
rlabel metal1 237889 2074 237889 2074 0 net319
rlabel metal2 250010 7140 250010 7140 0 net32
rlabel metal2 243846 918 243846 918 0 net320
rlabel metal1 240511 2074 240511 2074 0 net321
rlabel metal2 241086 850 241086 850 0 net322
rlabel metal2 20838 7650 20838 7650 0 net323
rlabel metal2 248998 7803 248998 7803 0 net324
rlabel metal2 224066 6800 224066 6800 0 net325
rlabel metal2 227562 5984 227562 5984 0 net326
rlabel metal1 226366 3570 226366 3570 0 net327
rlabel metal2 255346 8432 255346 8432 0 net328
rlabel metal2 249090 8568 249090 8568 0 net329
rlabel metal1 270802 7344 270802 7344 0 net33
rlabel metal2 249090 3672 249090 3672 0 net330
rlabel metal2 249826 8602 249826 8602 0 net331
rlabel metal2 244950 7072 244950 7072 0 net332
rlabel metal2 229034 4828 229034 4828 0 net333
rlabel metal2 39238 5576 39238 5576 0 net334
rlabel metal2 229862 1734 229862 1734 0 net335
rlabel metal2 229770 7208 229770 7208 0 net336
rlabel metal2 228252 3604 228252 3604 0 net337
rlabel metal2 214682 1054 214682 1054 0 net338
rlabel metal2 214406 5287 214406 5287 0 net339
rlabel metal1 270618 6698 270618 6698 0 net34
rlabel metal2 213762 5797 213762 5797 0 net340
rlabel metal2 246330 6953 246330 6953 0 net341
rlabel metal2 213394 697 213394 697 0 net342
rlabel metal1 213992 1870 213992 1870 0 net343
rlabel metal2 211002 765 211002 765 0 net344
rlabel metal1 15341 9554 15341 9554 0 net345
rlabel metal1 210220 2958 210220 2958 0 net346
rlabel metal2 207966 4046 207966 4046 0 net347
rlabel metal2 209162 6375 209162 6375 0 net348
rlabel via2 208426 5117 208426 5117 0 net349
rlabel metal2 18722 952 18722 952 0 net35
rlabel metal2 38778 5712 38778 5712 0 net350
rlabel metal2 7682 9214 7682 9214 0 net351
rlabel metal2 15778 952 15778 952 0 net352
rlabel metal2 40986 2587 40986 2587 0 net353
rlabel metal1 39744 2006 39744 2006 0 net354
rlabel metal1 38916 2414 38916 2414 0 net355
rlabel metal1 36846 4148 36846 4148 0 net356
rlabel metal1 37582 3060 37582 3060 0 net357
rlabel metal2 36754 3706 36754 3706 0 net358
rlabel metal2 19366 7021 19366 7021 0 net359
rlabel metal2 117254 3689 117254 3689 0 net36
rlabel metal2 36478 6698 36478 6698 0 net360
rlabel metal1 52486 1190 52486 1190 0 net361
rlabel metal2 51934 2924 51934 2924 0 net362
rlabel metal1 37582 2040 37582 2040 0 net363
rlabel metal1 51152 1190 51152 1190 0 net364
rlabel metal1 50508 3366 50508 3366 0 net365
rlabel metal1 49588 1190 49588 1190 0 net366
rlabel metal1 48990 1224 48990 1224 0 net367
rlabel metal1 48116 1190 48116 1190 0 net368
rlabel metal1 46920 4454 46920 4454 0 net369
rlabel metal2 115230 1224 115230 1224 0 net37
rlabel metal1 46138 1190 46138 1190 0 net370
rlabel metal1 45586 1190 45586 1190 0 net371
rlabel metal1 44896 4454 44896 4454 0 net372
rlabel metal1 44482 1224 44482 1224 0 net373
rlabel metal2 15134 2941 15134 2941 0 net374
rlabel metal1 43516 1190 43516 1190 0 net375
rlabel metal1 42688 1190 42688 1190 0 net376
rlabel metal1 41768 1190 41768 1190 0 net377
rlabel metal1 41032 3366 41032 3366 0 net378
rlabel metal1 40434 1190 40434 1190 0 net379
rlabel metal2 92414 1173 92414 1173 0 net38
rlabel metal2 39330 1598 39330 1598 0 net380
rlabel metal1 38502 1190 38502 1190 0 net381
rlabel metal1 37950 1190 37950 1190 0 net382
rlabel metal1 37812 2074 37812 2074 0 net383
rlabel metal1 36570 1190 36570 1190 0 net384
rlabel metal2 14398 2567 14398 2567 0 net385
rlabel metal1 35834 5338 35834 5338 0 net386
rlabel metal1 35604 4454 35604 4454 0 net387
rlabel metal2 52302 7514 52302 7514 0 net388
rlabel metal2 51290 7276 51290 7276 0 net389
rlabel metal1 109986 3468 109986 3468 0 net39
rlabel metal2 51842 6766 51842 6766 0 net390
rlabel metal1 50646 3502 50646 3502 0 net391
rlabel metal1 48714 4114 48714 4114 0 net392
rlabel metal1 48484 3434 48484 3434 0 net393
rlabel metal1 48158 3026 48158 3026 0 net394
rlabel metal2 47058 6970 47058 6970 0 net395
rlabel metal2 13570 850 13570 850 0 net396
rlabel metal1 46092 5270 46092 5270 0 net397
rlabel metal2 45678 7514 45678 7514 0 net398
rlabel metal2 44758 6460 44758 6460 0 net399
rlabel metal1 265420 3910 265420 3910 0 net4
rlabel metal2 92322 1360 92322 1360 0 net40
rlabel metal1 43746 3502 43746 3502 0 net400
rlabel metal2 43286 6222 43286 6222 0 net401
rlabel metal1 42734 2414 42734 2414 0 net402
rlabel metal2 41814 6970 41814 6970 0 net403
rlabel metal2 41078 6426 41078 6426 0 net404
rlabel metal1 40572 9350 40572 9350 0 net405
rlabel metal1 39790 8806 39790 8806 0 net406
rlabel metal2 12834 3060 12834 3060 0 net407
rlabel metal1 38318 2414 38318 2414 0 net408
rlabel metal1 37950 4148 37950 4148 0 net409
rlabel metal2 109986 1020 109986 1020 0 net41
rlabel metal2 37950 6222 37950 6222 0 net410
rlabel metal2 36662 6426 36662 6426 0 net411
rlabel metal2 35834 7310 35834 7310 0 net412
rlabel metal1 35834 4590 35834 4590 0 net413
rlabel metal1 91494 3978 91494 3978 0 net414
rlabel metal1 86618 1938 86618 1938 0 net415
rlabel metal2 117806 1618 117806 1618 0 net416
rlabel via2 117714 1955 117714 1955 0 net417
rlabel metal2 35558 5304 35558 5304 0 net418
rlabel metal1 195638 8908 195638 8908 0 net419
rlabel metal2 112378 1241 112378 1241 0 net42
rlabel metal1 197846 9010 197846 9010 0 net420
rlabel metal1 196374 1972 196374 1972 0 net421
rlabel metal2 198398 1598 198398 1598 0 net422
rlabel metal1 161276 8466 161276 8466 0 net423
rlabel metal1 168038 7888 168038 7888 0 net424
rlabel metal1 134366 8500 134366 8500 0 net425
rlabel metal1 132894 8976 132894 8976 0 net426
rlabel metal2 122682 2108 122682 2108 0 net427
rlabel metal2 134366 2176 134366 2176 0 net428
rlabel metal1 94622 8942 94622 8942 0 net429
rlabel metal2 78982 1462 78982 1462 0 net43
rlabel metal2 100970 8126 100970 8126 0 net430
rlabel metal2 59938 9146 59938 9146 0 net431
rlabel metal1 64262 8976 64262 8976 0 net432
rlabel metal2 59846 2108 59846 2108 0 net433
rlabel metal1 60674 1904 60674 1904 0 net434
rlabel metal1 25760 8942 25760 8942 0 net435
rlabel metal1 32982 8432 32982 8432 0 net436
rlabel metal1 263626 8908 263626 8908 0 net437
rlabel metal1 267444 7854 267444 7854 0 net438
rlabel metal1 264362 1904 264362 1904 0 net439
rlabel metal2 77602 1088 77602 1088 0 net44
rlabel metal2 265190 2176 265190 2176 0 net440
rlabel metal2 232346 8449 232346 8449 0 net441
rlabel metal1 230552 8942 230552 8942 0 net442
rlabel metal1 157182 1360 157182 1360 0 net443
rlabel metal1 167302 1972 167302 1972 0 net444
rlabel metal2 93334 1241 93334 1241 0 net445
rlabel metal1 96324 1938 96324 1938 0 net446
rlabel metal2 26082 1904 26082 1904 0 net447
rlabel metal1 27140 1938 27140 1938 0 net448
rlabel metal2 230782 2244 230782 2244 0 net449
rlabel metal2 77510 1428 77510 1428 0 net45
rlabel metal1 233404 2346 233404 2346 0 net450
rlabel metal1 38272 2346 38272 2346 0 net451
rlabel metal2 43378 2754 43378 2754 0 net452
rlabel metal2 51382 4964 51382 4964 0 net453
rlabel metal1 105938 1394 105938 1394 0 net454
rlabel metal2 116334 6188 116334 6188 0 net455
rlabel metal2 105662 3298 105662 3298 0 net456
rlabel metal2 154606 3706 154606 3706 0 net457
rlabel metal2 137034 6188 137034 6188 0 net458
rlabel metal1 153870 6256 153870 6256 0 net459
rlabel metal2 14306 1054 14306 1054 0 net46
rlabel metal2 226458 6052 226458 6052 0 net460
rlabel metal1 216936 6766 216936 6766 0 net461
rlabel metal1 213440 1394 213440 1394 0 net462
rlabel metal2 137310 5423 137310 5423 0 net463
rlabel metal1 41315 2482 41315 2482 0 net464
rlabel metal1 43661 2482 43661 2482 0 net465
rlabel metal2 47150 4097 47150 4097 0 net466
rlabel metal1 94898 2550 94898 2550 0 net467
rlabel metal2 111366 1666 111366 1666 0 net468
rlabel metal1 116610 1802 116610 1802 0 net469
rlabel metal1 89838 2516 89838 2516 0 net47
rlabel metal1 148580 1870 148580 1870 0 net470
rlabel metal1 137126 6256 137126 6256 0 net471
rlabel metal1 154146 5746 154146 5746 0 net472
rlabel metal1 220570 1870 220570 1870 0 net473
rlabel metal2 214130 5236 214130 5236 0 net474
rlabel metal1 213348 1870 213348 1870 0 net475
rlabel metal1 109940 1938 109940 1938 0 net476
rlabel metal1 58742 1938 58742 1938 0 net477
rlabel metal1 264132 1938 264132 1938 0 net478
rlabel metal1 25116 1394 25116 1394 0 net479
rlabel metal1 77326 1938 77326 1938 0 net48
rlabel metal1 231150 1938 231150 1938 0 net480
rlabel metal1 25806 1394 25806 1394 0 net481
rlabel metal1 264730 1938 264730 1938 0 net482
rlabel metal1 27140 1394 27140 1394 0 net483
rlabel metal1 232162 1938 232162 1938 0 net484
rlabel metal1 62146 8466 62146 8466 0 net485
rlabel metal1 266616 1938 266616 1938 0 net486
rlabel metal1 62422 8908 62422 8908 0 net487
rlabel metal1 233864 1938 233864 1938 0 net488
rlabel metal1 29440 1870 29440 1870 0 net489
rlabel metal2 75026 1122 75026 1122 0 net49
rlabel metal3 267697 2108 267697 2108 0 net490
rlabel metal1 30084 1870 30084 1870 0 net491
rlabel metal1 235704 1938 235704 1938 0 net492
rlabel metal1 31188 1870 31188 1870 0 net493
rlabel metal1 235888 1394 235888 1394 0 net494
rlabel metal1 28980 1428 28980 1428 0 net495
rlabel metal1 192326 2040 192326 2040 0 net496
rlabel metal1 23736 1394 23736 1394 0 net497
rlabel metal1 191176 1394 191176 1394 0 net498
rlabel metal1 23000 1870 23000 1870 0 net499
rlabel metal1 268640 7854 268640 7854 0 net5
rlabel metal2 74106 816 74106 816 0 net50
rlabel metal2 191866 1921 191866 1921 0 net500
rlabel metal2 27646 1700 27646 1700 0 net501
rlabel metal2 192878 2210 192878 2210 0 net502
rlabel metal1 22540 2482 22540 2482 0 net503
rlabel metal1 193614 1938 193614 1938 0 net504
rlabel metal1 125258 1938 125258 1938 0 net505
rlabel metal1 194672 1870 194672 1870 0 net506
rlabel metal1 22770 1394 22770 1394 0 net507
rlabel metal2 195362 4419 195362 4419 0 net508
rlabel metal1 58972 1394 58972 1394 0 net509
rlabel metal1 94438 1462 94438 1462 0 net51
rlabel metal1 196098 1938 196098 1938 0 net510
rlabel metal1 32108 1870 32108 1870 0 net511
rlabel metal1 236348 1938 236348 1938 0 net512
rlabel metal2 267582 5100 267582 5100 0 net513
rlabel metal1 267122 6766 267122 6766 0 net514
rlabel metal1 265098 5576 265098 5576 0 net515
rlabel metal1 253092 6290 253092 6290 0 net516
rlabel metal3 272121 8772 272121 8772 0 net517
rlabel metal1 265834 4148 265834 4148 0 net518
rlabel metal3 272305 1020 272305 1020 0 net519
rlabel metal2 72818 918 72818 918 0 net52
rlabel metal4 828 1459 828 1459 0 net520
rlabel metal1 1610 9146 1610 9146 0 net521
rlabel metal4 34960 371 34960 371 0 net522
rlabel metal2 35190 9707 35190 9707 0 net523
rlabel metal4 69092 507 69092 507 0 net524
rlabel via2 69138 9571 69138 9571 0 net525
rlabel metal4 103224 235 103224 235 0 net526
rlabel metal2 103270 9911 103270 9911 0 net527
rlabel metal4 137356 779 137356 779 0 net528
rlabel metal4 137356 10169 137356 10169 0 net529
rlabel metal1 94116 3502 94116 3502 0 net53
rlabel metal4 171488 371 171488 371 0 net530
rlabel metal2 171718 9911 171718 9911 0 net531
rlabel metal4 205620 507 205620 507 0 net532
rlabel metal2 205850 9911 205850 9911 0 net533
rlabel metal4 239752 371 239752 371 0 net534
rlabel metal2 239982 9911 239982 9911 0 net535
rlabel metal1 32154 2958 32154 2958 0 net536
rlabel metal2 32890 8194 32890 8194 0 net537
rlabel metal2 66378 2448 66378 2448 0 net538
rlabel metal1 67344 7922 67344 7922 0 net539
rlabel metal2 81466 3162 81466 3162 0 net54
rlabel metal1 96002 1938 96002 1938 0 net540
rlabel metal1 101246 7922 101246 7922 0 net541
rlabel metal1 135010 2482 135010 2482 0 net542
rlabel metal2 134274 8194 134274 8194 0 net543
rlabel metal2 167946 2686 167946 2686 0 net544
rlabel metal1 169326 7922 169326 7922 0 net545
rlabel metal2 203182 2686 203182 2686 0 net546
rlabel metal2 202998 8126 202998 8126 0 net547
rlabel metal1 235796 2958 235796 2958 0 net548
rlabel metal2 235842 8058 235842 8058 0 net549
rlabel metal1 74382 1326 74382 1326 0 net55
rlabel metal1 269238 2482 269238 2482 0 net550
rlabel metal2 268594 6868 268594 6868 0 net551
rlabel metal1 265972 3570 265972 3570 0 net552
rlabel metal1 74198 1224 74198 1224 0 net56
rlabel metal2 10626 1088 10626 1088 0 net57
rlabel metal1 92690 9656 92690 9656 0 net58
rlabel metal2 115046 6375 115046 6375 0 net59
rlabel metal1 269514 8364 269514 8364 0 net6
rlabel metal2 117346 7905 117346 7905 0 net60
rlabel metal1 117484 1938 117484 1938 0 net61
rlabel metal2 117070 7004 117070 7004 0 net62
rlabel metal2 115046 2074 115046 2074 0 net63
rlabel metal2 114954 1105 114954 1105 0 net64
rlabel metal2 109434 5134 109434 5134 0 net65
rlabel metal1 110630 1938 110630 1938 0 net66
rlabel metal2 94530 7344 94530 7344 0 net67
rlabel metal1 25070 1972 25070 1972 0 net68
rlabel metal2 110354 1598 110354 1598 0 net69
rlabel metal2 263074 6392 263074 6392 0 net7
rlabel metal2 78982 7633 78982 7633 0 net70
rlabel metal2 77602 8772 77602 8772 0 net71
rlabel via2 94438 5525 94438 5525 0 net72
rlabel metal2 82754 7497 82754 7497 0 net73
rlabel metal2 75854 8585 75854 8585 0 net74
rlabel metal2 75026 8466 75026 8466 0 net75
rlabel metal2 74566 9452 74566 9452 0 net76
rlabel metal2 73738 8432 73738 8432 0 net77
rlabel metal1 78706 9554 78706 9554 0 net78
rlabel metal2 43378 2125 43378 2125 0 net79
rlabel metal1 265742 7752 265742 7752 0 net8
rlabel metal2 72358 7684 72358 7684 0 net80
rlabel metal1 79258 9384 79258 9384 0 net81
rlabel metal2 69874 10132 69874 10132 0 net82
rlabel metal2 91126 7548 91126 7548 0 net83
rlabel metal1 120934 1224 120934 1224 0 net84
rlabel metal1 120152 1530 120152 1530 0 net85
rlabel metal1 119048 1190 119048 1190 0 net86
rlabel metal2 118542 1700 118542 1700 0 net87
rlabel metal1 117944 1190 117944 1190 0 net88
rlabel via1 116070 1938 116070 1938 0 net89
rlabel metal2 268502 5423 268502 5423 0 net9
rlabel metal2 36570 4250 36570 4250 0 net90
rlabel metal1 116357 1394 116357 1394 0 net91
rlabel metal1 114034 2040 114034 2040 0 net92
rlabel metal1 112585 1870 112585 1870 0 net93
rlabel metal2 118174 1207 118174 1207 0 net94
rlabel metal2 113298 1122 113298 1122 0 net95
rlabel metal1 109066 952 109066 952 0 net96
rlabel metal1 111182 6834 111182 6834 0 net97
rlabel metal2 110998 1601 110998 1601 0 net98
rlabel metal2 107870 5712 107870 5712 0 net99
rlabel metal2 262338 7327 262338 7327 0 spine_iw[10]
rlabel metal2 263258 6953 263258 6953 0 spine_iw[11]
rlabel metal2 267950 7225 267950 7225 0 spine_iw[12]
rlabel metal3 270166 6868 270166 6868 0 spine_iw[13]
rlabel metal3 271684 6732 271684 6732 0 spine_iw[14]
rlabel metal3 272236 6596 272236 6596 0 spine_iw[15]
rlabel metal3 272144 6460 272144 6460 0 spine_iw[16]
rlabel metal3 271868 6324 271868 6324 0 spine_iw[17]
rlabel metal3 271477 6188 271477 6188 0 spine_iw[18]
rlabel metal3 272052 6052 272052 6052 0 spine_iw[19]
rlabel metal3 270350 8500 270350 8500 0 spine_iw[1]
rlabel metal3 271776 5916 271776 5916 0 spine_iw[20]
rlabel metal3 271661 5780 271661 5780 0 spine_iw[21]
rlabel metal3 271569 5644 271569 5644 0 spine_iw[22]
rlabel metal3 272098 5508 272098 5508 0 spine_iw[23]
rlabel metal3 272098 5372 272098 5372 0 spine_iw[24]
rlabel metal3 270718 5236 270718 5236 0 spine_iw[25]
rlabel metal3 270442 5100 270442 5100 0 spine_iw[26]
rlabel metal3 272190 4964 272190 4964 0 spine_iw[27]
rlabel metal3 270672 4828 270672 4828 0 spine_iw[28]
rlabel metal1 268088 2414 268088 2414 0 spine_iw[29]
rlabel metal3 270212 8364 270212 8364 0 spine_iw[2]
rlabel metal3 272213 8228 272213 8228 0 spine_iw[3]
rlabel metal3 272282 8092 272282 8092 0 spine_iw[4]
rlabel metal3 272282 7956 272282 7956 0 spine_iw[5]
rlabel metal3 268648 7820 268648 7820 0 spine_iw[6]
rlabel metal3 272098 7684 272098 7684 0 spine_iw[7]
rlabel metal3 272121 7548 272121 7548 0 spine_iw[8]
rlabel metal2 263994 7531 263994 7531 0 spine_iw[9]
rlabel metal3 270166 3060 270166 3060 0 spine_ow[10]
rlabel metal2 249642 3077 249642 3077 0 spine_ow[11]
rlabel metal3 252264 2992 252264 2992 0 spine_ow[12]
rlabel metal1 250654 2550 250654 2550 0 spine_ow[13]
rlabel metal3 270396 2516 270396 2516 0 spine_ow[14]
rlabel metal1 247618 3026 247618 3026 0 spine_ow[15]
rlabel metal2 246698 1785 246698 1785 0 spine_ow[16]
rlabel metal2 253138 1938 253138 1938 0 spine_ow[17]
rlabel metal3 272236 1972 272236 1972 0 spine_ow[18]
rlabel metal2 250562 1666 250562 1666 0 spine_ow[19]
rlabel metal2 252678 4709 252678 4709 0 spine_ow[1]
rlabel metal2 252402 2176 252402 2176 0 spine_ow[20]
rlabel metal3 272282 1564 272282 1564 0 spine_ow[21]
rlabel metal1 250700 4046 250700 4046 0 spine_ow[22]
rlabel metal3 272190 1292 272190 1292 0 spine_ow[23]
rlabel metal3 272121 1156 272121 1156 0 spine_ow[24]
rlabel metal3 272121 4148 272121 4148 0 spine_ow[2]
rlabel metal3 272213 4012 272213 4012 0 spine_ow[3]
rlabel metal3 272282 3876 272282 3876 0 spine_ow[4]
rlabel metal3 270212 3740 270212 3740 0 spine_ow[5]
rlabel metal2 263994 2176 263994 2176 0 spine_ow[6]
rlabel metal3 272213 3468 272213 3468 0 spine_ow[7]
rlabel metal3 272121 3332 272121 3332 0 spine_ow[8]
rlabel metal3 272098 3196 272098 3196 0 spine_ow[9]
rlabel metal4 32476 847 32476 847 0 um_ena[0]
rlabel metal4 203136 303 203136 303 0 um_ena[10]
rlabel metal2 204102 9707 204102 9707 0 um_ena[11]
rlabel metal4 237268 847 237268 847 0 um_ena[12]
rlabel via2 236302 8619 236302 8619 0 um_ena[13]
rlabel metal4 271400 371 271400 371 0 um_ena[14]
rlabel metal1 270388 3706 270388 3706 0 um_ena[15]
rlabel via2 33074 9163 33074 9163 0 um_ena[1]
rlabel metal4 66608 303 66608 303 0 um_ena[2]
rlabel metal2 67206 9537 67206 9537 0 um_ena[3]
rlabel via3 100763 3196 100763 3196 0 um_ena[4]
rlabel via2 101246 9163 101246 9163 0 um_ena[5]
rlabel metal4 134872 235 134872 235 0 um_ena[6]
rlabel metal2 134734 9707 134734 9707 0 um_ena[7]
rlabel metal4 169004 371 169004 371 0 um_ena[8]
rlabel metal1 169786 9452 169786 9452 0 um_ena[9]
rlabel metal4 31740 371 31740 371 0 um_iw[0]
rlabel via2 92782 9707 92782 9707 0 um_iw[100]
rlabel via2 91770 9163 91770 9163 0 um_iw[101]
rlabel metal1 91770 9486 91770 9486 0 um_iw[102]
rlabel via2 90850 8619 90850 8619 0 um_iw[103]
rlabel metal2 90390 9843 90390 9843 0 um_iw[104]
rlabel metal2 89746 7905 89746 7905 0 um_iw[105]
rlabel metal1 88366 9146 88366 9146 0 um_iw[106]
rlabel metal1 88274 8602 88274 8602 0 um_iw[107]
rlabel metal4 134136 371 134136 371 0 um_iw[108]
rlabel metal4 133400 235 133400 235 0 um_iw[109]
rlabel metal4 24380 711 24380 711 0 um_iw[10]
rlabel metal4 132664 235 132664 235 0 um_iw[110]
rlabel metal4 131928 235 131928 235 0 um_iw[111]
rlabel metal4 131192 371 131192 371 0 um_iw[112]
rlabel metal4 130456 371 130456 371 0 um_iw[113]
rlabel metal4 129720 235 129720 235 0 um_iw[114]
rlabel metal4 128984 371 128984 371 0 um_iw[115]
rlabel metal4 128248 235 128248 235 0 um_iw[116]
rlabel metal4 127512 303 127512 303 0 um_iw[117]
rlabel metal4 126776 235 126776 235 0 um_iw[118]
rlabel metal4 126040 371 126040 371 0 um_iw[119]
rlabel metal4 23644 711 23644 711 0 um_iw[11]
rlabel metal4 125304 371 125304 371 0 um_iw[120]
rlabel metal4 124568 371 124568 371 0 um_iw[121]
rlabel metal4 123832 235 123832 235 0 um_iw[122]
rlabel metal4 123096 303 123096 303 0 um_iw[123]
rlabel metal4 122360 303 122360 303 0 um_iw[124]
rlabel metal4 121624 303 121624 303 0 um_iw[125]
rlabel metal2 134182 9979 134182 9979 0 um_iw[126]
rlabel metal2 133446 9979 133446 9979 0 um_iw[127]
rlabel metal2 132986 9163 132986 9163 0 um_iw[128]
rlabel metal2 132158 9435 132158 9435 0 um_iw[129]
rlabel metal1 22448 2618 22448 2618 0 um_iw[12]
rlabel metal2 131514 9979 131514 9979 0 um_iw[130]
rlabel metal2 130778 9979 130778 9979 0 um_iw[131]
rlabel metal1 129628 9690 129628 9690 0 um_iw[132]
rlabel metal2 129306 9163 129306 9163 0 um_iw[133]
rlabel metal2 128294 9435 128294 9435 0 um_iw[134]
rlabel metal2 127742 9435 127742 9435 0 um_iw[135]
rlabel metal2 127006 9435 127006 9435 0 um_iw[136]
rlabel metal2 126362 9979 126362 9979 0 um_iw[137]
rlabel metal2 125626 9503 125626 9503 0 um_iw[138]
rlabel metal2 125258 9979 125258 9979 0 um_iw[139]
rlabel metal4 22172 915 22172 915 0 um_iw[13]
rlabel metal2 124062 9435 124062 9435 0 um_iw[140]
rlabel metal2 123234 9435 123234 9435 0 um_iw[141]
rlabel metal2 122406 9435 122406 9435 0 um_iw[142]
rlabel metal2 121762 9979 121762 9979 0 um_iw[143]
rlabel metal4 168268 779 168268 779 0 um_iw[144]
rlabel metal4 167532 235 167532 235 0 um_iw[145]
rlabel metal4 166796 643 166796 643 0 um_iw[146]
rlabel metal4 166060 643 166060 643 0 um_iw[147]
rlabel metal4 165324 643 165324 643 0 um_iw[148]
rlabel metal4 164588 371 164588 371 0 um_iw[149]
rlabel metal4 21436 371 21436 371 0 um_iw[14]
rlabel metal4 163852 643 163852 643 0 um_iw[150]
rlabel metal4 163116 371 163116 371 0 um_iw[151]
rlabel metal4 162380 371 162380 371 0 um_iw[152]
rlabel metal4 161644 643 161644 643 0 um_iw[153]
rlabel metal4 160908 235 160908 235 0 um_iw[154]
rlabel metal4 160172 643 160172 643 0 um_iw[155]
rlabel metal4 159436 371 159436 371 0 um_iw[156]
rlabel metal4 158700 643 158700 643 0 um_iw[157]
rlabel metal4 157964 711 157964 711 0 um_iw[158]
rlabel metal4 157228 779 157228 779 0 um_iw[159]
rlabel metal4 20700 779 20700 779 0 um_iw[15]
rlabel metal1 156124 2618 156124 2618 0 um_iw[160]
rlabel metal4 155756 779 155756 779 0 um_iw[161]
rlabel metal1 170016 9078 170016 9078 0 um_iw[162]
rlabel metal1 168728 9690 168728 9690 0 um_iw[163]
rlabel metal2 166934 7939 166934 7939 0 um_iw[164]
rlabel metal1 166704 7718 166704 7718 0 um_iw[165]
rlabel metal1 165738 8058 165738 8058 0 um_iw[166]
rlabel metal1 165324 7718 165324 7718 0 um_iw[167]
rlabel metal1 164312 8058 164312 8058 0 um_iw[168]
rlabel metal2 163898 8211 163898 8211 0 um_iw[169]
rlabel metal4 19964 847 19964 847 0 um_iw[16]
rlabel metal1 162794 7514 162794 7514 0 um_iw[170]
rlabel metal2 162426 8211 162426 8211 0 um_iw[171]
rlabel metal1 161368 8058 161368 8058 0 um_iw[172]
rlabel metal2 160954 8211 160954 8211 0 um_iw[173]
rlabel metal1 159850 8058 159850 8058 0 um_iw[174]
rlabel metal1 159436 7718 159436 7718 0 um_iw[175]
rlabel via2 158746 8075 158746 8075 0 um_iw[176]
rlabel metal2 157274 8211 157274 8211 0 um_iw[177]
rlabel via2 156722 9435 156722 9435 0 um_iw[178]
rlabel metal1 156124 8602 156124 8602 0 um_iw[179]
rlabel via3 19251 2788 19251 2788 0 um_iw[17]
rlabel metal4 202400 303 202400 303 0 um_iw[180]
rlabel metal4 201664 235 201664 235 0 um_iw[181]
rlabel metal4 200928 235 200928 235 0 um_iw[182]
rlabel metal4 200192 303 200192 303 0 um_iw[183]
rlabel metal4 199456 235 199456 235 0 um_iw[184]
rlabel metal4 198720 303 198720 303 0 um_iw[185]
rlabel metal4 197984 235 197984 235 0 um_iw[186]
rlabel metal4 197248 235 197248 235 0 um_iw[187]
rlabel metal4 196512 303 196512 303 0 um_iw[188]
rlabel metal4 195776 235 195776 235 0 um_iw[189]
rlabel metal2 32522 9979 32522 9979 0 um_iw[18]
rlabel metal4 195040 303 195040 303 0 um_iw[190]
rlabel metal4 194304 235 194304 235 0 um_iw[191]
rlabel metal4 193568 303 193568 303 0 um_iw[192]
rlabel metal4 192832 303 192832 303 0 um_iw[193]
rlabel metal4 192096 235 192096 235 0 um_iw[194]
rlabel metal4 191360 235 191360 235 0 um_iw[195]
rlabel metal4 190624 303 190624 303 0 um_iw[196]
rlabel metal1 190532 2618 190532 2618 0 um_iw[197]
rlabel metal1 202860 9350 202860 9350 0 um_iw[198]
rlabel metal2 202538 9843 202538 9843 0 um_iw[199]
rlabel via2 31050 8619 31050 8619 0 um_iw[19]
rlabel metal4 31004 371 31004 371 0 um_iw[1]
rlabel metal1 201250 8330 201250 8330 0 um_iw[200]
rlabel metal2 200790 9299 200790 9299 0 um_iw[201]
rlabel metal2 199962 9299 199962 9299 0 um_iw[202]
rlabel metal1 199180 8330 199180 8330 0 um_iw[203]
rlabel metal1 198582 9146 198582 9146 0 um_iw[204]
rlabel metal1 197892 9418 197892 9418 0 um_iw[205]
rlabel metal2 196558 9843 196558 9843 0 um_iw[206]
rlabel metal2 195822 9299 195822 9299 0 um_iw[207]
rlabel metal2 195546 9843 195546 9843 0 um_iw[208]
rlabel metal1 194580 9418 194580 9418 0 um_iw[209]
rlabel metal1 30360 9690 30360 9690 0 um_iw[20]
rlabel metal2 194074 9299 194074 9299 0 um_iw[210]
rlabel metal1 193108 8330 193108 8330 0 um_iw[211]
rlabel metal2 192970 9843 192970 9843 0 um_iw[212]
rlabel metal1 191820 9418 191820 9418 0 um_iw[213]
rlabel metal2 191314 9367 191314 9367 0 um_iw[214]
rlabel metal4 189888 10509 189888 10509 0 um_iw[215]
rlabel metal4 236532 643 236532 643 0 um_iw[216]
rlabel metal4 235796 371 235796 371 0 um_iw[217]
rlabel metal4 235060 643 235060 643 0 um_iw[218]
rlabel metal4 234324 371 234324 371 0 um_iw[219]
rlabel via2 29118 9707 29118 9707 0 um_iw[21]
rlabel metal4 233588 371 233588 371 0 um_iw[220]
rlabel metal4 232852 643 232852 643 0 um_iw[221]
rlabel metal4 232116 643 232116 643 0 um_iw[222]
rlabel metal4 231380 371 231380 371 0 um_iw[223]
rlabel metal4 230644 643 230644 643 0 um_iw[224]
rlabel metal4 229908 643 229908 643 0 um_iw[225]
rlabel metal4 229172 371 229172 371 0 um_iw[226]
rlabel metal4 228436 371 228436 371 0 um_iw[227]
rlabel metal4 227700 643 227700 643 0 um_iw[228]
rlabel metal4 226964 371 226964 371 0 um_iw[229]
rlabel via2 28934 8619 28934 8619 0 um_iw[22]
rlabel metal4 226228 779 226228 779 0 um_iw[230]
rlabel metal4 225492 643 225492 643 0 um_iw[231]
rlabel metal4 224756 439 224756 439 0 um_iw[232]
rlabel metal4 224020 643 224020 643 0 um_iw[233]
rlabel via2 236854 9163 236854 9163 0 um_iw[234]
rlabel via2 236026 9435 236026 9435 0 um_iw[235]
rlabel metal2 234922 8041 234922 8041 0 um_iw[236]
rlabel via2 234462 8619 234462 8619 0 um_iw[237]
rlabel via2 233450 9435 233450 9435 0 um_iw[238]
rlabel via2 232622 8619 232622 8619 0 um_iw[239]
rlabel via2 28198 8619 28198 8619 0 um_iw[23]
rlabel via2 231978 9435 231978 9435 0 um_iw[240]
rlabel via2 231702 8619 231702 8619 0 um_iw[241]
rlabel via2 230966 8619 230966 8619 0 um_iw[242]
rlabel via2 229862 9435 229862 9435 0 um_iw[243]
rlabel via2 229218 8619 229218 8619 0 um_iw[244]
rlabel via2 229034 9435 229034 9435 0 um_iw[245]
rlabel via2 228298 9435 228298 9435 0 um_iw[246]
rlabel via2 227010 8619 227010 8619 0 um_iw[247]
rlabel via2 226274 8619 226274 8619 0 um_iw[248]
rlabel via2 225538 8619 225538 8619 0 um_iw[249]
rlabel via2 27462 8619 27462 8619 0 um_iw[24]
rlabel via2 224710 8619 224710 8619 0 um_iw[250]
rlabel metal2 224066 9401 224066 9401 0 um_iw[251]
rlabel metal4 270664 371 270664 371 0 um_iw[252]
rlabel metal4 269928 235 269928 235 0 um_iw[253]
rlabel metal4 269192 371 269192 371 0 um_iw[254]
rlabel metal4 268456 371 268456 371 0 um_iw[255]
rlabel metal4 267720 371 267720 371 0 um_iw[256]
rlabel metal4 266984 371 266984 371 0 um_iw[257]
rlabel metal4 266248 371 266248 371 0 um_iw[258]
rlabel metal4 265512 371 265512 371 0 um_iw[259]
rlabel via2 27370 9707 27370 9707 0 um_iw[25]
rlabel metal4 264776 371 264776 371 0 um_iw[260]
rlabel metal4 264040 371 264040 371 0 um_iw[261]
rlabel metal4 263304 371 263304 371 0 um_iw[262]
rlabel metal4 262568 371 262568 371 0 um_iw[263]
rlabel metal1 262430 2550 262430 2550 0 um_iw[264]
rlabel metal4 261096 371 261096 371 0 um_iw[265]
rlabel metal4 260360 371 260360 371 0 um_iw[266]
rlabel metal4 259624 371 259624 371 0 um_iw[267]
rlabel metal4 258888 371 258888 371 0 um_iw[268]
rlabel metal4 258152 371 258152 371 0 um_iw[269]
rlabel metal1 26220 9690 26220 9690 0 um_iw[26]
rlabel metal1 270388 3978 270388 3978 0 um_iw[270]
rlabel metal1 270526 4794 270526 4794 0 um_iw[271]
rlabel metal2 269514 4811 269514 4811 0 um_iw[272]
rlabel metal1 269744 5814 269744 5814 0 um_iw[273]
rlabel metal1 265420 7514 265420 7514 0 um_iw[274]
rlabel metal1 266248 6630 266248 6630 0 um_iw[275]
rlabel metal2 266202 8891 266202 8891 0 um_iw[276]
rlabel metal2 266294 10047 266294 10047 0 um_iw[277]
rlabel metal1 264960 8058 264960 8058 0 um_iw[278]
rlabel metal2 264362 8891 264362 8891 0 um_iw[279]
rlabel metal2 25254 8177 25254 8177 0 um_iw[27]
rlabel metal2 263350 9163 263350 9163 0 um_iw[280]
rlabel metal2 262522 9163 262522 9163 0 um_iw[281]
rlabel metal1 262108 8602 262108 8602 0 um_iw[282]
rlabel metal2 261786 9231 261786 9231 0 um_iw[283]
rlabel metal2 260498 9435 260498 9435 0 um_iw[284]
rlabel metal2 259946 9435 259946 9435 0 um_iw[285]
rlabel metal2 259210 9979 259210 9979 0 um_iw[286]
rlabel metal2 258290 9435 258290 9435 0 um_iw[287]
rlabel via2 23966 9163 23966 9163 0 um_iw[28]
rlabel metal2 23690 8177 23690 8177 0 um_iw[29]
rlabel metal4 30268 371 30268 371 0 um_iw[2]
rlabel metal2 22954 8177 22954 8177 0 um_iw[30]
rlabel metal2 21758 8959 21758 8959 0 um_iw[31]
rlabel via2 21390 8619 21390 8619 0 um_iw[32]
rlabel metal2 21942 8177 21942 8177 0 um_iw[33]
rlabel metal4 19964 10305 19964 10305 0 um_iw[34]
rlabel metal4 19228 8809 19228 8809 0 um_iw[35]
rlabel metal4 65872 303 65872 303 0 um_iw[36]
rlabel metal4 65136 235 65136 235 0 um_iw[37]
rlabel metal4 64400 235 64400 235 0 um_iw[38]
rlabel metal4 63664 235 63664 235 0 um_iw[39]
rlabel metal4 29532 643 29532 643 0 um_iw[3]
rlabel metal4 62928 303 62928 303 0 um_iw[40]
rlabel metal4 62192 303 62192 303 0 um_iw[41]
rlabel metal4 61456 303 61456 303 0 um_iw[42]
rlabel metal4 60720 303 60720 303 0 um_iw[43]
rlabel metal4 59984 303 59984 303 0 um_iw[44]
rlabel metal4 59248 235 59248 235 0 um_iw[45]
rlabel metal4 58512 303 58512 303 0 um_iw[46]
rlabel metal4 57776 235 57776 235 0 um_iw[47]
rlabel metal4 57040 303 57040 303 0 um_iw[48]
rlabel metal4 56304 303 56304 303 0 um_iw[49]
rlabel metal4 28796 235 28796 235 0 um_iw[4]
rlabel metal4 55568 303 55568 303 0 um_iw[50]
rlabel metal1 55476 2618 55476 2618 0 um_iw[51]
rlabel metal4 54096 371 54096 371 0 um_iw[52]
rlabel metal4 53360 371 53360 371 0 um_iw[53]
rlabel metal1 66102 8330 66102 8330 0 um_iw[54]
rlabel metal2 65550 9299 65550 9299 0 um_iw[55]
rlabel metal2 64722 9435 64722 9435 0 um_iw[56]
rlabel metal2 63986 9435 63986 9435 0 um_iw[57]
rlabel metal2 63434 9979 63434 9979 0 um_iw[58]
rlabel metal2 62514 9979 62514 9979 0 um_iw[59]
rlabel metal4 28060 371 28060 371 0 um_iw[5]
rlabel metal2 61778 9979 61778 9979 0 um_iw[60]
rlabel metal2 61042 9265 61042 9265 0 um_iw[61]
rlabel metal2 60306 9435 60306 9435 0 um_iw[62]
rlabel metal1 59432 8602 59432 8602 0 um_iw[63]
rlabel metal2 58834 9435 58834 9435 0 um_iw[64]
rlabel metal1 58052 9690 58052 9690 0 um_iw[65]
rlabel metal2 57362 9979 57362 9979 0 um_iw[66]
rlabel metal2 56534 9979 56534 9979 0 um_iw[67]
rlabel metal2 55706 9707 55706 9707 0 um_iw[68]
rlabel metal1 55292 9690 55292 9690 0 um_iw[69]
rlabel metal3 27439 2788 27439 2788 0 um_iw[6]
rlabel metal2 53866 9707 53866 9707 0 um_iw[70]
rlabel metal2 53314 9707 53314 9707 0 um_iw[71]
rlabel metal2 99314 901 99314 901 0 um_iw[72]
rlabel metal4 99268 507 99268 507 0 um_iw[73]
rlabel metal4 98532 847 98532 847 0 um_iw[74]
rlabel metal3 97681 3740 97681 3740 0 um_iw[75]
rlabel via3 97037 2788 97037 2788 0 um_iw[76]
rlabel metal4 96324 847 96324 847 0 um_iw[77]
rlabel metal3 95519 2788 95519 2788 0 um_iw[78]
rlabel metal4 94852 371 94852 371 0 um_iw[79]
rlabel metal4 26588 711 26588 711 0 um_iw[7]
rlabel metal3 94047 3060 94047 3060 0 um_iw[80]
rlabel metal4 93380 711 93380 711 0 um_iw[81]
rlabel metal4 92644 371 92644 371 0 um_iw[82]
rlabel metal4 91908 711 91908 711 0 um_iw[83]
rlabel metal4 91172 847 91172 847 0 um_iw[84]
rlabel metal4 90436 711 90436 711 0 um_iw[85]
rlabel metal4 89884 816 89884 816 0 um_iw[86]
rlabel metal4 88964 711 88964 711 0 um_iw[87]
rlabel metal4 88228 779 88228 779 0 um_iw[88]
rlabel metal4 87492 303 87492 303 0 um_iw[89]
rlabel metal4 25852 711 25852 711 0 um_iw[8]
rlabel via2 100510 9707 100510 9707 0 um_iw[90]
rlabel metal4 99268 9693 99268 9693 0 um_iw[91]
rlabel metal4 98532 10237 98532 10237 0 um_iw[92]
rlabel metal1 98164 8602 98164 8602 0 um_iw[93]
rlabel via2 97566 8619 97566 8619 0 um_iw[94]
rlabel metal1 96646 9690 96646 9690 0 um_iw[95]
rlabel via2 96094 9707 96094 9707 0 um_iw[96]
rlabel via2 95082 8619 95082 8619 0 um_iw[97]
rlabel via2 94622 8619 94622 8619 0 um_iw[98]
rlabel via2 93518 9707 93518 9707 0 um_iw[99]
rlabel metal1 24840 2618 24840 2618 0 um_iw[9]
rlabel metal4 18492 235 18492 235 0 um_ow[0]
rlabel metal4 83812 711 83812 711 0 um_ow[100]
rlabel metal4 83076 507 83076 507 0 um_ow[101]
rlabel metal4 82340 575 82340 575 0 um_ow[102]
rlabel metal4 81604 711 81604 711 0 um_ow[103]
rlabel metal4 80868 575 80868 575 0 um_ow[104]
rlabel metal2 79994 1105 79994 1105 0 um_ow[105]
rlabel metal4 79396 575 79396 575 0 um_ow[106]
rlabel metal4 78660 711 78660 711 0 um_ow[107]
rlabel metal4 77924 507 77924 507 0 um_ow[108]
rlabel metal4 77188 575 77188 575 0 um_ow[109]
rlabel metal4 11132 439 11132 439 0 um_ow[10]
rlabel metal4 76452 711 76452 711 0 um_ow[110]
rlabel metal4 75716 575 75716 575 0 um_ow[111]
rlabel metal4 74980 507 74980 507 0 um_ow[112]
rlabel metal4 74244 507 74244 507 0 um_ow[113]
rlabel metal4 73508 575 73508 575 0 um_ow[114]
rlabel metal4 72772 507 72772 507 0 um_ow[115]
rlabel metal4 72036 575 72036 575 0 um_ow[116]
rlabel metal4 71300 575 71300 575 0 um_ow[117]
rlabel metal4 70564 507 70564 507 0 um_ow[118]
rlabel metal4 69828 507 69828 507 0 um_ow[119]
rlabel metal4 10396 439 10396 439 0 um_ow[11]
rlabel metal4 86756 10645 86756 10645 0 um_ow[120]
rlabel metal4 86020 10305 86020 10305 0 um_ow[121]
rlabel metal4 85284 10441 85284 10441 0 um_ow[122]
rlabel metal4 84548 10441 84548 10441 0 um_ow[123]
rlabel metal4 83812 10441 83812 10441 0 um_ow[124]
rlabel metal4 83076 10441 83076 10441 0 um_ow[125]
rlabel metal4 82340 10645 82340 10645 0 um_ow[126]
rlabel metal4 81604 10645 81604 10645 0 um_ow[127]
rlabel metal4 80868 10305 80868 10305 0 um_ow[128]
rlabel metal1 79948 9554 79948 9554 0 um_ow[129]
rlabel metal4 9660 575 9660 575 0 um_ow[12]
rlabel metal4 79396 10441 79396 10441 0 um_ow[130]
rlabel metal4 78660 10305 78660 10305 0 um_ow[131]
rlabel via2 77326 9571 77326 9571 0 um_ow[132]
rlabel metal4 77188 10305 77188 10305 0 um_ow[133]
rlabel metal4 76452 10169 76452 10169 0 um_ow[134]
rlabel via2 74750 9571 74750 9571 0 um_ow[135]
rlabel metal2 74750 8993 74750 8993 0 um_ow[136]
rlabel metal4 74244 10169 74244 10169 0 um_ow[137]
rlabel via2 73462 9027 73462 9027 0 um_ow[138]
rlabel via2 72174 9571 72174 9571 0 um_ow[139]
rlabel metal4 8924 235 8924 235 0 um_ow[13]
rlabel metal4 72036 10577 72036 10577 0 um_ow[140]
rlabel metal4 71300 10441 71300 10441 0 um_ow[141]
rlabel metal1 69966 9554 69966 9554 0 um_ow[142]
rlabel metal4 69828 10305 69828 10305 0 um_ow[143]
rlabel metal4 120888 303 120888 303 0 um_ow[144]
rlabel metal4 120152 303 120152 303 0 um_ow[145]
rlabel metal4 119416 303 119416 303 0 um_ow[146]
rlabel metal2 118726 901 118726 901 0 um_ow[147]
rlabel metal4 117944 303 117944 303 0 um_ow[148]
rlabel metal4 117208 235 117208 235 0 um_ow[149]
rlabel metal4 8188 303 8188 303 0 um_ow[14]
rlabel metal1 117760 2550 117760 2550 0 um_ow[150]
rlabel metal4 115736 235 115736 235 0 um_ow[151]
rlabel metal4 115000 235 115000 235 0 um_ow[152]
rlabel metal4 114264 235 114264 235 0 um_ow[153]
rlabel metal2 120750 1700 120750 1700 0 um_ow[154]
rlabel metal4 112792 235 112792 235 0 um_ow[155]
rlabel metal4 112056 235 112056 235 0 um_ow[156]
rlabel metal4 111320 235 111320 235 0 um_ow[157]
rlabel metal4 110584 235 110584 235 0 um_ow[158]
rlabel metal4 109848 235 109848 235 0 um_ow[159]
rlabel metal4 7452 575 7452 575 0 um_ow[15]
rlabel metal4 109112 235 109112 235 0 um_ow[160]
rlabel metal4 108376 235 108376 235 0 um_ow[161]
rlabel metal4 107640 235 107640 235 0 um_ow[162]
rlabel metal4 106904 235 106904 235 0 um_ow[163]
rlabel metal4 106168 235 106168 235 0 um_ow[164]
rlabel metal4 105432 235 105432 235 0 um_ow[165]
rlabel metal4 104696 235 104696 235 0 um_ow[166]
rlabel metal4 103960 235 103960 235 0 um_ow[167]
rlabel metal4 120888 10509 120888 10509 0 um_ow[168]
rlabel metal4 120152 10509 120152 10509 0 um_ow[169]
rlabel metal4 6716 711 6716 711 0 um_ow[16]
rlabel metal4 119416 10509 119416 10509 0 um_ow[170]
rlabel metal4 118680 10509 118680 10509 0 um_ow[171]
rlabel metal4 117944 10509 117944 10509 0 um_ow[172]
rlabel metal4 117208 10509 117208 10509 0 um_ow[173]
rlabel metal4 116472 10509 116472 10509 0 um_ow[174]
rlabel metal4 115736 10509 115736 10509 0 um_ow[175]
rlabel metal4 115000 10509 115000 10509 0 um_ow[176]
rlabel metal4 114264 10509 114264 10509 0 um_ow[177]
rlabel metal4 113528 10509 113528 10509 0 um_ow[178]
rlabel metal4 112792 10509 112792 10509 0 um_ow[179]
rlabel metal4 5980 439 5980 439 0 um_ow[17]
rlabel metal4 112056 10509 112056 10509 0 um_ow[180]
rlabel metal4 111320 10509 111320 10509 0 um_ow[181]
rlabel metal4 110584 10509 110584 10509 0 um_ow[182]
rlabel metal4 109848 10509 109848 10509 0 um_ow[183]
rlabel metal4 109112 10509 109112 10509 0 um_ow[184]
rlabel metal4 108376 10509 108376 10509 0 um_ow[185]
rlabel metal4 107640 10509 107640 10509 0 um_ow[186]
rlabel metal4 106904 10509 106904 10509 0 um_ow[187]
rlabel metal4 106168 10509 106168 10509 0 um_ow[188]
rlabel metal4 105432 10509 105432 10509 0 um_ow[189]
rlabel metal4 5244 575 5244 575 0 um_ow[18]
rlabel metal4 104696 10509 104696 10509 0 um_ow[190]
rlabel metal4 103960 10509 103960 10509 0 um_ow[191]
rlabel via3 155043 2924 155043 2924 0 um_ow[192]
rlabel via3 154307 3332 154307 3332 0 um_ow[193]
rlabel metal3 153617 2924 153617 2924 0 um_ow[194]
rlabel metal4 152812 711 152812 711 0 um_ow[195]
rlabel metal4 152076 779 152076 779 0 um_ow[196]
rlabel metal4 151340 371 151340 371 0 um_ow[197]
rlabel metal4 150604 779 150604 779 0 um_ow[198]
rlabel metal4 149868 439 149868 439 0 um_ow[199]
rlabel metal4 4508 711 4508 711 0 um_ow[19]
rlabel metal4 17756 575 17756 575 0 um_ow[1]
rlabel metal1 151386 2346 151386 2346 0 um_ow[200]
rlabel metal4 148396 439 148396 439 0 um_ow[201]
rlabel metal2 147890 663 147890 663 0 um_ow[202]
rlabel metal1 147890 510 147890 510 0 um_ow[203]
rlabel metal2 147706 867 147706 867 0 um_ow[204]
rlabel metal1 150742 1394 150742 1394 0 um_ow[205]
rlabel via3 144739 3196 144739 3196 0 um_ow[206]
rlabel metal2 151018 1054 151018 1054 0 um_ow[207]
rlabel metal4 143244 371 143244 371 0 um_ow[208]
rlabel metal4 142508 439 142508 439 0 um_ow[209]
rlabel metal4 3772 575 3772 575 0 um_ow[20]
rlabel metal4 141772 439 141772 439 0 um_ow[210]
rlabel metal4 141036 779 141036 779 0 um_ow[211]
rlabel metal4 140300 983 140300 983 0 um_ow[212]
rlabel metal4 139564 575 139564 575 0 um_ow[213]
rlabel metal4 138828 439 138828 439 0 um_ow[214]
rlabel metal4 138092 371 138092 371 0 um_ow[215]
rlabel metal4 155020 10305 155020 10305 0 um_ow[216]
rlabel metal4 154284 10577 154284 10577 0 um_ow[217]
rlabel metal4 153548 10441 153548 10441 0 um_ow[218]
rlabel metal4 152812 10441 152812 10441 0 um_ow[219]
rlabel metal4 3036 439 3036 439 0 um_ow[21]
rlabel metal4 152076 10441 152076 10441 0 um_ow[220]
rlabel metal4 151340 10441 151340 10441 0 um_ow[221]
rlabel metal4 150604 10441 150604 10441 0 um_ow[222]
rlabel metal4 149868 10305 149868 10305 0 um_ow[223]
rlabel metal4 149132 10441 149132 10441 0 um_ow[224]
rlabel metal4 148396 10509 148396 10509 0 um_ow[225]
rlabel metal2 148442 10047 148442 10047 0 um_ow[226]
rlabel metal4 146924 10441 146924 10441 0 um_ow[227]
rlabel metal4 146188 10441 146188 10441 0 um_ow[228]
rlabel metal4 145452 10441 145452 10441 0 um_ow[229]
rlabel metal4 2300 371 2300 371 0 um_ow[22]
rlabel metal4 144716 10305 144716 10305 0 um_ow[230]
rlabel metal4 143980 10441 143980 10441 0 um_ow[231]
rlabel metal4 143244 10441 143244 10441 0 um_ow[232]
rlabel metal4 142508 10509 142508 10509 0 um_ow[233]
rlabel metal4 141772 10441 141772 10441 0 um_ow[234]
rlabel metal4 141036 10441 141036 10441 0 um_ow[235]
rlabel metal4 140300 10441 140300 10441 0 um_ow[236]
rlabel metal4 139564 10305 139564 10305 0 um_ow[237]
rlabel metal4 138828 10441 138828 10441 0 um_ow[238]
rlabel metal4 138092 10509 138092 10509 0 um_ow[239]
rlabel metal4 1564 575 1564 575 0 um_ow[23]
rlabel metal4 189152 303 189152 303 0 um_ow[240]
rlabel metal4 188416 303 188416 303 0 um_ow[241]
rlabel metal4 187680 303 187680 303 0 um_ow[242]
rlabel metal4 186944 303 186944 303 0 um_ow[243]
rlabel metal4 186208 235 186208 235 0 um_ow[244]
rlabel metal4 185472 303 185472 303 0 um_ow[245]
rlabel metal4 184736 303 184736 303 0 um_ow[246]
rlabel metal4 184000 303 184000 303 0 um_ow[247]
rlabel metal4 183264 303 183264 303 0 um_ow[248]
rlabel metal4 182528 303 182528 303 0 um_ow[249]
rlabel metal4 18492 10441 18492 10441 0 um_ow[24]
rlabel metal4 181792 303 181792 303 0 um_ow[250]
rlabel metal4 181056 235 181056 235 0 um_ow[251]
rlabel metal4 180320 371 180320 371 0 um_ow[252]
rlabel metal4 179584 371 179584 371 0 um_ow[253]
rlabel metal4 178848 371 178848 371 0 um_ow[254]
rlabel metal4 178112 371 178112 371 0 um_ow[255]
rlabel metal4 177376 371 177376 371 0 um_ow[256]
rlabel metal4 176640 371 176640 371 0 um_ow[257]
rlabel metal4 175904 303 175904 303 0 um_ow[258]
rlabel metal4 175168 371 175168 371 0 um_ow[259]
rlabel metal4 17756 10441 17756 10441 0 um_ow[25]
rlabel metal4 174432 371 174432 371 0 um_ow[260]
rlabel metal4 173696 371 173696 371 0 um_ow[261]
rlabel metal4 172960 371 172960 371 0 um_ow[262]
rlabel metal4 172224 371 172224 371 0 um_ow[263]
rlabel metal4 189152 10509 189152 10509 0 um_ow[264]
rlabel metal4 188416 10509 188416 10509 0 um_ow[265]
rlabel metal4 187680 10509 187680 10509 0 um_ow[266]
rlabel metal4 186944 10509 186944 10509 0 um_ow[267]
rlabel metal4 186208 10509 186208 10509 0 um_ow[268]
rlabel metal4 185472 10509 185472 10509 0 um_ow[269]
rlabel metal4 17020 10441 17020 10441 0 um_ow[26]
rlabel metal4 184736 10509 184736 10509 0 um_ow[270]
rlabel metal4 184000 10509 184000 10509 0 um_ow[271]
rlabel metal4 183264 10509 183264 10509 0 um_ow[272]
rlabel metal4 182528 10509 182528 10509 0 um_ow[273]
rlabel metal4 181792 10509 181792 10509 0 um_ow[274]
rlabel metal4 181056 10577 181056 10577 0 um_ow[275]
rlabel metal4 180320 10509 180320 10509 0 um_ow[276]
rlabel metal4 179584 10645 179584 10645 0 um_ow[277]
rlabel metal4 178848 10509 178848 10509 0 um_ow[278]
rlabel metal1 177882 9554 177882 9554 0 um_ow[279]
rlabel metal4 16284 10441 16284 10441 0 um_ow[27]
rlabel metal4 177376 10509 177376 10509 0 um_ow[280]
rlabel metal2 176778 9605 176778 9605 0 um_ow[281]
rlabel metal4 175904 10509 175904 10509 0 um_ow[282]
rlabel metal4 175168 10509 175168 10509 0 um_ow[283]
rlabel metal4 174432 10509 174432 10509 0 um_ow[284]
rlabel metal4 173696 10509 173696 10509 0 um_ow[285]
rlabel metal4 172960 10577 172960 10577 0 um_ow[286]
rlabel metal4 172224 10645 172224 10645 0 um_ow[287]
rlabel metal3 223399 3740 223399 3740 0 um_ow[288]
rlabel metal1 227194 2448 227194 2448 0 um_ow[289]
rlabel metal4 15548 10441 15548 10441 0 um_ow[28]
rlabel metal4 221812 371 221812 371 0 um_ow[290]
rlabel metal2 225906 3196 225906 3196 0 um_ow[291]
rlabel metal2 226458 1054 226458 1054 0 um_ow[292]
rlabel metal1 224986 2380 224986 2380 0 um_ow[293]
rlabel via3 218891 3740 218891 3740 0 um_ow[294]
rlabel metal4 218132 779 218132 779 0 um_ow[295]
rlabel metal3 217557 3196 217557 3196 0 um_ow[296]
rlabel metal3 216913 2924 216913 2924 0 um_ow[297]
rlabel metal4 215924 439 215924 439 0 um_ow[298]
rlabel via3 215211 4012 215211 4012 0 um_ow[299]
rlabel metal4 14812 10441 14812 10441 0 um_ow[29]
rlabel metal4 17020 439 17020 439 0 um_ow[2]
rlabel metal4 214452 235 214452 235 0 um_ow[300]
rlabel metal4 213716 303 213716 303 0 um_ow[301]
rlabel metal4 212980 235 212980 235 0 um_ow[302]
rlabel metal4 212244 983 212244 983 0 um_ow[303]
rlabel via3 211531 3060 211531 3060 0 um_ow[304]
rlabel metal1 209024 2482 209024 2482 0 um_ow[305]
rlabel metal4 210036 779 210036 779 0 um_ow[306]
rlabel metal4 209300 303 209300 303 0 um_ow[307]
rlabel metal4 208564 507 208564 507 0 um_ow[308]
rlabel metal4 207828 235 207828 235 0 um_ow[309]
rlabel metal4 14076 10441 14076 10441 0 um_ow[30]
rlabel metal4 207092 507 207092 507 0 um_ow[310]
rlabel metal4 206356 507 206356 507 0 um_ow[311]
rlabel metal4 223284 10441 223284 10441 0 um_ow[312]
rlabel metal4 222548 10441 222548 10441 0 um_ow[313]
rlabel metal4 221812 10305 221812 10305 0 um_ow[314]
rlabel metal4 221076 10577 221076 10577 0 um_ow[315]
rlabel metal4 220340 10509 220340 10509 0 um_ow[316]
rlabel metal4 219604 10441 219604 10441 0 um_ow[317]
rlabel metal4 218868 10441 218868 10441 0 um_ow[318]
rlabel metal4 218132 10645 218132 10645 0 um_ow[319]
rlabel metal4 13340 10305 13340 10305 0 um_ow[31]
rlabel metal4 217396 10441 217396 10441 0 um_ow[320]
rlabel metal4 216660 10305 216660 10305 0 um_ow[321]
rlabel metal4 215924 10441 215924 10441 0 um_ow[322]
rlabel metal4 215188 10169 215188 10169 0 um_ow[323]
rlabel metal4 214452 10441 214452 10441 0 um_ow[324]
rlabel metal4 213716 10441 213716 10441 0 um_ow[325]
rlabel metal4 212980 10645 212980 10645 0 um_ow[326]
rlabel metal4 212244 10441 212244 10441 0 um_ow[327]
rlabel metal4 211508 10305 211508 10305 0 um_ow[328]
rlabel metal4 210772 10441 210772 10441 0 um_ow[329]
rlabel metal4 12604 10441 12604 10441 0 um_ow[32]
rlabel metal4 210036 10577 210036 10577 0 um_ow[330]
rlabel metal4 209300 10441 209300 10441 0 um_ow[331]
rlabel metal4 208564 10441 208564 10441 0 um_ow[332]
rlabel metal4 207828 10645 207828 10645 0 um_ow[333]
rlabel metal4 207092 10441 207092 10441 0 um_ow[334]
rlabel metal4 206356 10441 206356 10441 0 um_ow[335]
rlabel metal4 257416 235 257416 235 0 um_ow[336]
rlabel metal4 256680 235 256680 235 0 um_ow[337]
rlabel metal4 255944 371 255944 371 0 um_ow[338]
rlabel metal4 255208 371 255208 371 0 um_ow[339]
rlabel metal4 11868 10441 11868 10441 0 um_ow[33]
rlabel metal4 254472 371 254472 371 0 um_ow[340]
rlabel metal4 253736 235 253736 235 0 um_ow[341]
rlabel metal4 253000 303 253000 303 0 um_ow[342]
rlabel metal4 252264 235 252264 235 0 um_ow[343]
rlabel metal4 251528 235 251528 235 0 um_ow[344]
rlabel metal4 250792 371 250792 371 0 um_ow[345]
rlabel metal4 250056 371 250056 371 0 um_ow[346]
rlabel metal4 249320 235 249320 235 0 um_ow[347]
rlabel metal4 248584 235 248584 235 0 um_ow[348]
rlabel metal4 247848 371 247848 371 0 um_ow[349]
rlabel metal4 11132 10441 11132 10441 0 um_ow[34]
rlabel metal4 247112 371 247112 371 0 um_ow[350]
rlabel metal4 246376 371 246376 371 0 um_ow[351]
rlabel metal4 245640 235 245640 235 0 um_ow[352]
rlabel metal4 244904 371 244904 371 0 um_ow[353]
rlabel metal4 244168 371 244168 371 0 um_ow[354]
rlabel metal4 243432 371 243432 371 0 um_ow[355]
rlabel metal4 242696 235 242696 235 0 um_ow[356]
rlabel metal4 241960 371 241960 371 0 um_ow[357]
rlabel metal4 241224 371 241224 371 0 um_ow[358]
rlabel metal4 240488 371 240488 371 0 um_ow[359]
rlabel metal4 10396 10441 10396 10441 0 um_ow[35]
rlabel metal4 257416 10509 257416 10509 0 um_ow[360]
rlabel metal4 256680 10509 256680 10509 0 um_ow[361]
rlabel metal4 255944 10509 255944 10509 0 um_ow[362]
rlabel metal4 255208 10509 255208 10509 0 um_ow[363]
rlabel metal4 254472 10509 254472 10509 0 um_ow[364]
rlabel metal4 253736 10509 253736 10509 0 um_ow[365]
rlabel metal4 253000 10577 253000 10577 0 um_ow[366]
rlabel metal4 252264 10509 252264 10509 0 um_ow[367]
rlabel metal4 251528 10509 251528 10509 0 um_ow[368]
rlabel metal4 250792 10509 250792 10509 0 um_ow[369]
rlabel metal4 9660 10441 9660 10441 0 um_ow[36]
rlabel metal4 250056 10509 250056 10509 0 um_ow[370]
rlabel metal4 249320 10509 249320 10509 0 um_ow[371]
rlabel metal4 248584 10509 248584 10509 0 um_ow[372]
rlabel metal4 247848 10509 247848 10509 0 um_ow[373]
rlabel metal4 247112 10509 247112 10509 0 um_ow[374]
rlabel metal4 246376 10509 246376 10509 0 um_ow[375]
rlabel metal4 245640 10577 245640 10577 0 um_ow[376]
rlabel metal4 244904 10509 244904 10509 0 um_ow[377]
rlabel metal1 245134 9520 245134 9520 0 um_ow[378]
rlabel metal4 243432 10509 243432 10509 0 um_ow[379]
rlabel metal4 8924 10441 8924 10441 0 um_ow[37]
rlabel metal4 242696 10509 242696 10509 0 um_ow[380]
rlabel metal4 241960 10509 241960 10509 0 um_ow[381]
rlabel metal4 241224 10509 241224 10509 0 um_ow[382]
rlabel metal4 240488 10509 240488 10509 0 um_ow[383]
rlabel metal4 8188 10305 8188 10305 0 um_ow[38]
rlabel metal4 7452 10441 7452 10441 0 um_ow[39]
rlabel metal4 16284 439 16284 439 0 um_ow[3]
rlabel metal4 6716 10441 6716 10441 0 um_ow[40]
rlabel metal4 5980 10441 5980 10441 0 um_ow[41]
rlabel metal4 5244 10441 5244 10441 0 um_ow[42]
rlabel metal4 4508 10441 4508 10441 0 um_ow[43]
rlabel metal4 3772 10441 3772 10441 0 um_ow[44]
rlabel metal4 3036 10305 3036 10305 0 um_ow[45]
rlabel metal4 2300 10441 2300 10441 0 um_ow[46]
rlabel metal4 1564 10441 1564 10441 0 um_ow[47]
rlabel metal4 52624 235 52624 235 0 um_ow[48]
rlabel metal4 51888 371 51888 371 0 um_ow[49]
rlabel metal4 15548 575 15548 575 0 um_ow[4]
rlabel metal4 51152 371 51152 371 0 um_ow[50]
rlabel metal4 50416 371 50416 371 0 um_ow[51]
rlabel metal4 49680 371 49680 371 0 um_ow[52]
rlabel metal4 48944 371 48944 371 0 um_ow[53]
rlabel metal4 48208 371 48208 371 0 um_ow[54]
rlabel metal4 47472 371 47472 371 0 um_ow[55]
rlabel metal4 46736 371 46736 371 0 um_ow[56]
rlabel metal4 46000 371 46000 371 0 um_ow[57]
rlabel metal4 45264 371 45264 371 0 um_ow[58]
rlabel metal4 44528 371 44528 371 0 um_ow[59]
rlabel metal4 14812 711 14812 711 0 um_ow[5]
rlabel metal4 43792 371 43792 371 0 um_ow[60]
rlabel metal4 43056 371 43056 371 0 um_ow[61]
rlabel metal4 42320 371 42320 371 0 um_ow[62]
rlabel metal4 41584 371 41584 371 0 um_ow[63]
rlabel metal4 40848 371 40848 371 0 um_ow[64]
rlabel metal4 40112 371 40112 371 0 um_ow[65]
rlabel metal4 39376 235 39376 235 0 um_ow[66]
rlabel metal4 38640 371 38640 371 0 um_ow[67]
rlabel metal4 37904 371 37904 371 0 um_ow[68]
rlabel metal4 37168 371 37168 371 0 um_ow[69]
rlabel metal4 14076 575 14076 575 0 um_ow[6]
rlabel metal4 36432 371 36432 371 0 um_ow[70]
rlabel metal4 35696 371 35696 371 0 um_ow[71]
rlabel metal4 52624 10645 52624 10645 0 um_ow[72]
rlabel metal4 51888 10509 51888 10509 0 um_ow[73]
rlabel metal4 51152 10509 51152 10509 0 um_ow[74]
rlabel metal4 50416 10509 50416 10509 0 um_ow[75]
rlabel metal4 49680 10509 49680 10509 0 um_ow[76]
rlabel metal4 48944 10509 48944 10509 0 um_ow[77]
rlabel metal4 48208 10509 48208 10509 0 um_ow[78]
rlabel metal4 47472 10509 47472 10509 0 um_ow[79]
rlabel metal4 13340 371 13340 371 0 um_ow[7]
rlabel metal4 46736 10509 46736 10509 0 um_ow[80]
rlabel metal4 46000 10509 46000 10509 0 um_ow[81]
rlabel metal4 45264 10509 45264 10509 0 um_ow[82]
rlabel metal4 44528 10509 44528 10509 0 um_ow[83]
rlabel metal4 43792 10509 43792 10509 0 um_ow[84]
rlabel metal4 43056 10509 43056 10509 0 um_ow[85]
rlabel metal4 42320 10509 42320 10509 0 um_ow[86]
rlabel metal4 41584 10509 41584 10509 0 um_ow[87]
rlabel metal4 40848 10509 40848 10509 0 um_ow[88]
rlabel metal4 40112 10509 40112 10509 0 um_ow[89]
rlabel metal4 12604 575 12604 575 0 um_ow[8]
rlabel metal4 39376 10509 39376 10509 0 um_ow[90]
rlabel metal4 38640 10509 38640 10509 0 um_ow[91]
rlabel metal4 37904 10509 37904 10509 0 um_ow[92]
rlabel metal4 37168 10509 37168 10509 0 um_ow[93]
rlabel metal4 36432 10509 36432 10509 0 um_ow[94]
rlabel metal4 35696 10509 35696 10509 0 um_ow[95]
rlabel metal4 86756 507 86756 507 0 um_ow[96]
rlabel metal4 86020 575 86020 575 0 um_ow[97]
rlabel metal4 85284 235 85284 235 0 um_ow[98]
rlabel metal4 84548 575 84548 575 0 um_ow[99]
rlabel metal4 11868 575 11868 575 0 um_ow[9]
rlabel metal1 252816 4794 252816 4794 0 zbuf_bus_ena_I.e
rlabel metal2 253138 6562 253138 6562 0 zbuf_bus_ena_I.genblk1.l
rlabel metal1 185610 6154 185610 6154 0 zbuf_bus_ena_I.z
rlabel metal2 268042 7242 268042 7242 0 zbuf_bus_iw_I\[0\].genblk1.l
rlabel metal2 263166 6086 263166 6086 0 zbuf_bus_iw_I\[10\].genblk1.l
rlabel metal2 262522 5814 262522 5814 0 zbuf_bus_iw_I\[11\].genblk1.l
rlabel metal2 261694 5882 261694 5882 0 zbuf_bus_iw_I\[12\].genblk1.l
rlabel metal2 260406 5882 260406 5882 0 zbuf_bus_iw_I\[13\].genblk1.l
rlabel via2 266938 5253 266938 5253 0 zbuf_bus_iw_I\[14\].genblk1.l
rlabel metal1 266892 4250 266892 4250 0 zbuf_bus_iw_I\[15\].genblk1.l
rlabel metal1 267950 3910 267950 3910 0 zbuf_bus_iw_I\[16\].genblk1.l
rlabel metal1 268594 4624 268594 4624 0 zbuf_bus_iw_I\[17\].genblk1.l
rlabel metal1 269560 5338 269560 5338 0 zbuf_bus_iw_I\[1\].genblk1.l
rlabel metal1 268410 5712 268410 5712 0 zbuf_bus_iw_I\[2\].genblk1.l
rlabel metal2 267858 6732 267858 6732 0 zbuf_bus_iw_I\[3\].genblk1.l
rlabel metal2 266938 6426 266938 6426 0 zbuf_bus_iw_I\[4\].genblk1.l
rlabel metal2 266662 6460 266662 6460 0 zbuf_bus_iw_I\[5\].genblk1.l
rlabel metal1 266708 5338 266708 5338 0 zbuf_bus_iw_I\[6\].genblk1.l
rlabel metal2 267766 6018 267766 6018 0 zbuf_bus_iw_I\[7\].genblk1.l
rlabel metal1 268502 5338 268502 5338 0 zbuf_bus_iw_I\[8\].genblk1.l
rlabel metal2 265282 6086 265282 6086 0 zbuf_bus_iw_I\[9\].genblk1.l
rlabel metal2 248446 6970 248446 6970 0 zbuf_bus_sel_I\[0\].genblk1.l
rlabel metal2 227010 7004 227010 7004 0 zbuf_bus_sel_I\[0\].z
rlabel metal1 225446 7480 225446 7480 0 zbuf_bus_sel_I\[1\].genblk1.l
rlabel metal1 225446 7378 225446 7378 0 zbuf_bus_sel_I\[1\].z
rlabel via2 213486 7395 213486 7395 0 zbuf_bus_sel_I\[2\].genblk1.l
rlabel viali 117622 6289 117622 6289 0 zbuf_bus_sel_I\[2\].z
rlabel metal2 213210 7021 213210 7021 0 zbuf_bus_sel_I\[3\].genblk1.l
rlabel metal2 168866 6154 168866 6154 0 zbuf_bus_sel_I\[3\].z
rlabel via2 213118 6307 213118 6307 0 zbuf_bus_sel_I\[4\].genblk1.l
rlabel metal2 116518 5831 116518 5831 0 zbuf_bus_sel_I\[4\].z
<< properties >>
string FIXED_BBOX 0 0 272600 11000
<< end >>
