VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_urish_dffram
  CLASS BLOCK ;
  FOREIGN tt_um_urish_dffram ;
  ORIGIN 0.000 0.000 ;
  SIZE 679.880 BY 220.320 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 206.850 158.850 220.320 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 162.230 219.320 162.530 220.320 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 217.420 155.170 220.320 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 218.780 151.490 220.320 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 215.380 147.810 220.320 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 216.740 144.130 220.320 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 217.420 140.450 220.320 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 215.380 136.770 220.320 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 218.780 133.090 220.320 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 215.380 129.410 220.320 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 214.020 125.730 220.320 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 215.380 122.050 220.320 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 216.740 118.370 220.320 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 216.740 114.690 220.320 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 216.740 111.010 220.320 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 218.100 107.330 220.320 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 218.780 103.650 220.320 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 216.740 99.970 220.320 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 215.380 96.290 220.320 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 218.780 33.730 220.320 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 214.700 30.050 220.320 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 214.700 26.370 220.320 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 216.060 22.690 220.320 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 211.300 19.010 220.320 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 214.700 15.330 220.320 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 214.700 11.650 220.320 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 214.700 7.970 220.320 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 214.700 63.170 220.320 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 214.700 59.490 220.320 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 214.700 55.810 220.320 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 214.700 52.130 220.320 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 214.700 48.450 220.320 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 211.300 44.770 220.320 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 218.780 41.090 220.320 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 214.700 37.410 220.320 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 199.740 92.610 220.320 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 199.060 88.930 220.320 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 199.740 85.250 220.320 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 199.740 81.570 220.320 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 199.740 77.890 220.320 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 199.060 74.210 220.320 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 199.740 70.530 220.320 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 199.740 66.850 220.320 ;
    END
  END uo_out[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 5.200 22.640 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 5.200 176.240 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 5.200 329.840 29.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 136.540 329.840 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 5.200 483.440 29.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 136.540 483.440 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 5.200 637.040 56.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 134.085 637.040 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.460 13.360 659.060 152.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 5.200 99.440 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 5.200 253.040 29.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 136.540 253.040 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 5.200 406.640 29.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 136.540 406.640 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 5.200 560.240 29.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 136.540 560.240 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 660.220 13.360 661.820 152.560 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 213.465 674.550 215.070 ;
        RECT 5.330 208.025 674.550 210.855 ;
        RECT 5.330 202.585 674.550 205.415 ;
        RECT 5.330 197.145 674.550 199.975 ;
        RECT 5.330 191.705 674.550 194.535 ;
        RECT 5.330 186.265 674.550 189.095 ;
        RECT 5.330 180.825 674.550 183.655 ;
        RECT 5.330 175.385 674.550 178.215 ;
        RECT 5.330 169.945 674.550 172.775 ;
        RECT 5.330 164.505 674.550 167.335 ;
        RECT 5.330 159.065 674.550 161.895 ;
        RECT 5.330 153.625 674.550 156.455 ;
        RECT 5.330 149.410 674.550 151.015 ;
        RECT 5.330 148.185 223.290 149.410 ;
        RECT 5.330 142.745 223.290 145.575 ;
        RECT 5.330 137.305 223.290 140.135 ;
        RECT 5.330 131.865 223.290 134.695 ;
        RECT 5.330 126.425 223.290 129.255 ;
        RECT 5.330 120.985 223.290 123.815 ;
        RECT 5.330 115.545 223.290 118.375 ;
        RECT 5.330 110.105 223.290 112.935 ;
        RECT 5.330 104.665 223.290 107.495 ;
        RECT 5.330 99.225 223.290 102.055 ;
        RECT 5.330 93.785 223.290 96.615 ;
        RECT 5.330 88.345 223.290 91.175 ;
        RECT 5.330 82.905 223.290 85.735 ;
        RECT 5.330 77.465 223.290 80.295 ;
        RECT 5.330 72.025 223.290 74.855 ;
        RECT 5.330 66.585 223.290 69.415 ;
        RECT 5.330 61.145 223.290 63.975 ;
        RECT 5.330 55.705 223.290 58.535 ;
        RECT 5.330 50.265 223.290 53.095 ;
        RECT 5.330 44.825 223.290 47.655 ;
        RECT 5.330 39.385 223.290 42.215 ;
        RECT 5.330 33.945 223.290 36.775 ;
        RECT 5.330 28.505 223.290 31.335 ;
        RECT 5.330 23.065 223.290 25.895 ;
        RECT 5.330 17.625 223.290 20.455 ;
        RECT 5.330 12.185 674.550 15.015 ;
        RECT 5.330 6.745 674.550 9.575 ;
      LAYER li1 ;
        RECT 5.520 5.355 674.360 214.965 ;
      LAYER met1 ;
        RECT 5.520 5.200 674.360 215.120 ;
      LAYER met2 ;
        RECT 8.830 5.255 661.790 218.805 ;
      LAYER met3 ;
        RECT 7.630 5.275 661.810 218.785 ;
      LAYER met4 ;
        RECT 8.370 214.300 10.950 218.785 ;
        RECT 12.050 214.300 14.630 218.785 ;
        RECT 15.730 214.300 18.310 218.785 ;
        RECT 7.655 210.900 18.310 214.300 ;
        RECT 19.410 215.660 21.990 218.785 ;
        RECT 23.090 215.660 25.670 218.785 ;
        RECT 19.410 215.520 25.670 215.660 ;
        RECT 19.410 210.900 20.640 215.520 ;
        RECT 7.655 29.680 20.640 210.900 ;
        RECT 23.040 214.300 25.670 215.520 ;
        RECT 26.770 214.300 29.350 218.785 ;
        RECT 30.450 218.380 33.030 218.785 ;
        RECT 34.130 218.380 36.710 218.785 ;
        RECT 30.450 214.300 36.710 218.380 ;
        RECT 37.810 218.380 40.390 218.785 ;
        RECT 41.490 218.380 44.070 218.785 ;
        RECT 37.810 214.300 44.070 218.380 ;
        RECT 23.040 210.900 44.070 214.300 ;
        RECT 45.170 214.300 47.750 218.785 ;
        RECT 48.850 214.300 51.430 218.785 ;
        RECT 52.530 214.300 55.110 218.785 ;
        RECT 56.210 214.300 58.790 218.785 ;
        RECT 59.890 214.300 62.470 218.785 ;
        RECT 63.570 214.300 66.150 218.785 ;
        RECT 45.170 210.900 66.150 214.300 ;
        RECT 23.040 199.340 66.150 210.900 ;
        RECT 67.250 199.340 69.830 218.785 ;
        RECT 70.930 199.340 73.510 218.785 ;
        RECT 23.040 198.660 73.510 199.340 ;
        RECT 74.610 199.340 77.190 218.785 ;
        RECT 78.290 199.340 80.870 218.785 ;
        RECT 81.970 199.340 84.550 218.785 ;
        RECT 85.650 199.340 88.230 218.785 ;
        RECT 74.610 198.660 88.230 199.340 ;
        RECT 89.330 199.340 91.910 218.785 ;
        RECT 93.010 214.980 95.590 218.785 ;
        RECT 96.690 216.340 99.270 218.785 ;
        RECT 100.370 218.380 102.950 218.785 ;
        RECT 104.050 218.380 106.630 218.785 ;
        RECT 100.370 217.700 106.630 218.380 ;
        RECT 107.730 217.700 110.310 218.785 ;
        RECT 100.370 216.340 110.310 217.700 ;
        RECT 111.410 216.340 113.990 218.785 ;
        RECT 115.090 216.340 117.670 218.785 ;
        RECT 118.770 216.340 121.350 218.785 ;
        RECT 96.690 215.520 121.350 216.340 ;
        RECT 96.690 214.980 97.440 215.520 ;
        RECT 93.010 199.340 97.440 214.980 ;
        RECT 89.330 198.660 97.440 199.340 ;
        RECT 23.040 29.680 97.440 198.660 ;
        RECT 99.840 214.980 121.350 215.520 ;
        RECT 122.450 214.980 125.030 218.785 ;
        RECT 99.840 213.620 125.030 214.980 ;
        RECT 126.130 214.980 128.710 218.785 ;
        RECT 129.810 218.380 132.390 218.785 ;
        RECT 133.490 218.380 136.070 218.785 ;
        RECT 129.810 214.980 136.070 218.380 ;
        RECT 137.170 217.020 139.750 218.785 ;
        RECT 140.850 217.020 143.430 218.785 ;
        RECT 137.170 216.340 143.430 217.020 ;
        RECT 144.530 216.340 147.110 218.785 ;
        RECT 137.170 214.980 147.110 216.340 ;
        RECT 148.210 218.380 150.790 218.785 ;
        RECT 151.890 218.380 154.470 218.785 ;
        RECT 148.210 217.020 154.470 218.380 ;
        RECT 155.570 217.020 158.150 218.785 ;
        RECT 148.210 214.980 158.150 217.020 ;
        RECT 126.130 213.620 158.150 214.980 ;
        RECT 99.840 206.450 158.150 213.620 ;
        RECT 159.250 215.520 626.625 218.785 ;
        RECT 159.250 206.450 174.240 215.520 ;
        RECT 99.840 29.680 174.240 206.450 ;
        RECT 176.640 136.140 251.040 215.520 ;
        RECT 253.440 136.140 327.840 215.520 ;
        RECT 330.240 136.140 404.640 215.520 ;
        RECT 407.040 136.140 481.440 215.520 ;
        RECT 483.840 136.140 558.240 215.520 ;
        RECT 560.640 136.140 626.625 215.520 ;
        RECT 176.640 29.780 626.625 136.140 ;
        RECT 176.640 29.680 251.040 29.780 ;
        RECT 253.440 29.680 327.840 29.780 ;
        RECT 330.240 29.680 404.640 29.780 ;
        RECT 407.040 29.680 481.440 29.780 ;
        RECT 483.840 29.680 558.240 29.780 ;
        RECT 560.640 29.680 626.625 29.780 ;
  END
END tt_um_urish_dffram
END LIBRARY

