VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    PORT
      LAYER met3 ;
        RECT 2917.600 1431.820 2924.800 1433.020 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    PORT
      LAYER met2 ;
        RECT 2228.190 3517.600 2228.750 3524.800 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    PORT
      LAYER met2 ;
        RECT 1904.350 3517.600 1904.910 3524.800 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    PORT
      LAYER met2 ;
        RECT 1580.510 3517.600 1581.070 3524.800 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    PORT
      LAYER met2 ;
        RECT 1256.670 3517.600 1257.230 3524.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    PORT
      LAYER met2 ;
        RECT 932.830 3517.600 933.390 3524.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    PORT
      LAYER met2 ;
        RECT 608.990 3517.600 609.550 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    PORT
      LAYER met2 ;
        RECT 285.150 3517.600 285.710 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    PORT
      LAYER met3 ;
        RECT -4.800 3435.100 2.400 3436.300 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    PORT
      LAYER met3 ;
        RECT -4.800 3182.140 2.400 3183.340 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    PORT
      LAYER met3 ;
        RECT -4.800 2929.180 2.400 2930.380 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 1692.940 2924.800 1694.140 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    PORT
      LAYER met3 ;
        RECT -4.800 2676.220 2.400 2677.420 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    PORT
      LAYER met3 ;
        RECT -4.800 2423.260 2.400 2424.460 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    PORT
      LAYER met3 ;
        RECT -4.800 2170.300 2.400 2171.500 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    PORT
      LAYER met3 ;
        RECT -4.800 1917.340 2.400 1918.540 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    PORT
      LAYER met3 ;
        RECT -4.800 1664.380 2.400 1665.580 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    PORT
      LAYER met3 ;
        RECT -4.800 1411.420 2.400 1412.620 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    PORT
      LAYER met3 ;
        RECT -4.800 1158.460 2.400 1159.660 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    PORT
      LAYER met3 ;
        RECT -4.800 905.500 2.400 906.700 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    PORT
      LAYER met3 ;
        RECT -4.800 652.540 2.400 653.740 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    PORT
      LAYER met3 ;
        RECT 2917.600 1954.060 2924.800 1955.260 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    PORT
      LAYER met3 ;
        RECT 2917.600 2215.180 2924.800 2216.380 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    PORT
      LAYER met3 ;
        RECT 2917.600 2476.300 2924.800 2477.500 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    PORT
      LAYER met3 ;
        RECT 2917.600 2737.420 2924.800 2738.620 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 2998.540 2924.800 2999.740 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    PORT
      LAYER met3 ;
        RECT 2917.600 3259.660 2924.800 3260.860 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    PORT
      LAYER met2 ;
        RECT 2875.870 3517.600 2876.430 3524.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    PORT
      LAYER met2 ;
        RECT 2552.030 3517.600 2552.590 3524.800 ;
    END
  END analog_io[9]
  PIN io_in[0]
    PORT
      LAYER met3 ;
        RECT 2917.600 60.940 2924.800 62.140 ;
    END
  END io_in[0]
  PIN io_in[10]
    PORT
      LAYER met3 ;
        RECT 2917.600 2280.460 2924.800 2281.660 ;
    END
  END io_in[10]
  PIN io_in[11]
    PORT
      LAYER met3 ;
        RECT 2917.600 2541.580 2924.800 2542.780 ;
    END
  END io_in[11]
  PIN io_in[12]
    PORT
      LAYER met3 ;
        RECT 2917.600 2802.700 2924.800 2803.900 ;
    END
  END io_in[12]
  PIN io_in[13]
    PORT
      LAYER met3 ;
        RECT 2917.600 3063.820 2924.800 3065.020 ;
    END
  END io_in[13]
  PIN io_in[14]
    PORT
      LAYER met3 ;
        RECT 2917.600 3324.940 2924.800 3326.140 ;
    END
  END io_in[14]
  PIN io_in[15]
    PORT
      LAYER met2 ;
        RECT 2794.910 3517.600 2795.470 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    PORT
      LAYER met2 ;
        RECT 2471.070 3517.600 2471.630 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    PORT
      LAYER met2 ;
        RECT 2147.230 3517.600 2147.790 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    PORT
      LAYER met2 ;
        RECT 1823.390 3517.600 1823.950 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    PORT
      LAYER met2 ;
        RECT 1499.550 3517.600 1500.110 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 256.780 2924.800 257.980 ;
    END
  END io_in[1]
  PIN io_in[20]
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    PORT
      LAYER met2 ;
        RECT 851.870 3517.600 852.430 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    PORT
      LAYER met2 ;
        RECT 528.030 3517.600 528.590 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    PORT
      LAYER met2 ;
        RECT 204.190 3517.600 204.750 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    PORT
      LAYER met3 ;
        RECT -4.800 3371.860 2.400 3373.060 ;
    END
  END io_in[24]
  PIN io_in[25]
    PORT
      LAYER met3 ;
        RECT -4.800 3118.900 2.400 3120.100 ;
    END
  END io_in[25]
  PIN io_in[26]
    PORT
      LAYER met3 ;
        RECT -4.800 2865.940 2.400 2867.140 ;
    END
  END io_in[26]
  PIN io_in[27]
    PORT
      LAYER met3 ;
        RECT -4.800 2612.980 2.400 2614.180 ;
    END
  END io_in[27]
  PIN io_in[28]
    PORT
      LAYER met3 ;
        RECT -4.800 2360.020 2.400 2361.220 ;
    END
  END io_in[28]
  PIN io_in[29]
    PORT
      LAYER met3 ;
        RECT -4.800 2107.060 2.400 2108.260 ;
    END
  END io_in[29]
  PIN io_in[2]
    PORT
      LAYER met3 ;
        RECT 2917.600 452.620 2924.800 453.820 ;
    END
  END io_in[2]
  PIN io_in[30]
    PORT
      LAYER met3 ;
        RECT -4.800 1854.100 2.400 1855.300 ;
    END
  END io_in[30]
  PIN io_in[31]
    PORT
      LAYER met3 ;
        RECT -4.800 1601.140 2.400 1602.340 ;
    END
  END io_in[31]
  PIN io_in[32]
    PORT
      LAYER met3 ;
        RECT -4.800 1348.180 2.400 1349.380 ;
    END
  END io_in[32]
  PIN io_in[33]
    PORT
      LAYER met3 ;
        RECT -4.800 1095.220 2.400 1096.420 ;
    END
  END io_in[33]
  PIN io_in[34]
    PORT
      LAYER met3 ;
        RECT -4.800 842.260 2.400 843.460 ;
    END
  END io_in[34]
  PIN io_in[35]
    PORT
      LAYER met3 ;
        RECT -4.800 589.300 2.400 590.500 ;
    END
  END io_in[35]
  PIN io_in[36]
    PORT
      LAYER met3 ;
        RECT -4.800 399.580 2.400 400.780 ;
    END
  END io_in[36]
  PIN io_in[37]
    PORT
      LAYER met3 ;
        RECT -4.800 209.860 2.400 211.060 ;
    END
  END io_in[37]
  PIN io_in[3]
    PORT
      LAYER met3 ;
        RECT 2917.600 648.460 2924.800 649.660 ;
    END
  END io_in[3]
  PIN io_in[4]
    PORT
      LAYER met3 ;
        RECT 2917.600 844.300 2924.800 845.500 ;
    END
  END io_in[4]
  PIN io_in[5]
    PORT
      LAYER met3 ;
        RECT 2917.600 1040.140 2924.800 1041.340 ;
    END
  END io_in[5]
  PIN io_in[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 1235.980 2924.800 1237.180 ;
    END
  END io_in[6]
  PIN io_in[7]
    PORT
      LAYER met3 ;
        RECT 2917.600 1497.100 2924.800 1498.300 ;
    END
  END io_in[7]
  PIN io_in[8]
    PORT
      LAYER met3 ;
        RECT 2917.600 1758.220 2924.800 1759.420 ;
    END
  END io_in[8]
  PIN io_in[9]
    PORT
      LAYER met3 ;
        RECT 2917.600 2019.340 2924.800 2020.540 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    PORT
      LAYER met3 ;
        RECT 2917.600 191.500 2924.800 192.700 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    PORT
      LAYER met3 ;
        RECT 2917.600 2411.020 2924.800 2412.220 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    PORT
      LAYER met3 ;
        RECT 2917.600 2672.140 2924.800 2673.340 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    PORT
      LAYER met3 ;
        RECT 2917.600 2933.260 2924.800 2934.460 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    PORT
      LAYER met3 ;
        RECT 2917.600 3194.380 2924.800 3195.580 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    PORT
      LAYER met3 ;
        RECT 2917.600 3455.500 2924.800 3456.700 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    PORT
      LAYER met2 ;
        RECT 2632.990 3517.600 2633.550 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    PORT
      LAYER met2 ;
        RECT 2309.150 3517.600 2309.710 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    PORT
      LAYER met2 ;
        RECT 1985.310 3517.600 1985.870 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    PORT
      LAYER met2 ;
        RECT 1661.470 3517.600 1662.030 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    PORT
      LAYER met2 ;
        RECT 1337.630 3517.600 1338.190 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 387.340 2924.800 388.540 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    PORT
      LAYER met2 ;
        RECT 689.950 3517.600 690.510 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    PORT
      LAYER met2 ;
        RECT 366.110 3517.600 366.670 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    PORT
      LAYER met2 ;
        RECT 42.270 3517.600 42.830 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    PORT
      LAYER met3 ;
        RECT -4.800 3245.380 2.400 3246.580 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    PORT
      LAYER met3 ;
        RECT -4.800 2992.420 2.400 2993.620 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    PORT
      LAYER met3 ;
        RECT -4.800 2739.460 2.400 2740.660 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    PORT
      LAYER met3 ;
        RECT -4.800 2486.500 2.400 2487.700 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    PORT
      LAYER met3 ;
        RECT -4.800 2233.540 2.400 2234.740 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    PORT
      LAYER met3 ;
        RECT -4.800 1980.580 2.400 1981.780 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    PORT
      LAYER met3 ;
        RECT 2917.600 583.180 2924.800 584.380 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    PORT
      LAYER met3 ;
        RECT -4.800 1727.620 2.400 1728.820 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    PORT
      LAYER met3 ;
        RECT -4.800 1474.660 2.400 1475.860 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    PORT
      LAYER met3 ;
        RECT -4.800 1221.700 2.400 1222.900 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    PORT
      LAYER met3 ;
        RECT -4.800 968.740 2.400 969.940 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    PORT
      LAYER met3 ;
        RECT -4.800 715.780 2.400 716.980 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    PORT
      LAYER met3 ;
        RECT -4.800 462.820 2.400 464.020 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    PORT
      LAYER met3 ;
        RECT -4.800 273.100 2.400 274.300 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    PORT
      LAYER met3 ;
        RECT -4.800 83.380 2.400 84.580 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    PORT
      LAYER met3 ;
        RECT 2917.600 779.020 2924.800 780.220 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    PORT
      LAYER met3 ;
        RECT 2917.600 974.860 2924.800 976.060 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    PORT
      LAYER met3 ;
        RECT 2917.600 1170.700 2924.800 1171.900 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 1366.540 2924.800 1367.740 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    PORT
      LAYER met3 ;
        RECT 2917.600 1627.660 2924.800 1628.860 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    PORT
      LAYER met3 ;
        RECT 2917.600 1888.780 2924.800 1889.980 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    PORT
      LAYER met3 ;
        RECT 2917.600 2149.900 2924.800 2151.100 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    PORT
      LAYER met3 ;
        RECT 2917.600 126.220 2924.800 127.420 ;
    END
  END io_out[0]
  PIN io_out[10]
    PORT
      LAYER met3 ;
        RECT 2917.600 2345.740 2924.800 2346.940 ;
    END
  END io_out[10]
  PIN io_out[11]
    PORT
      LAYER met3 ;
        RECT 2917.600 2606.860 2924.800 2608.060 ;
    END
  END io_out[11]
  PIN io_out[12]
    PORT
      LAYER met3 ;
        RECT 2917.600 2867.980 2924.800 2869.180 ;
    END
  END io_out[12]
  PIN io_out[13]
    PORT
      LAYER met3 ;
        RECT 2917.600 3129.100 2924.800 3130.300 ;
    END
  END io_out[13]
  PIN io_out[14]
    PORT
      LAYER met3 ;
        RECT 2917.600 3390.220 2924.800 3391.420 ;
    END
  END io_out[14]
  PIN io_out[15]
    PORT
      LAYER met2 ;
        RECT 2713.950 3517.600 2714.510 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    PORT
      LAYER met2 ;
        RECT 2390.110 3517.600 2390.670 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    PORT
      LAYER met2 ;
        RECT 2066.270 3517.600 2066.830 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    PORT
      LAYER met2 ;
        RECT 1742.430 3517.600 1742.990 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    PORT
      LAYER met2 ;
        RECT 1418.590 3517.600 1419.150 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 322.060 2924.800 323.260 ;
    END
  END io_out[1]
  PIN io_out[20]
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    PORT
      LAYER met2 ;
        RECT 770.910 3517.600 771.470 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    PORT
      LAYER met2 ;
        RECT 447.070 3517.600 447.630 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    PORT
      LAYER met2 ;
        RECT 123.230 3517.600 123.790 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    PORT
      LAYER met3 ;
        RECT -4.800 3308.620 2.400 3309.820 ;
    END
  END io_out[24]
  PIN io_out[25]
    PORT
      LAYER met3 ;
        RECT -4.800 3055.660 2.400 3056.860 ;
    END
  END io_out[25]
  PIN io_out[26]
    PORT
      LAYER met3 ;
        RECT -4.800 2802.700 2.400 2803.900 ;
    END
  END io_out[26]
  PIN io_out[27]
    PORT
      LAYER met3 ;
        RECT -4.800 2549.740 2.400 2550.940 ;
    END
  END io_out[27]
  PIN io_out[28]
    PORT
      LAYER met3 ;
        RECT -4.800 2296.780 2.400 2297.980 ;
    END
  END io_out[28]
  PIN io_out[29]
    PORT
      LAYER met3 ;
        RECT -4.800 2043.820 2.400 2045.020 ;
    END
  END io_out[29]
  PIN io_out[2]
    PORT
      LAYER met3 ;
        RECT 2917.600 517.900 2924.800 519.100 ;
    END
  END io_out[2]
  PIN io_out[30]
    PORT
      LAYER met3 ;
        RECT -4.800 1790.860 2.400 1792.060 ;
    END
  END io_out[30]
  PIN io_out[31]
    PORT
      LAYER met3 ;
        RECT -4.800 1537.900 2.400 1539.100 ;
    END
  END io_out[31]
  PIN io_out[32]
    PORT
      LAYER met3 ;
        RECT -4.800 1284.940 2.400 1286.140 ;
    END
  END io_out[32]
  PIN io_out[33]
    PORT
      LAYER met3 ;
        RECT -4.800 1031.980 2.400 1033.180 ;
    END
  END io_out[33]
  PIN io_out[34]
    PORT
      LAYER met3 ;
        RECT -4.800 779.020 2.400 780.220 ;
    END
  END io_out[34]
  PIN io_out[35]
    PORT
      LAYER met3 ;
        RECT -4.800 526.060 2.400 527.260 ;
    END
  END io_out[35]
  PIN io_out[36]
    PORT
      LAYER met3 ;
        RECT -4.800 336.340 2.400 337.540 ;
    END
  END io_out[36]
  PIN io_out[37]
    PORT
      LAYER met3 ;
        RECT -4.800 146.620 2.400 147.820 ;
    END
  END io_out[37]
  PIN io_out[3]
    PORT
      LAYER met3 ;
        RECT 2917.600 713.740 2924.800 714.940 ;
    END
  END io_out[3]
  PIN io_out[4]
    PORT
      LAYER met3 ;
        RECT 2917.600 909.580 2924.800 910.780 ;
    END
  END io_out[4]
  PIN io_out[5]
    PORT
      LAYER met3 ;
        RECT 2917.600 1105.420 2924.800 1106.620 ;
    END
  END io_out[5]
  PIN io_out[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 1301.260 2924.800 1302.460 ;
    END
  END io_out[6]
  PIN io_out[7]
    PORT
      LAYER met3 ;
        RECT 2917.600 1562.380 2924.800 1563.580 ;
    END
  END io_out[7]
  PIN io_out[8]
    PORT
      LAYER met3 ;
        RECT 2917.600 1823.500 2924.800 1824.700 ;
    END
  END io_out[8]
  PIN io_out[9]
    PORT
      LAYER met3 ;
        RECT 2917.600 2084.620 2924.800 2085.820 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    PORT
      LAYER met2 ;
        RECT 683.510 -4.800 684.070 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    PORT
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    PORT
      LAYER met2 ;
        RECT 2356.070 -4.800 2356.630 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    PORT
      LAYER met2 ;
        RECT 2372.630 -4.800 2373.190 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    PORT
      LAYER met2 ;
        RECT 2389.190 -4.800 2389.750 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    PORT
      LAYER met2 ;
        RECT 2405.750 -4.800 2406.310 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    PORT
      LAYER met2 ;
        RECT 2422.310 -4.800 2422.870 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    PORT
      LAYER met2 ;
        RECT 2438.870 -4.800 2439.430 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    PORT
      LAYER met2 ;
        RECT 2455.430 -4.800 2455.990 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    PORT
      LAYER met2 ;
        RECT 2471.990 -4.800 2472.550 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    PORT
      LAYER met2 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    PORT
      LAYER met2 ;
        RECT 849.110 -4.800 849.670 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    PORT
      LAYER met2 ;
        RECT 2505.110 -4.800 2505.670 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    PORT
      LAYER met2 ;
        RECT 2521.670 -4.800 2522.230 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    PORT
      LAYER met2 ;
        RECT 2538.230 -4.800 2538.790 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    PORT
      LAYER met2 ;
        RECT 2554.790 -4.800 2555.350 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    PORT
      LAYER met2 ;
        RECT 2571.350 -4.800 2571.910 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    PORT
      LAYER met2 ;
        RECT 2587.910 -4.800 2588.470 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    PORT
      LAYER met2 ;
        RECT 2604.470 -4.800 2605.030 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    PORT
      LAYER met2 ;
        RECT 2621.030 -4.800 2621.590 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    PORT
      LAYER met2 ;
        RECT 2637.590 -4.800 2638.150 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    PORT
      LAYER met2 ;
        RECT 2654.150 -4.800 2654.710 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    PORT
      LAYER met2 ;
        RECT 865.670 -4.800 866.230 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    PORT
      LAYER met2 ;
        RECT 2670.710 -4.800 2671.270 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    PORT
      LAYER met2 ;
        RECT 2687.270 -4.800 2687.830 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    PORT
      LAYER met2 ;
        RECT 2703.830 -4.800 2704.390 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    PORT
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    PORT
      LAYER met2 ;
        RECT 2736.950 -4.800 2737.510 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    PORT
      LAYER met2 ;
        RECT 2753.510 -4.800 2754.070 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    PORT
      LAYER met2 ;
        RECT 2770.070 -4.800 2770.630 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    PORT
      LAYER met2 ;
        RECT 2786.630 -4.800 2787.190 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    PORT
      LAYER met2 ;
        RECT 882.230 -4.800 882.790 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    PORT
      LAYER met2 ;
        RECT 898.790 -4.800 899.350 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    PORT
      LAYER met2 ;
        RECT 915.350 -4.800 915.910 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    PORT
      LAYER met2 ;
        RECT 931.910 -4.800 932.470 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    PORT
      LAYER met2 ;
        RECT 948.470 -4.800 949.030 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    PORT
      LAYER met2 ;
        RECT 965.030 -4.800 965.590 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    PORT
      LAYER met2 ;
        RECT 981.590 -4.800 982.150 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    PORT
      LAYER met2 ;
        RECT 998.150 -4.800 998.710 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    PORT
      LAYER met2 ;
        RECT 700.070 -4.800 700.630 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    PORT
      LAYER met2 ;
        RECT 1014.710 -4.800 1015.270 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    PORT
      LAYER met2 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    PORT
      LAYER met2 ;
        RECT 1047.830 -4.800 1048.390 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    PORT
      LAYER met2 ;
        RECT 1064.390 -4.800 1064.950 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    PORT
      LAYER met2 ;
        RECT 1080.950 -4.800 1081.510 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    PORT
      LAYER met2 ;
        RECT 1097.510 -4.800 1098.070 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    PORT
      LAYER met2 ;
        RECT 1114.070 -4.800 1114.630 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    PORT
      LAYER met2 ;
        RECT 1130.630 -4.800 1131.190 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    PORT
      LAYER met2 ;
        RECT 1147.190 -4.800 1147.750 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    PORT
      LAYER met2 ;
        RECT 1163.750 -4.800 1164.310 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    PORT
      LAYER met2 ;
        RECT 716.630 -4.800 717.190 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    PORT
      LAYER met2 ;
        RECT 1180.310 -4.800 1180.870 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    PORT
      LAYER met2 ;
        RECT 1196.870 -4.800 1197.430 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    PORT
      LAYER met2 ;
        RECT 1213.430 -4.800 1213.990 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    PORT
      LAYER met2 ;
        RECT 1229.990 -4.800 1230.550 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    PORT
      LAYER met2 ;
        RECT 1246.550 -4.800 1247.110 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    PORT
      LAYER met2 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    PORT
      LAYER met2 ;
        RECT 1279.670 -4.800 1280.230 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    PORT
      LAYER met2 ;
        RECT 1296.230 -4.800 1296.790 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    PORT
      LAYER met2 ;
        RECT 1312.790 -4.800 1313.350 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    PORT
      LAYER met2 ;
        RECT 1329.350 -4.800 1329.910 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    PORT
      LAYER met2 ;
        RECT 733.190 -4.800 733.750 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    PORT
      LAYER met2 ;
        RECT 1345.910 -4.800 1346.470 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    PORT
      LAYER met2 ;
        RECT 1362.470 -4.800 1363.030 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    PORT
      LAYER met2 ;
        RECT 1379.030 -4.800 1379.590 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    PORT
      LAYER met2 ;
        RECT 1395.590 -4.800 1396.150 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    PORT
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    PORT
      LAYER met2 ;
        RECT 1428.710 -4.800 1429.270 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    PORT
      LAYER met2 ;
        RECT 1445.270 -4.800 1445.830 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    PORT
      LAYER met2 ;
        RECT 1461.830 -4.800 1462.390 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    PORT
      LAYER met2 ;
        RECT 1478.390 -4.800 1478.950 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    PORT
      LAYER met2 ;
        RECT 1494.950 -4.800 1495.510 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    PORT
      LAYER met2 ;
        RECT 749.750 -4.800 750.310 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    PORT
      LAYER met2 ;
        RECT 1511.510 -4.800 1512.070 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    PORT
      LAYER met2 ;
        RECT 1528.070 -4.800 1528.630 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    PORT
      LAYER met2 ;
        RECT 1544.630 -4.800 1545.190 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    PORT
      LAYER met2 ;
        RECT 1561.190 -4.800 1561.750 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    PORT
      LAYER met2 ;
        RECT 1577.750 -4.800 1578.310 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    PORT
      LAYER met2 ;
        RECT 1594.310 -4.800 1594.870 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    PORT
      LAYER met2 ;
        RECT 1610.870 -4.800 1611.430 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    PORT
      LAYER met2 ;
        RECT 1627.430 -4.800 1627.990 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    PORT
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    PORT
      LAYER met2 ;
        RECT 1660.550 -4.800 1661.110 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    PORT
      LAYER met2 ;
        RECT 766.310 -4.800 766.870 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    PORT
      LAYER met2 ;
        RECT 1677.110 -4.800 1677.670 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    PORT
      LAYER met2 ;
        RECT 1693.670 -4.800 1694.230 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    PORT
      LAYER met2 ;
        RECT 1710.230 -4.800 1710.790 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    PORT
      LAYER met2 ;
        RECT 1726.790 -4.800 1727.350 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    PORT
      LAYER met2 ;
        RECT 1743.350 -4.800 1743.910 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    PORT
      LAYER met2 ;
        RECT 1759.910 -4.800 1760.470 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    PORT
      LAYER met2 ;
        RECT 1776.470 -4.800 1777.030 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    PORT
      LAYER met2 ;
        RECT 1793.030 -4.800 1793.590 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    PORT
      LAYER met2 ;
        RECT 1809.590 -4.800 1810.150 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    PORT
      LAYER met2 ;
        RECT 1826.150 -4.800 1826.710 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    PORT
      LAYER met2 ;
        RECT 782.870 -4.800 783.430 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    PORT
      LAYER met2 ;
        RECT 1842.710 -4.800 1843.270 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    PORT
      LAYER met2 ;
        RECT 1859.270 -4.800 1859.830 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    PORT
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    PORT
      LAYER met2 ;
        RECT 1892.390 -4.800 1892.950 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    PORT
      LAYER met2 ;
        RECT 1908.950 -4.800 1909.510 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    PORT
      LAYER met2 ;
        RECT 1925.510 -4.800 1926.070 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    PORT
      LAYER met2 ;
        RECT 1942.070 -4.800 1942.630 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    PORT
      LAYER met2 ;
        RECT 1958.630 -4.800 1959.190 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    PORT
      LAYER met2 ;
        RECT 1975.190 -4.800 1975.750 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    PORT
      LAYER met2 ;
        RECT 1991.750 -4.800 1992.310 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    PORT
      LAYER met2 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    PORT
      LAYER met2 ;
        RECT 2008.310 -4.800 2008.870 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    PORT
      LAYER met2 ;
        RECT 2024.870 -4.800 2025.430 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    PORT
      LAYER met2 ;
        RECT 2041.430 -4.800 2041.990 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    PORT
      LAYER met2 ;
        RECT 2057.990 -4.800 2058.550 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    PORT
      LAYER met2 ;
        RECT 2074.550 -4.800 2075.110 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    PORT
      LAYER met2 ;
        RECT 2091.110 -4.800 2091.670 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    PORT
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    PORT
      LAYER met2 ;
        RECT 2124.230 -4.800 2124.790 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    PORT
      LAYER met2 ;
        RECT 2140.790 -4.800 2141.350 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    PORT
      LAYER met2 ;
        RECT 2157.350 -4.800 2157.910 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    PORT
      LAYER met2 ;
        RECT 815.990 -4.800 816.550 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    PORT
      LAYER met2 ;
        RECT 2173.910 -4.800 2174.470 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    PORT
      LAYER met2 ;
        RECT 2190.470 -4.800 2191.030 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    PORT
      LAYER met2 ;
        RECT 2207.030 -4.800 2207.590 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    PORT
      LAYER met2 ;
        RECT 2223.590 -4.800 2224.150 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    PORT
      LAYER met2 ;
        RECT 2240.150 -4.800 2240.710 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    PORT
      LAYER met2 ;
        RECT 2256.710 -4.800 2257.270 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    PORT
      LAYER met2 ;
        RECT 2273.270 -4.800 2273.830 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    PORT
      LAYER met2 ;
        RECT 2289.830 -4.800 2290.390 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    PORT
      LAYER met2 ;
        RECT 2306.390 -4.800 2306.950 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    PORT
      LAYER met2 ;
        RECT 2322.950 -4.800 2323.510 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    PORT
      LAYER met2 ;
        RECT 832.550 -4.800 833.110 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    PORT
      LAYER met2 ;
        RECT 689.030 -4.800 689.590 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    PORT
      LAYER met2 ;
        RECT 2345.030 -4.800 2345.590 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    PORT
      LAYER met2 ;
        RECT 2361.590 -4.800 2362.150 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    PORT
      LAYER met2 ;
        RECT 2378.150 -4.800 2378.710 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    PORT
      LAYER met2 ;
        RECT 2394.710 -4.800 2395.270 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    PORT
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    PORT
      LAYER met2 ;
        RECT 2427.830 -4.800 2428.390 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    PORT
      LAYER met2 ;
        RECT 2444.390 -4.800 2444.950 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    PORT
      LAYER met2 ;
        RECT 2460.950 -4.800 2461.510 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    PORT
      LAYER met2 ;
        RECT 2477.510 -4.800 2478.070 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    PORT
      LAYER met2 ;
        RECT 2494.070 -4.800 2494.630 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    PORT
      LAYER met2 ;
        RECT 854.630 -4.800 855.190 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    PORT
      LAYER met2 ;
        RECT 2510.630 -4.800 2511.190 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    PORT
      LAYER met2 ;
        RECT 2527.190 -4.800 2527.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    PORT
      LAYER met2 ;
        RECT 2543.750 -4.800 2544.310 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    PORT
      LAYER met2 ;
        RECT 2560.310 -4.800 2560.870 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    PORT
      LAYER met2 ;
        RECT 2576.870 -4.800 2577.430 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    PORT
      LAYER met2 ;
        RECT 2593.430 -4.800 2593.990 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    PORT
      LAYER met2 ;
        RECT 2609.990 -4.800 2610.550 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    PORT
      LAYER met2 ;
        RECT 2626.550 -4.800 2627.110 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    PORT
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    PORT
      LAYER met2 ;
        RECT 2659.670 -4.800 2660.230 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    PORT
      LAYER met2 ;
        RECT 871.190 -4.800 871.750 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    PORT
      LAYER met2 ;
        RECT 2676.230 -4.800 2676.790 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    PORT
      LAYER met2 ;
        RECT 2692.790 -4.800 2693.350 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    PORT
      LAYER met2 ;
        RECT 2709.350 -4.800 2709.910 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    PORT
      LAYER met2 ;
        RECT 2725.910 -4.800 2726.470 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    PORT
      LAYER met2 ;
        RECT 2742.470 -4.800 2743.030 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    PORT
      LAYER met2 ;
        RECT 2759.030 -4.800 2759.590 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    PORT
      LAYER met2 ;
        RECT 2775.590 -4.800 2776.150 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    PORT
      LAYER met2 ;
        RECT 2792.150 -4.800 2792.710 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    PORT
      LAYER met2 ;
        RECT 887.750 -4.800 888.310 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    PORT
      LAYER met2 ;
        RECT 904.310 -4.800 904.870 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    PORT
      LAYER met2 ;
        RECT 920.870 -4.800 921.430 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    PORT
      LAYER met2 ;
        RECT 937.430 -4.800 937.990 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    PORT
      LAYER met2 ;
        RECT 970.550 -4.800 971.110 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    PORT
      LAYER met2 ;
        RECT 987.110 -4.800 987.670 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    PORT
      LAYER met2 ;
        RECT 1003.670 -4.800 1004.230 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    PORT
      LAYER met2 ;
        RECT 705.590 -4.800 706.150 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    PORT
      LAYER met2 ;
        RECT 1020.230 -4.800 1020.790 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    PORT
      LAYER met2 ;
        RECT 1036.790 -4.800 1037.350 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    PORT
      LAYER met2 ;
        RECT 1053.350 -4.800 1053.910 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    PORT
      LAYER met2 ;
        RECT 1069.910 -4.800 1070.470 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    PORT
      LAYER met2 ;
        RECT 1086.470 -4.800 1087.030 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    PORT
      LAYER met2 ;
        RECT 1103.030 -4.800 1103.590 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    PORT
      LAYER met2 ;
        RECT 1119.590 -4.800 1120.150 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    PORT
      LAYER met2 ;
        RECT 1136.150 -4.800 1136.710 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    PORT
      LAYER met2 ;
        RECT 1152.710 -4.800 1153.270 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    PORT
      LAYER met2 ;
        RECT 1169.270 -4.800 1169.830 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    PORT
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    PORT
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    PORT
      LAYER met2 ;
        RECT 1202.390 -4.800 1202.950 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    PORT
      LAYER met2 ;
        RECT 1218.950 -4.800 1219.510 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    PORT
      LAYER met2 ;
        RECT 1235.510 -4.800 1236.070 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    PORT
      LAYER met2 ;
        RECT 1252.070 -4.800 1252.630 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    PORT
      LAYER met2 ;
        RECT 1268.630 -4.800 1269.190 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    PORT
      LAYER met2 ;
        RECT 1285.190 -4.800 1285.750 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    PORT
      LAYER met2 ;
        RECT 1301.750 -4.800 1302.310 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    PORT
      LAYER met2 ;
        RECT 1318.310 -4.800 1318.870 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    PORT
      LAYER met2 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    PORT
      LAYER met2 ;
        RECT 738.710 -4.800 739.270 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    PORT
      LAYER met2 ;
        RECT 1351.430 -4.800 1351.990 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    PORT
      LAYER met2 ;
        RECT 1367.990 -4.800 1368.550 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    PORT
      LAYER met2 ;
        RECT 1384.550 -4.800 1385.110 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    PORT
      LAYER met2 ;
        RECT 1401.110 -4.800 1401.670 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    PORT
      LAYER met2 ;
        RECT 1417.670 -4.800 1418.230 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    PORT
      LAYER met2 ;
        RECT 1434.230 -4.800 1434.790 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    PORT
      LAYER met2 ;
        RECT 1450.790 -4.800 1451.350 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    PORT
      LAYER met2 ;
        RECT 1467.350 -4.800 1467.910 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    PORT
      LAYER met2 ;
        RECT 1483.910 -4.800 1484.470 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    PORT
      LAYER met2 ;
        RECT 1500.470 -4.800 1501.030 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    PORT
      LAYER met2 ;
        RECT 755.270 -4.800 755.830 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    PORT
      LAYER met2 ;
        RECT 1517.030 -4.800 1517.590 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    PORT
      LAYER met2 ;
        RECT 1533.590 -4.800 1534.150 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    PORT
      LAYER met2 ;
        RECT 1550.150 -4.800 1550.710 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    PORT
      LAYER met2 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    PORT
      LAYER met2 ;
        RECT 1583.270 -4.800 1583.830 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    PORT
      LAYER met2 ;
        RECT 1599.830 -4.800 1600.390 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    PORT
      LAYER met2 ;
        RECT 1616.390 -4.800 1616.950 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    PORT
      LAYER met2 ;
        RECT 1632.950 -4.800 1633.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    PORT
      LAYER met2 ;
        RECT 1649.510 -4.800 1650.070 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    PORT
      LAYER met2 ;
        RECT 1666.070 -4.800 1666.630 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    PORT
      LAYER met2 ;
        RECT 771.830 -4.800 772.390 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    PORT
      LAYER met2 ;
        RECT 1682.630 -4.800 1683.190 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    PORT
      LAYER met2 ;
        RECT 1699.190 -4.800 1699.750 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    PORT
      LAYER met2 ;
        RECT 1715.750 -4.800 1716.310 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    PORT
      LAYER met2 ;
        RECT 1732.310 -4.800 1732.870 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    PORT
      LAYER met2 ;
        RECT 1748.870 -4.800 1749.430 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    PORT
      LAYER met2 ;
        RECT 1765.430 -4.800 1765.990 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    PORT
      LAYER met2 ;
        RECT 1781.990 -4.800 1782.550 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    PORT
      LAYER met2 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    PORT
      LAYER met2 ;
        RECT 1815.110 -4.800 1815.670 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    PORT
      LAYER met2 ;
        RECT 1831.670 -4.800 1832.230 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    PORT
      LAYER met2 ;
        RECT 788.390 -4.800 788.950 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    PORT
      LAYER met2 ;
        RECT 1848.230 -4.800 1848.790 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    PORT
      LAYER met2 ;
        RECT 1864.790 -4.800 1865.350 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    PORT
      LAYER met2 ;
        RECT 1881.350 -4.800 1881.910 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    PORT
      LAYER met2 ;
        RECT 1897.910 -4.800 1898.470 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    PORT
      LAYER met2 ;
        RECT 1914.470 -4.800 1915.030 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    PORT
      LAYER met2 ;
        RECT 1931.030 -4.800 1931.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    PORT
      LAYER met2 ;
        RECT 1947.590 -4.800 1948.150 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    PORT
      LAYER met2 ;
        RECT 1964.150 -4.800 1964.710 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    PORT
      LAYER met2 ;
        RECT 1980.710 -4.800 1981.270 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    PORT
      LAYER met2 ;
        RECT 1997.270 -4.800 1997.830 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    PORT
      LAYER met2 ;
        RECT 804.950 -4.800 805.510 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    PORT
      LAYER met2 ;
        RECT 2013.830 -4.800 2014.390 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    PORT
      LAYER met2 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    PORT
      LAYER met2 ;
        RECT 2046.950 -4.800 2047.510 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    PORT
      LAYER met2 ;
        RECT 2063.510 -4.800 2064.070 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    PORT
      LAYER met2 ;
        RECT 2080.070 -4.800 2080.630 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    PORT
      LAYER met2 ;
        RECT 2096.630 -4.800 2097.190 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    PORT
      LAYER met2 ;
        RECT 2113.190 -4.800 2113.750 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    PORT
      LAYER met2 ;
        RECT 2129.750 -4.800 2130.310 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    PORT
      LAYER met2 ;
        RECT 2146.310 -4.800 2146.870 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    PORT
      LAYER met2 ;
        RECT 2162.870 -4.800 2163.430 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    PORT
      LAYER met2 ;
        RECT 821.510 -4.800 822.070 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    PORT
      LAYER met2 ;
        RECT 2179.430 -4.800 2179.990 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    PORT
      LAYER met2 ;
        RECT 2195.990 -4.800 2196.550 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    PORT
      LAYER met2 ;
        RECT 2212.550 -4.800 2213.110 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    PORT
      LAYER met2 ;
        RECT 2229.110 -4.800 2229.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    PORT
      LAYER met2 ;
        RECT 2245.670 -4.800 2246.230 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    PORT
      LAYER met2 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    PORT
      LAYER met2 ;
        RECT 2278.790 -4.800 2279.350 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    PORT
      LAYER met2 ;
        RECT 2295.350 -4.800 2295.910 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    PORT
      LAYER met2 ;
        RECT 2311.910 -4.800 2312.470 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    PORT
      LAYER met2 ;
        RECT 2328.470 -4.800 2329.030 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    PORT
      LAYER met2 ;
        RECT 838.070 -4.800 838.630 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    PORT
      LAYER met2 ;
        RECT 694.550 -4.800 695.110 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    PORT
      LAYER met2 ;
        RECT 2350.550 -4.800 2351.110 2.400 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    PORT
      LAYER met2 ;
        RECT 2367.110 -4.800 2367.670 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    PORT
      LAYER met2 ;
        RECT 2383.670 -4.800 2384.230 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    PORT
      LAYER met2 ;
        RECT 2400.230 -4.800 2400.790 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    PORT
      LAYER met2 ;
        RECT 2416.790 -4.800 2417.350 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    PORT
      LAYER met2 ;
        RECT 2433.350 -4.800 2433.910 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    PORT
      LAYER met2 ;
        RECT 2449.910 -4.800 2450.470 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    PORT
      LAYER met2 ;
        RECT 2466.470 -4.800 2467.030 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    PORT
      LAYER met2 ;
        RECT 2483.030 -4.800 2483.590 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    PORT
      LAYER met2 ;
        RECT 2499.590 -4.800 2500.150 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    PORT
      LAYER met2 ;
        RECT 860.150 -4.800 860.710 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    PORT
      LAYER met2 ;
        RECT 2516.150 -4.800 2516.710 2.400 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    PORT
      LAYER met2 ;
        RECT 2532.710 -4.800 2533.270 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    PORT
      LAYER met2 ;
        RECT 2549.270 -4.800 2549.830 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    PORT
      LAYER met2 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    PORT
      LAYER met2 ;
        RECT 2582.390 -4.800 2582.950 2.400 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    PORT
      LAYER met2 ;
        RECT 2598.950 -4.800 2599.510 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    PORT
      LAYER met2 ;
        RECT 2615.510 -4.800 2616.070 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    PORT
      LAYER met2 ;
        RECT 2632.070 -4.800 2632.630 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    PORT
      LAYER met2 ;
        RECT 2648.630 -4.800 2649.190 2.400 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    PORT
      LAYER met2 ;
        RECT 2665.190 -4.800 2665.750 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    PORT
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    PORT
      LAYER met2 ;
        RECT 2681.750 -4.800 2682.310 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    PORT
      LAYER met2 ;
        RECT 2698.310 -4.800 2698.870 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    PORT
      LAYER met2 ;
        RECT 2714.870 -4.800 2715.430 2.400 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    PORT
      LAYER met2 ;
        RECT 2731.430 -4.800 2731.990 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    PORT
      LAYER met2 ;
        RECT 2747.990 -4.800 2748.550 2.400 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    PORT
      LAYER met2 ;
        RECT 2764.550 -4.800 2765.110 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    PORT
      LAYER met2 ;
        RECT 2781.110 -4.800 2781.670 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    PORT
      LAYER met2 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    PORT
      LAYER met2 ;
        RECT 893.270 -4.800 893.830 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    PORT
      LAYER met2 ;
        RECT 909.830 -4.800 910.390 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    PORT
      LAYER met2 ;
        RECT 926.390 -4.800 926.950 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    PORT
      LAYER met2 ;
        RECT 942.950 -4.800 943.510 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    PORT
      LAYER met2 ;
        RECT 959.510 -4.800 960.070 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    PORT
      LAYER met2 ;
        RECT 976.070 -4.800 976.630 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    PORT
      LAYER met2 ;
        RECT 992.630 -4.800 993.190 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    PORT
      LAYER met2 ;
        RECT 1009.190 -4.800 1009.750 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    PORT
      LAYER met2 ;
        RECT 711.110 -4.800 711.670 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    PORT
      LAYER met2 ;
        RECT 1025.750 -4.800 1026.310 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    PORT
      LAYER met2 ;
        RECT 1042.310 -4.800 1042.870 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    PORT
      LAYER met2 ;
        RECT 1058.870 -4.800 1059.430 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    PORT
      LAYER met2 ;
        RECT 1075.430 -4.800 1075.990 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    PORT
      LAYER met2 ;
        RECT 1091.990 -4.800 1092.550 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    PORT
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    PORT
      LAYER met2 ;
        RECT 1125.110 -4.800 1125.670 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    PORT
      LAYER met2 ;
        RECT 1141.670 -4.800 1142.230 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    PORT
      LAYER met2 ;
        RECT 1158.230 -4.800 1158.790 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    PORT
      LAYER met2 ;
        RECT 1174.790 -4.800 1175.350 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    PORT
      LAYER met2 ;
        RECT 727.670 -4.800 728.230 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    PORT
      LAYER met2 ;
        RECT 1191.350 -4.800 1191.910 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    PORT
      LAYER met2 ;
        RECT 1207.910 -4.800 1208.470 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    PORT
      LAYER met2 ;
        RECT 1224.470 -4.800 1225.030 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    PORT
      LAYER met2 ;
        RECT 1241.030 -4.800 1241.590 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    PORT
      LAYER met2 ;
        RECT 1257.590 -4.800 1258.150 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    PORT
      LAYER met2 ;
        RECT 1274.150 -4.800 1274.710 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    PORT
      LAYER met2 ;
        RECT 1290.710 -4.800 1291.270 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    PORT
      LAYER met2 ;
        RECT 1307.270 -4.800 1307.830 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    PORT
      LAYER met2 ;
        RECT 1323.830 -4.800 1324.390 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    PORT
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    PORT
      LAYER met2 ;
        RECT 744.230 -4.800 744.790 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    PORT
      LAYER met2 ;
        RECT 1356.950 -4.800 1357.510 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    PORT
      LAYER met2 ;
        RECT 1373.510 -4.800 1374.070 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    PORT
      LAYER met2 ;
        RECT 1390.070 -4.800 1390.630 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    PORT
      LAYER met2 ;
        RECT 1406.630 -4.800 1407.190 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    PORT
      LAYER met2 ;
        RECT 1423.190 -4.800 1423.750 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    PORT
      LAYER met2 ;
        RECT 1439.750 -4.800 1440.310 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    PORT
      LAYER met2 ;
        RECT 1456.310 -4.800 1456.870 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    PORT
      LAYER met2 ;
        RECT 1472.870 -4.800 1473.430 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    PORT
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    PORT
      LAYER met2 ;
        RECT 1505.990 -4.800 1506.550 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    PORT
      LAYER met2 ;
        RECT 760.790 -4.800 761.350 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    PORT
      LAYER met2 ;
        RECT 1522.550 -4.800 1523.110 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    PORT
      LAYER met2 ;
        RECT 1539.110 -4.800 1539.670 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    PORT
      LAYER met2 ;
        RECT 1555.670 -4.800 1556.230 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    PORT
      LAYER met2 ;
        RECT 1572.230 -4.800 1572.790 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    PORT
      LAYER met2 ;
        RECT 1588.790 -4.800 1589.350 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    PORT
      LAYER met2 ;
        RECT 1605.350 -4.800 1605.910 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    PORT
      LAYER met2 ;
        RECT 1621.910 -4.800 1622.470 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    PORT
      LAYER met2 ;
        RECT 1638.470 -4.800 1639.030 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    PORT
      LAYER met2 ;
        RECT 1655.030 -4.800 1655.590 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    PORT
      LAYER met2 ;
        RECT 1671.590 -4.800 1672.150 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    PORT
      LAYER met2 ;
        RECT 777.350 -4.800 777.910 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    PORT
      LAYER met2 ;
        RECT 1688.150 -4.800 1688.710 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    PORT
      LAYER met2 ;
        RECT 1704.710 -4.800 1705.270 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    PORT
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    PORT
      LAYER met2 ;
        RECT 1737.830 -4.800 1738.390 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    PORT
      LAYER met2 ;
        RECT 1754.390 -4.800 1754.950 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    PORT
      LAYER met2 ;
        RECT 1770.950 -4.800 1771.510 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    PORT
      LAYER met2 ;
        RECT 1787.510 -4.800 1788.070 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    PORT
      LAYER met2 ;
        RECT 1804.070 -4.800 1804.630 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    PORT
      LAYER met2 ;
        RECT 1820.630 -4.800 1821.190 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    PORT
      LAYER met2 ;
        RECT 1837.190 -4.800 1837.750 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    PORT
      LAYER met2 ;
        RECT 793.910 -4.800 794.470 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    PORT
      LAYER met2 ;
        RECT 1853.750 -4.800 1854.310 2.400 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    PORT
      LAYER met2 ;
        RECT 1870.310 -4.800 1870.870 2.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    PORT
      LAYER met2 ;
        RECT 1886.870 -4.800 1887.430 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    PORT
      LAYER met2 ;
        RECT 1903.430 -4.800 1903.990 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    PORT
      LAYER met2 ;
        RECT 1919.990 -4.800 1920.550 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    PORT
      LAYER met2 ;
        RECT 1936.550 -4.800 1937.110 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    PORT
      LAYER met2 ;
        RECT 1969.670 -4.800 1970.230 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    PORT
      LAYER met2 ;
        RECT 1986.230 -4.800 1986.790 2.400 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    PORT
      LAYER met2 ;
        RECT 2002.790 -4.800 2003.350 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    PORT
      LAYER met2 ;
        RECT 810.470 -4.800 811.030 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    PORT
      LAYER met2 ;
        RECT 2019.350 -4.800 2019.910 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    PORT
      LAYER met2 ;
        RECT 2035.910 -4.800 2036.470 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    PORT
      LAYER met2 ;
        RECT 2052.470 -4.800 2053.030 2.400 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    PORT
      LAYER met2 ;
        RECT 2069.030 -4.800 2069.590 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    PORT
      LAYER met2 ;
        RECT 2085.590 -4.800 2086.150 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    PORT
      LAYER met2 ;
        RECT 2102.150 -4.800 2102.710 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    PORT
      LAYER met2 ;
        RECT 2118.710 -4.800 2119.270 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    PORT
      LAYER met2 ;
        RECT 2135.270 -4.800 2135.830 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    PORT
      LAYER met2 ;
        RECT 2151.830 -4.800 2152.390 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    PORT
      LAYER met2 ;
        RECT 2168.390 -4.800 2168.950 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    PORT
      LAYER met2 ;
        RECT 827.030 -4.800 827.590 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    PORT
      LAYER met2 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    PORT
      LAYER met2 ;
        RECT 2201.510 -4.800 2202.070 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    PORT
      LAYER met2 ;
        RECT 2218.070 -4.800 2218.630 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    PORT
      LAYER met2 ;
        RECT 2234.630 -4.800 2235.190 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    PORT
      LAYER met2 ;
        RECT 2251.190 -4.800 2251.750 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    PORT
      LAYER met2 ;
        RECT 2267.750 -4.800 2268.310 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    PORT
      LAYER met2 ;
        RECT 2284.310 -4.800 2284.870 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    PORT
      LAYER met2 ;
        RECT 2300.870 -4.800 2301.430 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    PORT
      LAYER met2 ;
        RECT 2317.430 -4.800 2317.990 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    PORT
      LAYER met2 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    PORT
      LAYER met2 ;
        RECT 843.590 -4.800 844.150 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    PORT
      LAYER met2 ;
        RECT 2803.190 -4.800 2803.750 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    PORT
      LAYER met2 ;
        RECT 2808.710 -4.800 2809.270 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    PORT
      LAYER met2 ;
        RECT 2814.230 -4.800 2814.790 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    PORT
      LAYER met2 ;
        RECT 2819.750 -4.800 2820.310 2.400 ;
    END
  END user_irq[2]
  PIN vccd1
    PORT
      LAYER met5 ;
        RECT -45.180 3459.160 2964.800 3462.260 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3403.130 2964.800 3406.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3347.100 2964.800 3350.200 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3291.070 2964.800 3294.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3235.040 2964.800 3238.140 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3179.010 2964.800 3182.110 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3122.980 2964.800 3126.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3066.950 2964.800 3070.050 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3010.920 2964.800 3014.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2954.890 2964.800 2957.990 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2898.860 2964.800 2901.960 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2842.830 2964.800 2845.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2786.800 2964.800 2789.900 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2730.770 2964.800 2733.870 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2674.740 2964.800 2677.840 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2618.710 2964.800 2621.810 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2562.680 2964.800 2565.780 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2506.650 2964.800 2509.750 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2450.620 2964.800 2453.720 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2394.590 2964.800 2397.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2338.560 2964.800 2341.660 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2282.530 2964.800 2285.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2226.500 2964.800 2229.600 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2170.470 2964.800 2173.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2114.440 2964.800 2117.540 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2058.410 2964.800 2061.510 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2002.380 2964.800 2005.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1946.350 2964.800 1949.450 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1890.320 2964.800 1893.420 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1834.290 2964.800 1837.390 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1778.260 2964.800 1781.360 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1722.230 2964.800 1725.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1666.200 2964.800 1669.300 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1610.170 2964.800 1613.270 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1554.140 2964.800 1557.240 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1498.110 2964.800 1501.210 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1442.080 2964.800 1445.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1386.050 2964.800 1389.150 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1330.020 2964.800 1333.120 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1273.990 2964.800 1277.090 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1217.960 2964.800 1221.060 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1161.930 2964.800 1165.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1105.900 2964.800 1109.000 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1049.870 2964.800 1052.970 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 993.840 2964.800 996.940 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 937.810 2964.800 940.910 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 881.780 2964.800 884.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 825.750 2964.800 828.850 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 769.720 2964.800 772.820 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 713.690 2964.800 716.790 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 657.660 2964.800 660.760 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 601.630 2964.800 604.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 545.600 2964.800 548.700 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 489.570 2964.800 492.670 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 433.540 2964.800 436.640 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 377.510 2964.800 380.610 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 321.480 2964.800 324.580 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 265.450 2964.800 268.550 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 209.420 2964.800 212.520 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 153.390 2964.800 156.490 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 97.360 2964.800 100.460 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 41.330 2964.800 44.430 ;
    END
    PORT
      LAYER met4 ;
        RECT 2928.100 -6.220 2931.200 3525.900 ;
    END
    PORT
      LAYER met5 ;
        RECT -11.580 3522.800 2931.200 3525.900 ;
    END
    PORT
      LAYER met5 ;
        RECT -11.580 -6.220 2931.200 -3.120 ;
    END
    PORT
      LAYER met4 ;
        RECT -11.580 -6.220 -8.480 3525.900 ;
    END
  END vccd1
  PIN vccd2
    PORT
      LAYER met4 ;
        RECT 2937.700 -15.820 2940.800 3535.500 ;
    END
    PORT
      LAYER met5 ;
        RECT -21.180 3532.400 2940.800 3535.500 ;
    END
    PORT
      LAYER met5 ;
        RECT -21.180 -15.820 2940.800 -12.720 ;
    END
    PORT
      LAYER met4 ;
        RECT -21.180 -15.820 -18.080 3535.500 ;
    END
  END vccd2
  PIN vdda1
    PORT
      LAYER met4 ;
        RECT 2947.300 -25.420 2950.400 3545.100 ;
    END
    PORT
      LAYER met5 ;
        RECT -30.780 3542.000 2950.400 3545.100 ;
    END
    PORT
      LAYER met5 ;
        RECT -30.780 -25.420 2950.400 -22.320 ;
    END
    PORT
      LAYER met4 ;
        RECT -30.780 -25.420 -27.680 3545.100 ;
    END
  END vdda1
  PIN vdda2
    PORT
      LAYER met4 ;
        RECT 2956.900 -35.020 2960.000 3554.700 ;
    END
    PORT
      LAYER met5 ;
        RECT -40.380 3551.600 2960.000 3554.700 ;
    END
    PORT
      LAYER met5 ;
        RECT -40.380 -35.020 2960.000 -31.920 ;
    END
    PORT
      LAYER met4 ;
        RECT -40.380 -35.020 -37.280 3554.700 ;
    END
  END vdda2
  PIN vssa1
    PORT
      LAYER met4 ;
        RECT 2952.100 -30.220 2955.200 3549.900 ;
    END
    PORT
      LAYER met5 ;
        RECT -35.580 3546.800 2955.200 3549.900 ;
    END
    PORT
      LAYER met5 ;
        RECT -35.580 -30.220 2955.200 -27.120 ;
    END
    PORT
      LAYER met4 ;
        RECT -35.580 -30.220 -32.480 3549.900 ;
    END
  END vssa1
  PIN vssa2
    PORT
      LAYER met4 ;
        RECT 2961.700 -39.820 2964.800 3559.500 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3556.400 2964.800 3559.500 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 -39.820 2964.800 -36.720 ;
    END
    PORT
      LAYER met4 ;
        RECT -45.180 -39.820 -42.080 3559.500 ;
    END
  END vssa2
  PIN vssd1
    PORT
      LAYER met5 ;
        RECT -45.180 3477.760 2964.800 3480.860 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3421.730 2964.800 3424.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3365.700 2964.800 3368.800 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3309.670 2964.800 3312.770 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3253.640 2964.800 3256.740 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3197.610 2964.800 3200.710 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3141.580 2964.800 3144.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3085.550 2964.800 3088.650 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3029.520 2964.800 3032.620 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2973.490 2964.800 2976.590 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2917.460 2964.800 2920.560 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2861.430 2964.800 2864.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2805.400 2964.800 2808.500 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2749.370 2964.800 2752.470 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2693.340 2964.800 2696.440 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2637.310 2964.800 2640.410 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2581.280 2964.800 2584.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2525.250 2964.800 2528.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2469.220 2964.800 2472.320 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2413.190 2964.800 2416.290 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2357.160 2964.800 2360.260 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2301.130 2964.800 2304.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2245.100 2964.800 2248.200 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2189.070 2964.800 2192.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2133.040 2964.800 2136.140 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2077.010 2964.800 2080.110 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2020.980 2964.800 2024.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1964.950 2964.800 1968.050 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1908.920 2964.800 1912.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1852.890 2964.800 1855.990 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1796.860 2964.800 1799.960 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1740.830 2964.800 1743.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1684.800 2964.800 1687.900 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1628.770 2964.800 1631.870 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1572.740 2964.800 1575.840 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1516.710 2964.800 1519.810 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1460.680 2964.800 1463.780 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1404.650 2964.800 1407.750 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1348.620 2964.800 1351.720 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1292.590 2964.800 1295.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1236.560 2964.800 1239.660 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1180.530 2964.800 1183.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1124.500 2964.800 1127.600 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1068.470 2964.800 1071.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1012.440 2964.800 1015.540 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 956.410 2964.800 959.510 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 900.380 2964.800 903.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 844.350 2964.800 847.450 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 788.320 2964.800 791.420 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 732.290 2964.800 735.390 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 676.260 2964.800 679.360 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 620.230 2964.800 623.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 564.200 2964.800 567.300 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 508.170 2964.800 511.270 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 452.140 2964.800 455.240 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 396.110 2964.800 399.210 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 340.080 2964.800 343.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 284.050 2964.800 287.150 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 228.020 2964.800 231.120 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 171.990 2964.800 175.090 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 115.960 2964.800 119.060 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 59.930 2964.800 63.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 2932.900 -11.020 2936.000 3530.700 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3527.600 2936.000 3530.700 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 -11.020 2936.000 -7.920 ;
    END
    PORT
      LAYER met4 ;
        RECT -16.380 -11.020 -13.280 3530.700 ;
    END
  END vssd1
  PIN vssd2
    PORT
      LAYER met4 ;
        RECT 2942.500 -20.620 2945.600 3540.300 ;
    END
    PORT
      LAYER met5 ;
        RECT -25.980 3537.200 2945.600 3540.300 ;
    END
    PORT
      LAYER met5 ;
        RECT -25.980 -20.620 2945.600 -17.520 ;
    END
    PORT
      LAYER met4 ;
        RECT -25.980 -20.620 -22.880 3540.300 ;
    END
  END vssd2
  PIN wb_clk_i
    PORT
      LAYER met2 ;
        RECT 98.390 -4.800 98.950 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    PORT
      LAYER met2 ;
        RECT 103.910 -4.800 104.470 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    PORT
      LAYER met2 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    PORT
      LAYER met2 ;
        RECT 131.510 -4.800 132.070 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    PORT
      LAYER met2 ;
        RECT 319.190 -4.800 319.750 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    PORT
      LAYER met2 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    PORT
      LAYER met2 ;
        RECT 352.310 -4.800 352.870 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    PORT
      LAYER met2 ;
        RECT 368.870 -4.800 369.430 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    PORT
      LAYER met2 ;
        RECT 385.430 -4.800 385.990 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    PORT
      LAYER met2 ;
        RECT 401.990 -4.800 402.550 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    PORT
      LAYER met2 ;
        RECT 418.550 -4.800 419.110 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    PORT
      LAYER met2 ;
        RECT 435.110 -4.800 435.670 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    PORT
      LAYER met2 ;
        RECT 451.670 -4.800 452.230 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    PORT
      LAYER met2 ;
        RECT 468.230 -4.800 468.790 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    PORT
      LAYER met2 ;
        RECT 153.590 -4.800 154.150 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    PORT
      LAYER met2 ;
        RECT 484.790 -4.800 485.350 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    PORT
      LAYER met2 ;
        RECT 501.350 -4.800 501.910 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    PORT
      LAYER met2 ;
        RECT 517.910 -4.800 518.470 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    PORT
      LAYER met2 ;
        RECT 534.470 -4.800 535.030 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    PORT
      LAYER met2 ;
        RECT 551.030 -4.800 551.590 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    PORT
      LAYER met2 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    PORT
      LAYER met2 ;
        RECT 584.150 -4.800 584.710 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    PORT
      LAYER met2 ;
        RECT 600.710 -4.800 601.270 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    PORT
      LAYER met2 ;
        RECT 617.270 -4.800 617.830 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    PORT
      LAYER met2 ;
        RECT 633.830 -4.800 634.390 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    PORT
      LAYER met2 ;
        RECT 175.670 -4.800 176.230 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    PORT
      LAYER met2 ;
        RECT 650.390 -4.800 650.950 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    PORT
      LAYER met2 ;
        RECT 666.950 -4.800 667.510 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    PORT
      LAYER met2 ;
        RECT 197.750 -4.800 198.310 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    PORT
      LAYER met2 ;
        RECT 219.830 -4.800 220.390 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    PORT
      LAYER met2 ;
        RECT 236.390 -4.800 236.950 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    PORT
      LAYER met2 ;
        RECT 252.950 -4.800 253.510 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    PORT
      LAYER met2 ;
        RECT 269.510 -4.800 270.070 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    PORT
      LAYER met2 ;
        RECT 286.070 -4.800 286.630 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    PORT
      LAYER met2 ;
        RECT 302.630 -4.800 303.190 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    PORT
      LAYER met2 ;
        RECT 114.950 -4.800 115.510 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    PORT
      LAYER met2 ;
        RECT 137.030 -4.800 137.590 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    PORT
      LAYER met2 ;
        RECT 324.710 -4.800 325.270 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    PORT
      LAYER met2 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    PORT
      LAYER met2 ;
        RECT 357.830 -4.800 358.390 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    PORT
      LAYER met2 ;
        RECT 374.390 -4.800 374.950 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    PORT
      LAYER met2 ;
        RECT 390.950 -4.800 391.510 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    PORT
      LAYER met2 ;
        RECT 407.510 -4.800 408.070 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    PORT
      LAYER met2 ;
        RECT 424.070 -4.800 424.630 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    PORT
      LAYER met2 ;
        RECT 440.630 -4.800 441.190 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    PORT
      LAYER met2 ;
        RECT 457.190 -4.800 457.750 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    PORT
      LAYER met2 ;
        RECT 473.750 -4.800 474.310 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    PORT
      LAYER met2 ;
        RECT 159.110 -4.800 159.670 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    PORT
      LAYER met2 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    PORT
      LAYER met2 ;
        RECT 506.870 -4.800 507.430 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    PORT
      LAYER met2 ;
        RECT 523.430 -4.800 523.990 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    PORT
      LAYER met2 ;
        RECT 539.990 -4.800 540.550 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    PORT
      LAYER met2 ;
        RECT 556.550 -4.800 557.110 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    PORT
      LAYER met2 ;
        RECT 573.110 -4.800 573.670 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    PORT
      LAYER met2 ;
        RECT 589.670 -4.800 590.230 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    PORT
      LAYER met2 ;
        RECT 606.230 -4.800 606.790 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    PORT
      LAYER met2 ;
        RECT 622.790 -4.800 623.350 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    PORT
      LAYER met2 ;
        RECT 639.350 -4.800 639.910 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    PORT
      LAYER met2 ;
        RECT 181.190 -4.800 181.750 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    PORT
      LAYER met2 ;
        RECT 655.910 -4.800 656.470 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    PORT
      LAYER met2 ;
        RECT 672.470 -4.800 673.030 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    PORT
      LAYER met2 ;
        RECT 203.270 -4.800 203.830 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    PORT
      LAYER met2 ;
        RECT 225.350 -4.800 225.910 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    PORT
      LAYER met2 ;
        RECT 241.910 -4.800 242.470 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    PORT
      LAYER met2 ;
        RECT 258.470 -4.800 259.030 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    PORT
      LAYER met2 ;
        RECT 275.030 -4.800 275.590 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    PORT
      LAYER met2 ;
        RECT 291.590 -4.800 292.150 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    PORT
      LAYER met2 ;
        RECT 308.150 -4.800 308.710 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    PORT
      LAYER met2 ;
        RECT 142.550 -4.800 143.110 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    PORT
      LAYER met2 ;
        RECT 330.230 -4.800 330.790 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    PORT
      LAYER met2 ;
        RECT 346.790 -4.800 347.350 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    PORT
      LAYER met2 ;
        RECT 363.350 -4.800 363.910 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    PORT
      LAYER met2 ;
        RECT 379.910 -4.800 380.470 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    PORT
      LAYER met2 ;
        RECT 396.470 -4.800 397.030 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    PORT
      LAYER met2 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    PORT
      LAYER met2 ;
        RECT 429.590 -4.800 430.150 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    PORT
      LAYER met2 ;
        RECT 446.150 -4.800 446.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    PORT
      LAYER met2 ;
        RECT 462.710 -4.800 463.270 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    PORT
      LAYER met2 ;
        RECT 479.270 -4.800 479.830 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    PORT
      LAYER met2 ;
        RECT 164.630 -4.800 165.190 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    PORT
      LAYER met2 ;
        RECT 495.830 -4.800 496.390 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    PORT
      LAYER met2 ;
        RECT 512.390 -4.800 512.950 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    PORT
      LAYER met2 ;
        RECT 528.950 -4.800 529.510 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    PORT
      LAYER met2 ;
        RECT 545.510 -4.800 546.070 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    PORT
      LAYER met2 ;
        RECT 562.070 -4.800 562.630 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    PORT
      LAYER met2 ;
        RECT 578.630 -4.800 579.190 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    PORT
      LAYER met2 ;
        RECT 595.190 -4.800 595.750 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    PORT
      LAYER met2 ;
        RECT 611.750 -4.800 612.310 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    PORT
      LAYER met2 ;
        RECT 628.310 -4.800 628.870 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    PORT
      LAYER met2 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    PORT
      LAYER met2 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    PORT
      LAYER met2 ;
        RECT 661.430 -4.800 661.990 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    PORT
      LAYER met2 ;
        RECT 677.990 -4.800 678.550 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    PORT
      LAYER met2 ;
        RECT 208.790 -4.800 209.350 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    PORT
      LAYER met2 ;
        RECT 230.870 -4.800 231.430 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    PORT
      LAYER met2 ;
        RECT 247.430 -4.800 247.990 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    PORT
      LAYER met2 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    PORT
      LAYER met2 ;
        RECT 280.550 -4.800 281.110 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    PORT
      LAYER met2 ;
        RECT 297.110 -4.800 297.670 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    PORT
      LAYER met2 ;
        RECT 313.670 -4.800 314.230 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    PORT
      LAYER met2 ;
        RECT 148.070 -4.800 148.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    PORT
      LAYER met2 ;
        RECT 170.150 -4.800 170.710 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    PORT
      LAYER met2 ;
        RECT 192.230 -4.800 192.790 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    PORT
      LAYER met2 ;
        RECT 214.310 -4.800 214.870 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    PORT
      LAYER met2 ;
        RECT 120.470 -4.800 121.030 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    PORT
      LAYER met2 ;
        RECT 125.990 -4.800 126.550 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 4.560 83.035 2915.440 3436.965 ;
      LAYER met1 ;
        RECT 0.530 1.060 2918.170 3505.020 ;
      LAYER met2 ;
        RECT 0.550 3517.320 41.990 3517.600 ;
        RECT 43.110 3517.320 122.950 3517.600 ;
        RECT 124.070 3517.320 203.910 3517.600 ;
        RECT 205.030 3517.320 284.870 3517.600 ;
        RECT 285.990 3517.320 365.830 3517.600 ;
        RECT 366.950 3517.320 446.790 3517.600 ;
        RECT 447.910 3517.320 527.750 3517.600 ;
        RECT 528.870 3517.320 608.710 3517.600 ;
        RECT 609.830 3517.320 689.670 3517.600 ;
        RECT 690.790 3517.320 770.630 3517.600 ;
        RECT 771.750 3517.320 851.590 3517.600 ;
        RECT 852.710 3517.320 932.550 3517.600 ;
        RECT 933.670 3517.320 1013.510 3517.600 ;
        RECT 1014.630 3517.320 1094.470 3517.600 ;
        RECT 1095.590 3517.320 1175.430 3517.600 ;
        RECT 1176.550 3517.320 1256.390 3517.600 ;
        RECT 1257.510 3517.320 1337.350 3517.600 ;
        RECT 1338.470 3517.320 1418.310 3517.600 ;
        RECT 1419.430 3517.320 1499.270 3517.600 ;
        RECT 1500.390 3517.320 1580.230 3517.600 ;
        RECT 1581.350 3517.320 1661.190 3517.600 ;
        RECT 1662.310 3517.320 1742.150 3517.600 ;
        RECT 1743.270 3517.320 1823.110 3517.600 ;
        RECT 1824.230 3517.320 1904.070 3517.600 ;
        RECT 1905.190 3517.320 1985.030 3517.600 ;
        RECT 1986.150 3517.320 2065.990 3517.600 ;
        RECT 2067.110 3517.320 2146.950 3517.600 ;
        RECT 2148.070 3517.320 2227.910 3517.600 ;
        RECT 2229.030 3517.320 2308.870 3517.600 ;
        RECT 2309.990 3517.320 2389.830 3517.600 ;
        RECT 2390.950 3517.320 2470.790 3517.600 ;
        RECT 2471.910 3517.320 2551.750 3517.600 ;
        RECT 2552.870 3517.320 2632.710 3517.600 ;
        RECT 2633.830 3517.320 2713.670 3517.600 ;
        RECT 2714.790 3517.320 2794.630 3517.600 ;
        RECT 2795.750 3517.320 2875.590 3517.600 ;
        RECT 2876.710 3517.320 2918.150 3517.600 ;
        RECT 0.550 2.680 2918.150 3517.320 ;
        RECT 0.550 0.950 98.110 2.680 ;
        RECT 99.230 0.950 103.630 2.680 ;
        RECT 104.750 0.950 109.150 2.680 ;
        RECT 110.270 0.950 114.670 2.680 ;
        RECT 115.790 0.950 120.190 2.680 ;
        RECT 121.310 0.950 125.710 2.680 ;
        RECT 126.830 0.950 131.230 2.680 ;
        RECT 132.350 0.950 136.750 2.680 ;
        RECT 137.870 0.950 142.270 2.680 ;
        RECT 143.390 0.950 147.790 2.680 ;
        RECT 148.910 0.950 153.310 2.680 ;
        RECT 154.430 0.950 158.830 2.680 ;
        RECT 159.950 0.950 164.350 2.680 ;
        RECT 165.470 0.950 169.870 2.680 ;
        RECT 170.990 0.950 175.390 2.680 ;
        RECT 176.510 0.950 180.910 2.680 ;
        RECT 182.030 0.950 186.430 2.680 ;
        RECT 187.550 0.950 191.950 2.680 ;
        RECT 193.070 0.950 197.470 2.680 ;
        RECT 198.590 0.950 202.990 2.680 ;
        RECT 204.110 0.950 208.510 2.680 ;
        RECT 209.630 0.950 214.030 2.680 ;
        RECT 215.150 0.950 219.550 2.680 ;
        RECT 220.670 0.950 225.070 2.680 ;
        RECT 226.190 0.950 230.590 2.680 ;
        RECT 231.710 0.950 236.110 2.680 ;
        RECT 237.230 0.950 241.630 2.680 ;
        RECT 242.750 0.950 247.150 2.680 ;
        RECT 248.270 0.950 252.670 2.680 ;
        RECT 253.790 0.950 258.190 2.680 ;
        RECT 259.310 0.950 263.710 2.680 ;
        RECT 264.830 0.950 269.230 2.680 ;
        RECT 270.350 0.950 274.750 2.680 ;
        RECT 275.870 0.950 280.270 2.680 ;
        RECT 281.390 0.950 285.790 2.680 ;
        RECT 286.910 0.950 291.310 2.680 ;
        RECT 292.430 0.950 296.830 2.680 ;
        RECT 297.950 0.950 302.350 2.680 ;
        RECT 303.470 0.950 307.870 2.680 ;
        RECT 308.990 0.950 313.390 2.680 ;
        RECT 314.510 0.950 318.910 2.680 ;
        RECT 320.030 0.950 324.430 2.680 ;
        RECT 325.550 0.950 329.950 2.680 ;
        RECT 331.070 0.950 335.470 2.680 ;
        RECT 336.590 0.950 340.990 2.680 ;
        RECT 342.110 0.950 346.510 2.680 ;
        RECT 347.630 0.950 352.030 2.680 ;
        RECT 353.150 0.950 357.550 2.680 ;
        RECT 358.670 0.950 363.070 2.680 ;
        RECT 364.190 0.950 368.590 2.680 ;
        RECT 369.710 0.950 374.110 2.680 ;
        RECT 375.230 0.950 379.630 2.680 ;
        RECT 380.750 0.950 385.150 2.680 ;
        RECT 386.270 0.950 390.670 2.680 ;
        RECT 391.790 0.950 396.190 2.680 ;
        RECT 397.310 0.950 401.710 2.680 ;
        RECT 402.830 0.950 407.230 2.680 ;
        RECT 408.350 0.950 412.750 2.680 ;
        RECT 413.870 0.950 418.270 2.680 ;
        RECT 419.390 0.950 423.790 2.680 ;
        RECT 424.910 0.950 429.310 2.680 ;
        RECT 430.430 0.950 434.830 2.680 ;
        RECT 435.950 0.950 440.350 2.680 ;
        RECT 441.470 0.950 445.870 2.680 ;
        RECT 446.990 0.950 451.390 2.680 ;
        RECT 452.510 0.950 456.910 2.680 ;
        RECT 458.030 0.950 462.430 2.680 ;
        RECT 463.550 0.950 467.950 2.680 ;
        RECT 469.070 0.950 473.470 2.680 ;
        RECT 474.590 0.950 478.990 2.680 ;
        RECT 480.110 0.950 484.510 2.680 ;
        RECT 485.630 0.950 490.030 2.680 ;
        RECT 491.150 0.950 495.550 2.680 ;
        RECT 496.670 0.950 501.070 2.680 ;
        RECT 502.190 0.950 506.590 2.680 ;
        RECT 507.710 0.950 512.110 2.680 ;
        RECT 513.230 0.950 517.630 2.680 ;
        RECT 518.750 0.950 523.150 2.680 ;
        RECT 524.270 0.950 528.670 2.680 ;
        RECT 529.790 0.950 534.190 2.680 ;
        RECT 535.310 0.950 539.710 2.680 ;
        RECT 540.830 0.950 545.230 2.680 ;
        RECT 546.350 0.950 550.750 2.680 ;
        RECT 551.870 0.950 556.270 2.680 ;
        RECT 557.390 0.950 561.790 2.680 ;
        RECT 562.910 0.950 567.310 2.680 ;
        RECT 568.430 0.950 572.830 2.680 ;
        RECT 573.950 0.950 578.350 2.680 ;
        RECT 579.470 0.950 583.870 2.680 ;
        RECT 584.990 0.950 589.390 2.680 ;
        RECT 590.510 0.950 594.910 2.680 ;
        RECT 596.030 0.950 600.430 2.680 ;
        RECT 601.550 0.950 605.950 2.680 ;
        RECT 607.070 0.950 611.470 2.680 ;
        RECT 612.590 0.950 616.990 2.680 ;
        RECT 618.110 0.950 622.510 2.680 ;
        RECT 623.630 0.950 628.030 2.680 ;
        RECT 629.150 0.950 633.550 2.680 ;
        RECT 634.670 0.950 639.070 2.680 ;
        RECT 640.190 0.950 644.590 2.680 ;
        RECT 645.710 0.950 650.110 2.680 ;
        RECT 651.230 0.950 655.630 2.680 ;
        RECT 656.750 0.950 661.150 2.680 ;
        RECT 662.270 0.950 666.670 2.680 ;
        RECT 667.790 0.950 672.190 2.680 ;
        RECT 673.310 0.950 677.710 2.680 ;
        RECT 678.830 0.950 683.230 2.680 ;
        RECT 684.350 0.950 688.750 2.680 ;
        RECT 689.870 0.950 694.270 2.680 ;
        RECT 695.390 0.950 699.790 2.680 ;
        RECT 700.910 0.950 705.310 2.680 ;
        RECT 706.430 0.950 710.830 2.680 ;
        RECT 711.950 0.950 716.350 2.680 ;
        RECT 717.470 0.950 721.870 2.680 ;
        RECT 722.990 0.950 727.390 2.680 ;
        RECT 728.510 0.950 732.910 2.680 ;
        RECT 734.030 0.950 738.430 2.680 ;
        RECT 739.550 0.950 743.950 2.680 ;
        RECT 745.070 0.950 749.470 2.680 ;
        RECT 750.590 0.950 754.990 2.680 ;
        RECT 756.110 0.950 760.510 2.680 ;
        RECT 761.630 0.950 766.030 2.680 ;
        RECT 767.150 0.950 771.550 2.680 ;
        RECT 772.670 0.950 777.070 2.680 ;
        RECT 778.190 0.950 782.590 2.680 ;
        RECT 783.710 0.950 788.110 2.680 ;
        RECT 789.230 0.950 793.630 2.680 ;
        RECT 794.750 0.950 799.150 2.680 ;
        RECT 800.270 0.950 804.670 2.680 ;
        RECT 805.790 0.950 810.190 2.680 ;
        RECT 811.310 0.950 815.710 2.680 ;
        RECT 816.830 0.950 821.230 2.680 ;
        RECT 822.350 0.950 826.750 2.680 ;
        RECT 827.870 0.950 832.270 2.680 ;
        RECT 833.390 0.950 837.790 2.680 ;
        RECT 838.910 0.950 843.310 2.680 ;
        RECT 844.430 0.950 848.830 2.680 ;
        RECT 849.950 0.950 854.350 2.680 ;
        RECT 855.470 0.950 859.870 2.680 ;
        RECT 860.990 0.950 865.390 2.680 ;
        RECT 866.510 0.950 870.910 2.680 ;
        RECT 872.030 0.950 876.430 2.680 ;
        RECT 877.550 0.950 881.950 2.680 ;
        RECT 883.070 0.950 887.470 2.680 ;
        RECT 888.590 0.950 892.990 2.680 ;
        RECT 894.110 0.950 898.510 2.680 ;
        RECT 899.630 0.950 904.030 2.680 ;
        RECT 905.150 0.950 909.550 2.680 ;
        RECT 910.670 0.950 915.070 2.680 ;
        RECT 916.190 0.950 920.590 2.680 ;
        RECT 921.710 0.950 926.110 2.680 ;
        RECT 927.230 0.950 931.630 2.680 ;
        RECT 932.750 0.950 937.150 2.680 ;
        RECT 938.270 0.950 942.670 2.680 ;
        RECT 943.790 0.950 948.190 2.680 ;
        RECT 949.310 0.950 953.710 2.680 ;
        RECT 954.830 0.950 959.230 2.680 ;
        RECT 960.350 0.950 964.750 2.680 ;
        RECT 965.870 0.950 970.270 2.680 ;
        RECT 971.390 0.950 975.790 2.680 ;
        RECT 976.910 0.950 981.310 2.680 ;
        RECT 982.430 0.950 986.830 2.680 ;
        RECT 987.950 0.950 992.350 2.680 ;
        RECT 993.470 0.950 997.870 2.680 ;
        RECT 998.990 0.950 1003.390 2.680 ;
        RECT 1004.510 0.950 1008.910 2.680 ;
        RECT 1010.030 0.950 1014.430 2.680 ;
        RECT 1015.550 0.950 1019.950 2.680 ;
        RECT 1021.070 0.950 1025.470 2.680 ;
        RECT 1026.590 0.950 1030.990 2.680 ;
        RECT 1032.110 0.950 1036.510 2.680 ;
        RECT 1037.630 0.950 1042.030 2.680 ;
        RECT 1043.150 0.950 1047.550 2.680 ;
        RECT 1048.670 0.950 1053.070 2.680 ;
        RECT 1054.190 0.950 1058.590 2.680 ;
        RECT 1059.710 0.950 1064.110 2.680 ;
        RECT 1065.230 0.950 1069.630 2.680 ;
        RECT 1070.750 0.950 1075.150 2.680 ;
        RECT 1076.270 0.950 1080.670 2.680 ;
        RECT 1081.790 0.950 1086.190 2.680 ;
        RECT 1087.310 0.950 1091.710 2.680 ;
        RECT 1092.830 0.950 1097.230 2.680 ;
        RECT 1098.350 0.950 1102.750 2.680 ;
        RECT 1103.870 0.950 1108.270 2.680 ;
        RECT 1109.390 0.950 1113.790 2.680 ;
        RECT 1114.910 0.950 1119.310 2.680 ;
        RECT 1120.430 0.950 1124.830 2.680 ;
        RECT 1125.950 0.950 1130.350 2.680 ;
        RECT 1131.470 0.950 1135.870 2.680 ;
        RECT 1136.990 0.950 1141.390 2.680 ;
        RECT 1142.510 0.950 1146.910 2.680 ;
        RECT 1148.030 0.950 1152.430 2.680 ;
        RECT 1153.550 0.950 1157.950 2.680 ;
        RECT 1159.070 0.950 1163.470 2.680 ;
        RECT 1164.590 0.950 1168.990 2.680 ;
        RECT 1170.110 0.950 1174.510 2.680 ;
        RECT 1175.630 0.950 1180.030 2.680 ;
        RECT 1181.150 0.950 1185.550 2.680 ;
        RECT 1186.670 0.950 1191.070 2.680 ;
        RECT 1192.190 0.950 1196.590 2.680 ;
        RECT 1197.710 0.950 1202.110 2.680 ;
        RECT 1203.230 0.950 1207.630 2.680 ;
        RECT 1208.750 0.950 1213.150 2.680 ;
        RECT 1214.270 0.950 1218.670 2.680 ;
        RECT 1219.790 0.950 1224.190 2.680 ;
        RECT 1225.310 0.950 1229.710 2.680 ;
        RECT 1230.830 0.950 1235.230 2.680 ;
        RECT 1236.350 0.950 1240.750 2.680 ;
        RECT 1241.870 0.950 1246.270 2.680 ;
        RECT 1247.390 0.950 1251.790 2.680 ;
        RECT 1252.910 0.950 1257.310 2.680 ;
        RECT 1258.430 0.950 1262.830 2.680 ;
        RECT 1263.950 0.950 1268.350 2.680 ;
        RECT 1269.470 0.950 1273.870 2.680 ;
        RECT 1274.990 0.950 1279.390 2.680 ;
        RECT 1280.510 0.950 1284.910 2.680 ;
        RECT 1286.030 0.950 1290.430 2.680 ;
        RECT 1291.550 0.950 1295.950 2.680 ;
        RECT 1297.070 0.950 1301.470 2.680 ;
        RECT 1302.590 0.950 1306.990 2.680 ;
        RECT 1308.110 0.950 1312.510 2.680 ;
        RECT 1313.630 0.950 1318.030 2.680 ;
        RECT 1319.150 0.950 1323.550 2.680 ;
        RECT 1324.670 0.950 1329.070 2.680 ;
        RECT 1330.190 0.950 1334.590 2.680 ;
        RECT 1335.710 0.950 1340.110 2.680 ;
        RECT 1341.230 0.950 1345.630 2.680 ;
        RECT 1346.750 0.950 1351.150 2.680 ;
        RECT 1352.270 0.950 1356.670 2.680 ;
        RECT 1357.790 0.950 1362.190 2.680 ;
        RECT 1363.310 0.950 1367.710 2.680 ;
        RECT 1368.830 0.950 1373.230 2.680 ;
        RECT 1374.350 0.950 1378.750 2.680 ;
        RECT 1379.870 0.950 1384.270 2.680 ;
        RECT 1385.390 0.950 1389.790 2.680 ;
        RECT 1390.910 0.950 1395.310 2.680 ;
        RECT 1396.430 0.950 1400.830 2.680 ;
        RECT 1401.950 0.950 1406.350 2.680 ;
        RECT 1407.470 0.950 1411.870 2.680 ;
        RECT 1412.990 0.950 1417.390 2.680 ;
        RECT 1418.510 0.950 1422.910 2.680 ;
        RECT 1424.030 0.950 1428.430 2.680 ;
        RECT 1429.550 0.950 1433.950 2.680 ;
        RECT 1435.070 0.950 1439.470 2.680 ;
        RECT 1440.590 0.950 1444.990 2.680 ;
        RECT 1446.110 0.950 1450.510 2.680 ;
        RECT 1451.630 0.950 1456.030 2.680 ;
        RECT 1457.150 0.950 1461.550 2.680 ;
        RECT 1462.670 0.950 1467.070 2.680 ;
        RECT 1468.190 0.950 1472.590 2.680 ;
        RECT 1473.710 0.950 1478.110 2.680 ;
        RECT 1479.230 0.950 1483.630 2.680 ;
        RECT 1484.750 0.950 1489.150 2.680 ;
        RECT 1490.270 0.950 1494.670 2.680 ;
        RECT 1495.790 0.950 1500.190 2.680 ;
        RECT 1501.310 0.950 1505.710 2.680 ;
        RECT 1506.830 0.950 1511.230 2.680 ;
        RECT 1512.350 0.950 1516.750 2.680 ;
        RECT 1517.870 0.950 1522.270 2.680 ;
        RECT 1523.390 0.950 1527.790 2.680 ;
        RECT 1528.910 0.950 1533.310 2.680 ;
        RECT 1534.430 0.950 1538.830 2.680 ;
        RECT 1539.950 0.950 1544.350 2.680 ;
        RECT 1545.470 0.950 1549.870 2.680 ;
        RECT 1550.990 0.950 1555.390 2.680 ;
        RECT 1556.510 0.950 1560.910 2.680 ;
        RECT 1562.030 0.950 1566.430 2.680 ;
        RECT 1567.550 0.950 1571.950 2.680 ;
        RECT 1573.070 0.950 1577.470 2.680 ;
        RECT 1578.590 0.950 1582.990 2.680 ;
        RECT 1584.110 0.950 1588.510 2.680 ;
        RECT 1589.630 0.950 1594.030 2.680 ;
        RECT 1595.150 0.950 1599.550 2.680 ;
        RECT 1600.670 0.950 1605.070 2.680 ;
        RECT 1606.190 0.950 1610.590 2.680 ;
        RECT 1611.710 0.950 1616.110 2.680 ;
        RECT 1617.230 0.950 1621.630 2.680 ;
        RECT 1622.750 0.950 1627.150 2.680 ;
        RECT 1628.270 0.950 1632.670 2.680 ;
        RECT 1633.790 0.950 1638.190 2.680 ;
        RECT 1639.310 0.950 1643.710 2.680 ;
        RECT 1644.830 0.950 1649.230 2.680 ;
        RECT 1650.350 0.950 1654.750 2.680 ;
        RECT 1655.870 0.950 1660.270 2.680 ;
        RECT 1661.390 0.950 1665.790 2.680 ;
        RECT 1666.910 0.950 1671.310 2.680 ;
        RECT 1672.430 0.950 1676.830 2.680 ;
        RECT 1677.950 0.950 1682.350 2.680 ;
        RECT 1683.470 0.950 1687.870 2.680 ;
        RECT 1688.990 0.950 1693.390 2.680 ;
        RECT 1694.510 0.950 1698.910 2.680 ;
        RECT 1700.030 0.950 1704.430 2.680 ;
        RECT 1705.550 0.950 1709.950 2.680 ;
        RECT 1711.070 0.950 1715.470 2.680 ;
        RECT 1716.590 0.950 1720.990 2.680 ;
        RECT 1722.110 0.950 1726.510 2.680 ;
        RECT 1727.630 0.950 1732.030 2.680 ;
        RECT 1733.150 0.950 1737.550 2.680 ;
        RECT 1738.670 0.950 1743.070 2.680 ;
        RECT 1744.190 0.950 1748.590 2.680 ;
        RECT 1749.710 0.950 1754.110 2.680 ;
        RECT 1755.230 0.950 1759.630 2.680 ;
        RECT 1760.750 0.950 1765.150 2.680 ;
        RECT 1766.270 0.950 1770.670 2.680 ;
        RECT 1771.790 0.950 1776.190 2.680 ;
        RECT 1777.310 0.950 1781.710 2.680 ;
        RECT 1782.830 0.950 1787.230 2.680 ;
        RECT 1788.350 0.950 1792.750 2.680 ;
        RECT 1793.870 0.950 1798.270 2.680 ;
        RECT 1799.390 0.950 1803.790 2.680 ;
        RECT 1804.910 0.950 1809.310 2.680 ;
        RECT 1810.430 0.950 1814.830 2.680 ;
        RECT 1815.950 0.950 1820.350 2.680 ;
        RECT 1821.470 0.950 1825.870 2.680 ;
        RECT 1826.990 0.950 1831.390 2.680 ;
        RECT 1832.510 0.950 1836.910 2.680 ;
        RECT 1838.030 0.950 1842.430 2.680 ;
        RECT 1843.550 0.950 1847.950 2.680 ;
        RECT 1849.070 0.950 1853.470 2.680 ;
        RECT 1854.590 0.950 1858.990 2.680 ;
        RECT 1860.110 0.950 1864.510 2.680 ;
        RECT 1865.630 0.950 1870.030 2.680 ;
        RECT 1871.150 0.950 1875.550 2.680 ;
        RECT 1876.670 0.950 1881.070 2.680 ;
        RECT 1882.190 0.950 1886.590 2.680 ;
        RECT 1887.710 0.950 1892.110 2.680 ;
        RECT 1893.230 0.950 1897.630 2.680 ;
        RECT 1898.750 0.950 1903.150 2.680 ;
        RECT 1904.270 0.950 1908.670 2.680 ;
        RECT 1909.790 0.950 1914.190 2.680 ;
        RECT 1915.310 0.950 1919.710 2.680 ;
        RECT 1920.830 0.950 1925.230 2.680 ;
        RECT 1926.350 0.950 1930.750 2.680 ;
        RECT 1931.870 0.950 1936.270 2.680 ;
        RECT 1937.390 0.950 1941.790 2.680 ;
        RECT 1942.910 0.950 1947.310 2.680 ;
        RECT 1948.430 0.950 1952.830 2.680 ;
        RECT 1953.950 0.950 1958.350 2.680 ;
        RECT 1959.470 0.950 1963.870 2.680 ;
        RECT 1964.990 0.950 1969.390 2.680 ;
        RECT 1970.510 0.950 1974.910 2.680 ;
        RECT 1976.030 0.950 1980.430 2.680 ;
        RECT 1981.550 0.950 1985.950 2.680 ;
        RECT 1987.070 0.950 1991.470 2.680 ;
        RECT 1992.590 0.950 1996.990 2.680 ;
        RECT 1998.110 0.950 2002.510 2.680 ;
        RECT 2003.630 0.950 2008.030 2.680 ;
        RECT 2009.150 0.950 2013.550 2.680 ;
        RECT 2014.670 0.950 2019.070 2.680 ;
        RECT 2020.190 0.950 2024.590 2.680 ;
        RECT 2025.710 0.950 2030.110 2.680 ;
        RECT 2031.230 0.950 2035.630 2.680 ;
        RECT 2036.750 0.950 2041.150 2.680 ;
        RECT 2042.270 0.950 2046.670 2.680 ;
        RECT 2047.790 0.950 2052.190 2.680 ;
        RECT 2053.310 0.950 2057.710 2.680 ;
        RECT 2058.830 0.950 2063.230 2.680 ;
        RECT 2064.350 0.950 2068.750 2.680 ;
        RECT 2069.870 0.950 2074.270 2.680 ;
        RECT 2075.390 0.950 2079.790 2.680 ;
        RECT 2080.910 0.950 2085.310 2.680 ;
        RECT 2086.430 0.950 2090.830 2.680 ;
        RECT 2091.950 0.950 2096.350 2.680 ;
        RECT 2097.470 0.950 2101.870 2.680 ;
        RECT 2102.990 0.950 2107.390 2.680 ;
        RECT 2108.510 0.950 2112.910 2.680 ;
        RECT 2114.030 0.950 2118.430 2.680 ;
        RECT 2119.550 0.950 2123.950 2.680 ;
        RECT 2125.070 0.950 2129.470 2.680 ;
        RECT 2130.590 0.950 2134.990 2.680 ;
        RECT 2136.110 0.950 2140.510 2.680 ;
        RECT 2141.630 0.950 2146.030 2.680 ;
        RECT 2147.150 0.950 2151.550 2.680 ;
        RECT 2152.670 0.950 2157.070 2.680 ;
        RECT 2158.190 0.950 2162.590 2.680 ;
        RECT 2163.710 0.950 2168.110 2.680 ;
        RECT 2169.230 0.950 2173.630 2.680 ;
        RECT 2174.750 0.950 2179.150 2.680 ;
        RECT 2180.270 0.950 2184.670 2.680 ;
        RECT 2185.790 0.950 2190.190 2.680 ;
        RECT 2191.310 0.950 2195.710 2.680 ;
        RECT 2196.830 0.950 2201.230 2.680 ;
        RECT 2202.350 0.950 2206.750 2.680 ;
        RECT 2207.870 0.950 2212.270 2.680 ;
        RECT 2213.390 0.950 2217.790 2.680 ;
        RECT 2218.910 0.950 2223.310 2.680 ;
        RECT 2224.430 0.950 2228.830 2.680 ;
        RECT 2229.950 0.950 2234.350 2.680 ;
        RECT 2235.470 0.950 2239.870 2.680 ;
        RECT 2240.990 0.950 2245.390 2.680 ;
        RECT 2246.510 0.950 2250.910 2.680 ;
        RECT 2252.030 0.950 2256.430 2.680 ;
        RECT 2257.550 0.950 2261.950 2.680 ;
        RECT 2263.070 0.950 2267.470 2.680 ;
        RECT 2268.590 0.950 2272.990 2.680 ;
        RECT 2274.110 0.950 2278.510 2.680 ;
        RECT 2279.630 0.950 2284.030 2.680 ;
        RECT 2285.150 0.950 2289.550 2.680 ;
        RECT 2290.670 0.950 2295.070 2.680 ;
        RECT 2296.190 0.950 2300.590 2.680 ;
        RECT 2301.710 0.950 2306.110 2.680 ;
        RECT 2307.230 0.950 2311.630 2.680 ;
        RECT 2312.750 0.950 2317.150 2.680 ;
        RECT 2318.270 0.950 2322.670 2.680 ;
        RECT 2323.790 0.950 2328.190 2.680 ;
        RECT 2329.310 0.950 2333.710 2.680 ;
        RECT 2334.830 0.950 2339.230 2.680 ;
        RECT 2340.350 0.950 2344.750 2.680 ;
        RECT 2345.870 0.950 2350.270 2.680 ;
        RECT 2351.390 0.950 2355.790 2.680 ;
        RECT 2356.910 0.950 2361.310 2.680 ;
        RECT 2362.430 0.950 2366.830 2.680 ;
        RECT 2367.950 0.950 2372.350 2.680 ;
        RECT 2373.470 0.950 2377.870 2.680 ;
        RECT 2378.990 0.950 2383.390 2.680 ;
        RECT 2384.510 0.950 2388.910 2.680 ;
        RECT 2390.030 0.950 2394.430 2.680 ;
        RECT 2395.550 0.950 2399.950 2.680 ;
        RECT 2401.070 0.950 2405.470 2.680 ;
        RECT 2406.590 0.950 2410.990 2.680 ;
        RECT 2412.110 0.950 2416.510 2.680 ;
        RECT 2417.630 0.950 2422.030 2.680 ;
        RECT 2423.150 0.950 2427.550 2.680 ;
        RECT 2428.670 0.950 2433.070 2.680 ;
        RECT 2434.190 0.950 2438.590 2.680 ;
        RECT 2439.710 0.950 2444.110 2.680 ;
        RECT 2445.230 0.950 2449.630 2.680 ;
        RECT 2450.750 0.950 2455.150 2.680 ;
        RECT 2456.270 0.950 2460.670 2.680 ;
        RECT 2461.790 0.950 2466.190 2.680 ;
        RECT 2467.310 0.950 2471.710 2.680 ;
        RECT 2472.830 0.950 2477.230 2.680 ;
        RECT 2478.350 0.950 2482.750 2.680 ;
        RECT 2483.870 0.950 2488.270 2.680 ;
        RECT 2489.390 0.950 2493.790 2.680 ;
        RECT 2494.910 0.950 2499.310 2.680 ;
        RECT 2500.430 0.950 2504.830 2.680 ;
        RECT 2505.950 0.950 2510.350 2.680 ;
        RECT 2511.470 0.950 2515.870 2.680 ;
        RECT 2516.990 0.950 2521.390 2.680 ;
        RECT 2522.510 0.950 2526.910 2.680 ;
        RECT 2528.030 0.950 2532.430 2.680 ;
        RECT 2533.550 0.950 2537.950 2.680 ;
        RECT 2539.070 0.950 2543.470 2.680 ;
        RECT 2544.590 0.950 2548.990 2.680 ;
        RECT 2550.110 0.950 2554.510 2.680 ;
        RECT 2555.630 0.950 2560.030 2.680 ;
        RECT 2561.150 0.950 2565.550 2.680 ;
        RECT 2566.670 0.950 2571.070 2.680 ;
        RECT 2572.190 0.950 2576.590 2.680 ;
        RECT 2577.710 0.950 2582.110 2.680 ;
        RECT 2583.230 0.950 2587.630 2.680 ;
        RECT 2588.750 0.950 2593.150 2.680 ;
        RECT 2594.270 0.950 2598.670 2.680 ;
        RECT 2599.790 0.950 2604.190 2.680 ;
        RECT 2605.310 0.950 2609.710 2.680 ;
        RECT 2610.830 0.950 2615.230 2.680 ;
        RECT 2616.350 0.950 2620.750 2.680 ;
        RECT 2621.870 0.950 2626.270 2.680 ;
        RECT 2627.390 0.950 2631.790 2.680 ;
        RECT 2632.910 0.950 2637.310 2.680 ;
        RECT 2638.430 0.950 2642.830 2.680 ;
        RECT 2643.950 0.950 2648.350 2.680 ;
        RECT 2649.470 0.950 2653.870 2.680 ;
        RECT 2654.990 0.950 2659.390 2.680 ;
        RECT 2660.510 0.950 2664.910 2.680 ;
        RECT 2666.030 0.950 2670.430 2.680 ;
        RECT 2671.550 0.950 2675.950 2.680 ;
        RECT 2677.070 0.950 2681.470 2.680 ;
        RECT 2682.590 0.950 2686.990 2.680 ;
        RECT 2688.110 0.950 2692.510 2.680 ;
        RECT 2693.630 0.950 2698.030 2.680 ;
        RECT 2699.150 0.950 2703.550 2.680 ;
        RECT 2704.670 0.950 2709.070 2.680 ;
        RECT 2710.190 0.950 2714.590 2.680 ;
        RECT 2715.710 0.950 2720.110 2.680 ;
        RECT 2721.230 0.950 2725.630 2.680 ;
        RECT 2726.750 0.950 2731.150 2.680 ;
        RECT 2732.270 0.950 2736.670 2.680 ;
        RECT 2737.790 0.950 2742.190 2.680 ;
        RECT 2743.310 0.950 2747.710 2.680 ;
        RECT 2748.830 0.950 2753.230 2.680 ;
        RECT 2754.350 0.950 2758.750 2.680 ;
        RECT 2759.870 0.950 2764.270 2.680 ;
        RECT 2765.390 0.950 2769.790 2.680 ;
        RECT 2770.910 0.950 2775.310 2.680 ;
        RECT 2776.430 0.950 2780.830 2.680 ;
        RECT 2781.950 0.950 2786.350 2.680 ;
        RECT 2787.470 0.950 2791.870 2.680 ;
        RECT 2792.990 0.950 2797.390 2.680 ;
        RECT 2798.510 0.950 2802.910 2.680 ;
        RECT 2804.030 0.950 2808.430 2.680 ;
        RECT 2809.550 0.950 2813.950 2.680 ;
        RECT 2815.070 0.950 2819.470 2.680 ;
        RECT 2820.590 0.950 2918.150 2.680 ;
      LAYER met3 ;
        RECT 0.270 3457.100 2918.175 3501.825 ;
        RECT 0.270 3455.100 2917.200 3457.100 ;
        RECT 0.270 3436.700 2918.175 3455.100 ;
        RECT 2.800 3434.700 2918.175 3436.700 ;
        RECT 0.270 3391.820 2918.175 3434.700 ;
        RECT 0.270 3389.820 2917.200 3391.820 ;
        RECT 0.270 3373.460 2918.175 3389.820 ;
        RECT 2.800 3371.460 2918.175 3373.460 ;
        RECT 0.270 3326.540 2918.175 3371.460 ;
        RECT 0.270 3324.540 2917.200 3326.540 ;
        RECT 0.270 3310.220 2918.175 3324.540 ;
        RECT 2.800 3308.220 2918.175 3310.220 ;
        RECT 0.270 3261.260 2918.175 3308.220 ;
        RECT 0.270 3259.260 2917.200 3261.260 ;
        RECT 0.270 3246.980 2918.175 3259.260 ;
        RECT 2.800 3244.980 2918.175 3246.980 ;
        RECT 0.270 3195.980 2918.175 3244.980 ;
        RECT 0.270 3193.980 2917.200 3195.980 ;
        RECT 0.270 3183.740 2918.175 3193.980 ;
        RECT 2.800 3181.740 2918.175 3183.740 ;
        RECT 0.270 3130.700 2918.175 3181.740 ;
        RECT 0.270 3128.700 2917.200 3130.700 ;
        RECT 0.270 3120.500 2918.175 3128.700 ;
        RECT 2.800 3118.500 2918.175 3120.500 ;
        RECT 0.270 3065.420 2918.175 3118.500 ;
        RECT 0.270 3063.420 2917.200 3065.420 ;
        RECT 0.270 3057.260 2918.175 3063.420 ;
        RECT 2.800 3055.260 2918.175 3057.260 ;
        RECT 0.270 3000.140 2918.175 3055.260 ;
        RECT 0.270 2998.140 2917.200 3000.140 ;
        RECT 0.270 2994.020 2918.175 2998.140 ;
        RECT 2.800 2992.020 2918.175 2994.020 ;
        RECT 0.270 2934.860 2918.175 2992.020 ;
        RECT 0.270 2932.860 2917.200 2934.860 ;
        RECT 0.270 2930.780 2918.175 2932.860 ;
        RECT 2.800 2928.780 2918.175 2930.780 ;
        RECT 0.270 2869.580 2918.175 2928.780 ;
        RECT 0.270 2867.580 2917.200 2869.580 ;
        RECT 0.270 2867.540 2918.175 2867.580 ;
        RECT 2.800 2865.540 2918.175 2867.540 ;
        RECT 0.270 2804.300 2918.175 2865.540 ;
        RECT 2.800 2802.300 2917.200 2804.300 ;
        RECT 0.270 2741.060 2918.175 2802.300 ;
        RECT 2.800 2739.060 2918.175 2741.060 ;
        RECT 0.270 2739.020 2918.175 2739.060 ;
        RECT 0.270 2737.020 2917.200 2739.020 ;
        RECT 0.270 2677.820 2918.175 2737.020 ;
        RECT 2.800 2675.820 2918.175 2677.820 ;
        RECT 0.270 2673.740 2918.175 2675.820 ;
        RECT 0.270 2671.740 2917.200 2673.740 ;
        RECT 0.270 2614.580 2918.175 2671.740 ;
        RECT 2.800 2612.580 2918.175 2614.580 ;
        RECT 0.270 2608.460 2918.175 2612.580 ;
        RECT 0.270 2606.460 2917.200 2608.460 ;
        RECT 0.270 2551.340 2918.175 2606.460 ;
        RECT 2.800 2549.340 2918.175 2551.340 ;
        RECT 0.270 2543.180 2918.175 2549.340 ;
        RECT 0.270 2541.180 2917.200 2543.180 ;
        RECT 0.270 2488.100 2918.175 2541.180 ;
        RECT 2.800 2486.100 2918.175 2488.100 ;
        RECT 0.270 2477.900 2918.175 2486.100 ;
        RECT 0.270 2475.900 2917.200 2477.900 ;
        RECT 0.270 2424.860 2918.175 2475.900 ;
        RECT 2.800 2422.860 2918.175 2424.860 ;
        RECT 0.270 2412.620 2918.175 2422.860 ;
        RECT 0.270 2410.620 2917.200 2412.620 ;
        RECT 0.270 2361.620 2918.175 2410.620 ;
        RECT 2.800 2359.620 2918.175 2361.620 ;
        RECT 0.270 2347.340 2918.175 2359.620 ;
        RECT 0.270 2345.340 2917.200 2347.340 ;
        RECT 0.270 2298.380 2918.175 2345.340 ;
        RECT 2.800 2296.380 2918.175 2298.380 ;
        RECT 0.270 2282.060 2918.175 2296.380 ;
        RECT 0.270 2280.060 2917.200 2282.060 ;
        RECT 0.270 2235.140 2918.175 2280.060 ;
        RECT 2.800 2233.140 2918.175 2235.140 ;
        RECT 0.270 2216.780 2918.175 2233.140 ;
        RECT 0.270 2214.780 2917.200 2216.780 ;
        RECT 0.270 2171.900 2918.175 2214.780 ;
        RECT 2.800 2169.900 2918.175 2171.900 ;
        RECT 0.270 2151.500 2918.175 2169.900 ;
        RECT 0.270 2149.500 2917.200 2151.500 ;
        RECT 0.270 2108.660 2918.175 2149.500 ;
        RECT 2.800 2106.660 2918.175 2108.660 ;
        RECT 0.270 2086.220 2918.175 2106.660 ;
        RECT 0.270 2084.220 2917.200 2086.220 ;
        RECT 0.270 2045.420 2918.175 2084.220 ;
        RECT 2.800 2043.420 2918.175 2045.420 ;
        RECT 0.270 2020.940 2918.175 2043.420 ;
        RECT 0.270 2018.940 2917.200 2020.940 ;
        RECT 0.270 1982.180 2918.175 2018.940 ;
        RECT 2.800 1980.180 2918.175 1982.180 ;
        RECT 0.270 1955.660 2918.175 1980.180 ;
        RECT 0.270 1953.660 2917.200 1955.660 ;
        RECT 0.270 1918.940 2918.175 1953.660 ;
        RECT 2.800 1916.940 2918.175 1918.940 ;
        RECT 0.270 1890.380 2918.175 1916.940 ;
        RECT 0.270 1888.380 2917.200 1890.380 ;
        RECT 0.270 1855.700 2918.175 1888.380 ;
        RECT 2.800 1853.700 2918.175 1855.700 ;
        RECT 0.270 1825.100 2918.175 1853.700 ;
        RECT 0.270 1823.100 2917.200 1825.100 ;
        RECT 0.270 1792.460 2918.175 1823.100 ;
        RECT 2.800 1790.460 2918.175 1792.460 ;
        RECT 0.270 1759.820 2918.175 1790.460 ;
        RECT 0.270 1757.820 2917.200 1759.820 ;
        RECT 0.270 1729.220 2918.175 1757.820 ;
        RECT 2.800 1727.220 2918.175 1729.220 ;
        RECT 0.270 1694.540 2918.175 1727.220 ;
        RECT 0.270 1692.540 2917.200 1694.540 ;
        RECT 0.270 1665.980 2918.175 1692.540 ;
        RECT 2.800 1663.980 2918.175 1665.980 ;
        RECT 0.270 1629.260 2918.175 1663.980 ;
        RECT 0.270 1627.260 2917.200 1629.260 ;
        RECT 0.270 1602.740 2918.175 1627.260 ;
        RECT 2.800 1600.740 2918.175 1602.740 ;
        RECT 0.270 1563.980 2918.175 1600.740 ;
        RECT 0.270 1561.980 2917.200 1563.980 ;
        RECT 0.270 1539.500 2918.175 1561.980 ;
        RECT 2.800 1537.500 2918.175 1539.500 ;
        RECT 0.270 1498.700 2918.175 1537.500 ;
        RECT 0.270 1496.700 2917.200 1498.700 ;
        RECT 0.270 1476.260 2918.175 1496.700 ;
        RECT 2.800 1474.260 2918.175 1476.260 ;
        RECT 0.270 1433.420 2918.175 1474.260 ;
        RECT 0.270 1431.420 2917.200 1433.420 ;
        RECT 0.270 1413.020 2918.175 1431.420 ;
        RECT 2.800 1411.020 2918.175 1413.020 ;
        RECT 0.270 1368.140 2918.175 1411.020 ;
        RECT 0.270 1366.140 2917.200 1368.140 ;
        RECT 0.270 1349.780 2918.175 1366.140 ;
        RECT 2.800 1347.780 2918.175 1349.780 ;
        RECT 0.270 1302.860 2918.175 1347.780 ;
        RECT 0.270 1300.860 2917.200 1302.860 ;
        RECT 0.270 1286.540 2918.175 1300.860 ;
        RECT 2.800 1284.540 2918.175 1286.540 ;
        RECT 0.270 1237.580 2918.175 1284.540 ;
        RECT 0.270 1235.580 2917.200 1237.580 ;
        RECT 0.270 1223.300 2918.175 1235.580 ;
        RECT 2.800 1221.300 2918.175 1223.300 ;
        RECT 0.270 1172.300 2918.175 1221.300 ;
        RECT 0.270 1170.300 2917.200 1172.300 ;
        RECT 0.270 1160.060 2918.175 1170.300 ;
        RECT 2.800 1158.060 2918.175 1160.060 ;
        RECT 0.270 1107.020 2918.175 1158.060 ;
        RECT 0.270 1105.020 2917.200 1107.020 ;
        RECT 0.270 1096.820 2918.175 1105.020 ;
        RECT 2.800 1094.820 2918.175 1096.820 ;
        RECT 0.270 1041.740 2918.175 1094.820 ;
        RECT 0.270 1039.740 2917.200 1041.740 ;
        RECT 0.270 1033.580 2918.175 1039.740 ;
        RECT 2.800 1031.580 2918.175 1033.580 ;
        RECT 0.270 976.460 2918.175 1031.580 ;
        RECT 0.270 974.460 2917.200 976.460 ;
        RECT 0.270 970.340 2918.175 974.460 ;
        RECT 2.800 968.340 2918.175 970.340 ;
        RECT 0.270 911.180 2918.175 968.340 ;
        RECT 0.270 909.180 2917.200 911.180 ;
        RECT 0.270 907.100 2918.175 909.180 ;
        RECT 2.800 905.100 2918.175 907.100 ;
        RECT 0.270 845.900 2918.175 905.100 ;
        RECT 0.270 843.900 2917.200 845.900 ;
        RECT 0.270 843.860 2918.175 843.900 ;
        RECT 2.800 841.860 2918.175 843.860 ;
        RECT 0.270 780.620 2918.175 841.860 ;
        RECT 2.800 778.620 2917.200 780.620 ;
        RECT 0.270 717.380 2918.175 778.620 ;
        RECT 2.800 715.380 2918.175 717.380 ;
        RECT 0.270 715.340 2918.175 715.380 ;
        RECT 0.270 713.340 2917.200 715.340 ;
        RECT 0.270 654.140 2918.175 713.340 ;
        RECT 2.800 652.140 2918.175 654.140 ;
        RECT 0.270 650.060 2918.175 652.140 ;
        RECT 0.270 648.060 2917.200 650.060 ;
        RECT 0.270 590.900 2918.175 648.060 ;
        RECT 2.800 588.900 2918.175 590.900 ;
        RECT 0.270 584.780 2918.175 588.900 ;
        RECT 0.270 582.780 2917.200 584.780 ;
        RECT 0.270 527.660 2918.175 582.780 ;
        RECT 2.800 525.660 2918.175 527.660 ;
        RECT 0.270 519.500 2918.175 525.660 ;
        RECT 0.270 517.500 2917.200 519.500 ;
        RECT 0.270 464.420 2918.175 517.500 ;
        RECT 2.800 462.420 2918.175 464.420 ;
        RECT 0.270 454.220 2918.175 462.420 ;
        RECT 0.270 452.220 2917.200 454.220 ;
        RECT 0.270 401.180 2918.175 452.220 ;
        RECT 2.800 399.180 2918.175 401.180 ;
        RECT 0.270 388.940 2918.175 399.180 ;
        RECT 0.270 386.940 2917.200 388.940 ;
        RECT 0.270 337.940 2918.175 386.940 ;
        RECT 2.800 335.940 2918.175 337.940 ;
        RECT 0.270 323.660 2918.175 335.940 ;
        RECT 0.270 321.660 2917.200 323.660 ;
        RECT 0.270 274.700 2918.175 321.660 ;
        RECT 2.800 272.700 2918.175 274.700 ;
        RECT 0.270 258.380 2918.175 272.700 ;
        RECT 0.270 256.380 2917.200 258.380 ;
        RECT 0.270 211.460 2918.175 256.380 ;
        RECT 2.800 209.460 2918.175 211.460 ;
        RECT 0.270 193.100 2918.175 209.460 ;
        RECT 0.270 191.100 2917.200 193.100 ;
        RECT 0.270 148.220 2918.175 191.100 ;
        RECT 2.800 146.220 2918.175 148.220 ;
        RECT 0.270 127.820 2918.175 146.220 ;
        RECT 0.270 125.820 2917.200 127.820 ;
        RECT 0.270 84.980 2918.175 125.820 ;
        RECT 2.800 82.980 2918.175 84.980 ;
        RECT 0.270 62.540 2918.175 82.980 ;
        RECT 0.270 60.540 2917.200 62.540 ;
        RECT 0.270 16.495 2918.175 60.540 ;
      LAYER met4 ;
        RECT 0.295 16.495 2917.945 3499.105 ;
  END
END user_project_wrapper
END LIBRARY

